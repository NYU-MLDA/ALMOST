//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n803_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_;
  XOR2_X1   g000(.A(KEYINPUT99), .B(KEYINPUT0), .Z(new_n202_));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G225gat), .A2(G233gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT85), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT86), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT84), .ZN(new_n218_));
  INV_X1    g017(.A(new_n214_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n216_), .B(new_n218_), .C1(KEYINPUT1), .C2(new_n219_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n214_), .A2(KEYINPUT86), .A3(new_n215_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n209_), .B(new_n211_), .C1(new_n220_), .C2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT87), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n223_), .A2(KEYINPUT3), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n210_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT2), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n209_), .B1(new_n226_), .B2(KEYINPUT88), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT88), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n228_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n225_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n230_));
  OAI22_X1  g029(.A1(new_n224_), .A2(new_n210_), .B1(new_n228_), .B2(KEYINPUT2), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n219_), .B(new_n218_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n222_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G127gat), .B(G134gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G113gat), .B(G120gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n235_), .A2(new_n236_), .ZN(new_n239_));
  MUX2_X1   g038(.A(new_n237_), .B(new_n239_), .S(KEYINPUT83), .Z(new_n240_));
  NOR2_X1   g039(.A1(new_n234_), .A2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT4), .B1(new_n238_), .B2(new_n241_), .ZN(new_n242_));
  OR2_X1    g041(.A1(new_n241_), .A2(KEYINPUT4), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n208_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n234_), .A2(new_n237_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n245_), .B1(new_n240_), .B2(new_n234_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n208_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n207_), .B1(new_n244_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n248_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n241_), .A2(KEYINPUT4), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(new_n246_), .B2(KEYINPUT4), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n250_), .B(new_n206_), .C1(new_n252_), .C2(new_n208_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT100), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n249_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(KEYINPUT100), .B(new_n207_), .C1(new_n244_), .C2(new_n248_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT25), .B(G183gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT26), .B(G190gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT82), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT23), .ZN(new_n264_));
  OR2_X1    g063(.A1(G169gat), .A2(G176gat), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n265_), .A2(KEYINPUT24), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G169gat), .A2(G176gat), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n265_), .A2(KEYINPUT24), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n262_), .A2(new_n264_), .A3(new_n266_), .A4(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n264_), .B1(G183gat), .B2(G190gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT22), .B(G169gat), .ZN(new_n272_));
  INV_X1    g071(.A(G176gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n271_), .A2(new_n267_), .A3(new_n274_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n270_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G227gat), .A2(G233gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XOR2_X1   g077(.A(G71gat), .B(G99gat), .Z(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(KEYINPUT30), .B(G15gat), .Z(new_n281_));
  XNOR2_X1  g080(.A(new_n240_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(KEYINPUT31), .B(G43gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n280_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n280_), .A2(new_n284_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n258_), .A2(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G197gat), .B(G204gat), .Z(new_n289_));
  OR2_X1    g088(.A1(new_n289_), .A2(KEYINPUT21), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(KEYINPUT21), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G211gat), .B(G218gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n291_), .A2(new_n292_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n276_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT20), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G226gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT19), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n297_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT96), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n275_), .B(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n269_), .A2(new_n264_), .A3(new_n266_), .A4(new_n261_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n296_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT97), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT97), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n308_), .A3(new_n296_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n301_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n298_), .B1(new_n276_), .B2(new_n296_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(new_n296_), .B2(new_n305_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n300_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n310_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G8gat), .B(G36gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G64gat), .B(G92gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT27), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n275_), .A2(new_n304_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT20), .B1(new_n295_), .B2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n300_), .B1(new_n297_), .B2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n325_), .B1(new_n312_), .B2(new_n300_), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n320_), .B(KEYINPUT101), .Z(new_n327_));
  AOI21_X1  g126(.A(new_n322_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n321_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n314_), .B(new_n320_), .ZN(new_n330_));
  OAI211_X1 g129(.A(KEYINPUT102), .B(new_n329_), .C1(new_n330_), .C2(KEYINPUT27), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT102), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n330_), .A2(KEYINPUT27), .ZN(new_n333_));
  INV_X1    g132(.A(new_n329_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  XOR2_X1   g134(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n336_));
  AOI21_X1  g135(.A(new_n296_), .B1(new_n233_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(G233gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT91), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n339_), .A2(G228gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(G228gat), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n338_), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT92), .ZN(new_n343_));
  OR2_X1    g142(.A1(new_n337_), .A2(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G78gat), .B(G106gat), .Z(new_n345_));
  NAND2_X1  g144(.A1(new_n233_), .A2(KEYINPUT29), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(new_n295_), .A3(new_n343_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n344_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT94), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(new_n347_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n345_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT95), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n348_), .A2(new_n349_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT95), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n351_), .A2(new_n356_), .A3(new_n352_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n350_), .A2(new_n354_), .A3(new_n355_), .A4(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n233_), .A2(KEYINPUT29), .ZN(new_n359_));
  XOR2_X1   g158(.A(G22gat), .B(G50gat), .Z(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT90), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n359_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n358_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n348_), .A3(new_n353_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n288_), .A2(new_n331_), .A3(new_n335_), .A4(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT33), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n253_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n246_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n206_), .B1(new_n372_), .B2(new_n247_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(new_n252_), .B2(new_n247_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n330_), .A2(new_n371_), .A3(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n253_), .A2(new_n370_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n320_), .A2(KEYINPUT32), .ZN(new_n377_));
  MUX2_X1   g176(.A(new_n326_), .B(new_n315_), .S(new_n377_), .Z(new_n378_));
  OAI22_X1  g177(.A1(new_n375_), .A2(new_n376_), .B1(new_n257_), .B2(new_n378_), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n366_), .A2(new_n367_), .B1(new_n256_), .B2(new_n255_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n333_), .A2(new_n334_), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n379_), .A2(new_n368_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n287_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n369_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(G85gat), .ZN(new_n385_));
  INV_X1    g184(.A(G92gat), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n385_), .A2(new_n386_), .A3(KEYINPUT9), .ZN(new_n387_));
  XOR2_X1   g186(.A(KEYINPUT10), .B(G99gat), .Z(new_n388_));
  INV_X1    g187(.A(G106gat), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G85gat), .B(G92gat), .Z(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT9), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G99gat), .A2(G106gat), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT6), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT64), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT64), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT6), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n393_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n395_), .A2(new_n397_), .A3(new_n393_), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n390_), .B(new_n392_), .C1(new_n398_), .C2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(G99gat), .A2(G106gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT7), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(new_n399_), .B2(new_n398_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT8), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n404_), .A3(new_n391_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT65), .B1(new_n399_), .B2(new_n398_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n393_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n396_), .A2(KEYINPUT6), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n394_), .A2(KEYINPUT64), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT65), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n395_), .A2(new_n397_), .A3(new_n393_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n406_), .A2(new_n413_), .A3(new_n402_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n404_), .B1(new_n414_), .B2(new_n391_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT66), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n405_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  AOI211_X1 g216(.A(KEYINPUT66), .B(new_n404_), .C1(new_n414_), .C2(new_n391_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n400_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G71gat), .B(G78gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G57gat), .B(G64gat), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(KEYINPUT11), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n422_), .B1(KEYINPUT11), .B2(new_n421_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n420_), .A3(KEYINPUT11), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n419_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT68), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n419_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n429_), .A3(KEYINPUT12), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT12), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n419_), .B(new_n426_), .C1(new_n428_), .C2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n425_), .B(new_n400_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G230gat), .A2(G233gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT69), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT69), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n434_), .A2(new_n438_), .A3(new_n435_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n433_), .A2(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n427_), .A2(KEYINPUT67), .A3(new_n434_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n435_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT67), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n419_), .A2(new_n444_), .A3(new_n426_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n442_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n446_));
  XOR2_X1   g245(.A(KEYINPUT70), .B(KEYINPUT5), .Z(new_n447_));
  XNOR2_X1  g246(.A(G120gat), .B(G148gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G176gat), .B(G204gat), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n449_), .B(new_n450_), .Z(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n441_), .A2(new_n446_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n452_), .B1(new_n441_), .B2(new_n446_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n456_), .B(KEYINPUT13), .Z(new_n457_));
  INV_X1    g256(.A(KEYINPUT81), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G29gat), .B(G36gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G43gat), .B(G50gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT15), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G1gat), .B(G8gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT77), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G15gat), .B(G22gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G1gat), .A2(G8gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT14), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n465_), .A2(new_n467_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n464_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n464_), .A2(new_n468_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n462_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n470_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n461_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  MUX2_X1   g273(.A(new_n471_), .B(new_n474_), .S(KEYINPUT80), .Z(new_n475_));
  NAND2_X1  g274(.A1(G229gat), .A2(G233gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n473_), .A2(KEYINPUT79), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n472_), .A2(new_n461_), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n479_), .B(new_n480_), .Z(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n477_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G113gat), .B(G141gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G169gat), .B(G197gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n478_), .A2(new_n482_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n486_), .B1(new_n478_), .B2(new_n482_), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n458_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(KEYINPUT81), .A3(new_n487_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n457_), .A2(new_n494_), .ZN(new_n495_));
  AND2_X1   g294(.A1(new_n384_), .A2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n419_), .A2(new_n462_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G232gat), .A2(G233gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n498_), .B(KEYINPUT34), .Z(new_n499_));
  INV_X1    g298(.A(KEYINPUT35), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n497_), .A2(new_n501_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n461_), .B(new_n400_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n499_), .A2(new_n500_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT72), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n502_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G134gat), .B(G162gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT74), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G190gat), .B(G218gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT36), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT75), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT76), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT71), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n497_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n419_), .A2(new_n462_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT71), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n506_), .A3(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(KEYINPUT73), .A3(new_n501_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT73), .B1(new_n520_), .B2(new_n501_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n507_), .B(new_n515_), .C1(new_n522_), .C2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT37), .ZN(new_n525_));
  INV_X1    g324(.A(new_n523_), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n526_), .A2(new_n521_), .B1(new_n506_), .B2(new_n502_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n511_), .B(KEYINPUT36), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n524_), .B(new_n525_), .C1(new_n527_), .C2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n507_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(new_n528_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n525_), .B1(new_n533_), .B2(new_n524_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n531_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G231gat), .A2(G233gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n425_), .B(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n472_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(G127gat), .B(G155gat), .Z(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(G211gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(KEYINPUT16), .B(G183gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(KEYINPUT68), .A3(KEYINPUT17), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(KEYINPUT17), .B2(new_n543_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n538_), .A2(new_n544_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n548_), .B(KEYINPUT78), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n535_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n496_), .A2(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n552_), .B(KEYINPUT103), .Z(new_n553_));
  OR3_X1    g352(.A1(new_n553_), .A2(G1gat), .A3(new_n257_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT38), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n533_), .A2(new_n524_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n496_), .A2(new_n557_), .A3(new_n548_), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n558_), .B(KEYINPUT104), .Z(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n258_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(G1gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n554_), .A2(new_n555_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n561_), .A3(new_n562_), .ZN(G1324gat));
  AND2_X1   g362(.A1(new_n335_), .A2(new_n331_), .ZN(new_n564_));
  OAI21_X1  g363(.A(G8gat), .B1(new_n558_), .B2(new_n564_), .ZN(new_n565_));
  XOR2_X1   g364(.A(new_n565_), .B(KEYINPUT39), .Z(new_n566_));
  NOR3_X1   g365(.A1(new_n553_), .A2(G8gat), .A3(new_n564_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT40), .ZN(G1325gat));
  NAND2_X1  g368(.A1(new_n559_), .A2(new_n383_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(G15gat), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n571_), .A2(KEYINPUT41), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(KEYINPUT41), .ZN(new_n573_));
  OR3_X1    g372(.A1(new_n552_), .A2(G15gat), .A3(new_n287_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(new_n573_), .A3(new_n574_), .ZN(G1326gat));
  INV_X1    g374(.A(G22gat), .ZN(new_n576_));
  INV_X1    g375(.A(new_n368_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n576_), .B1(new_n559_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT42), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n576_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n552_), .B2(new_n581_), .ZN(G1327gat));
  NAND2_X1  g381(.A1(new_n384_), .A2(new_n535_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n535_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT105), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT43), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n384_), .A2(new_n585_), .A3(KEYINPUT43), .A4(new_n535_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n587_), .A2(new_n495_), .A3(new_n550_), .A4(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT44), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n549_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n592_), .A2(KEYINPUT44), .A3(new_n495_), .A4(new_n588_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n258_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(G29gat), .ZN(new_n595_));
  INV_X1    g394(.A(new_n557_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(new_n550_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n496_), .A2(new_n598_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n257_), .A2(G29gat), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n595_), .B1(new_n599_), .B2(new_n600_), .ZN(G1328gat));
  INV_X1    g400(.A(KEYINPUT46), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n602_), .A2(KEYINPUT108), .ZN(new_n603_));
  INV_X1    g402(.A(new_n564_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n591_), .A2(new_n604_), .A3(new_n593_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(G36gat), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT106), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n611_));
  OR4_X1    g410(.A1(G36gat), .A2(new_n599_), .A3(new_n564_), .A4(new_n611_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n564_), .A2(G36gat), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n611_), .B1(new_n599_), .B2(new_n613_), .ZN(new_n614_));
  AOI22_X1  g413(.A1(new_n612_), .A2(new_n614_), .B1(KEYINPUT108), .B2(new_n602_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n603_), .B1(new_n610_), .B2(new_n615_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n605_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT106), .B1(new_n605_), .B2(G36gat), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n603_), .B(new_n615_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n616_), .A2(new_n620_), .ZN(G1329gat));
  NOR3_X1   g420(.A1(new_n599_), .A2(G43gat), .A3(new_n287_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n591_), .A2(new_n383_), .A3(new_n593_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n623_), .B2(G43gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n624_), .B(new_n625_), .Z(G1330gat));
  NOR2_X1   g425(.A1(new_n368_), .A2(G50gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT110), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n599_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n591_), .A2(new_n577_), .A3(new_n593_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(G50gat), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT111), .Z(G1331gat));
  INV_X1    g431(.A(new_n457_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(new_n493_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n634_), .A2(new_n384_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n635_), .A2(new_n551_), .ZN(new_n636_));
  AOI21_X1  g435(.A(G57gat), .B1(new_n636_), .B2(new_n258_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n635_), .A2(new_n557_), .A3(new_n549_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n258_), .A2(G57gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n637_), .B1(new_n638_), .B2(new_n639_), .ZN(G1332gat));
  INV_X1    g439(.A(G64gat), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n641_), .B1(new_n638_), .B2(new_n604_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT48), .Z(new_n643_));
  NAND3_X1  g442(.A1(new_n636_), .A2(new_n641_), .A3(new_n604_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1333gat));
  INV_X1    g444(.A(G71gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n638_), .B2(new_n383_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT49), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n636_), .A2(new_n646_), .A3(new_n383_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1334gat));
  INV_X1    g449(.A(G78gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n638_), .B2(new_n577_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n636_), .A2(new_n651_), .A3(new_n577_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1335gat));
  AND2_X1   g455(.A1(new_n635_), .A2(new_n598_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n385_), .B1(new_n658_), .B2(new_n257_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n592_), .A2(new_n588_), .A3(new_n634_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n258_), .A2(G85gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n659_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT113), .Z(G1336gat));
  NOR3_X1   g462(.A1(new_n660_), .A2(new_n386_), .A3(new_n564_), .ZN(new_n664_));
  AOI21_X1  g463(.A(G92gat), .B1(new_n657_), .B2(new_n604_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(G1337gat));
  OAI21_X1  g465(.A(G99gat), .B1(new_n660_), .B2(new_n287_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n657_), .A2(new_n388_), .A3(new_n383_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n669_), .B(new_n670_), .Z(G1338gat));
  NAND3_X1  g470(.A1(new_n657_), .A2(new_n389_), .A3(new_n577_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT115), .Z(new_n673_));
  NAND4_X1  g472(.A1(new_n592_), .A2(new_n577_), .A3(new_n588_), .A4(new_n634_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(G106gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT116), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT116), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n674_), .A2(new_n677_), .A3(G106gat), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT52), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n676_), .A2(KEYINPUT52), .A3(new_n678_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n673_), .A2(new_n681_), .A3(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT53), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT53), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n673_), .A2(new_n681_), .A3(new_n685_), .A4(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1339gat));
  NOR2_X1   g486(.A1(new_n457_), .A2(new_n493_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT54), .ZN(new_n689_));
  AOI22_X1  g488(.A1(new_n551_), .A2(new_n688_), .B1(KEYINPUT117), .B2(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n690_), .B1(KEYINPUT117), .B2(new_n689_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT117), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n551_), .A2(new_n688_), .A3(new_n692_), .A4(KEYINPUT54), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n486_), .B1(new_n481_), .B2(new_n476_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n695_), .B1(new_n476_), .B2(new_n475_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n696_), .A2(new_n487_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n697_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT120), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n697_), .B(KEYINPUT120), .C1(new_n454_), .C2(new_n455_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n435_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT55), .B1(new_n433_), .B2(new_n440_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  AOI22_X1  g504(.A1(new_n432_), .A2(new_n430_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT55), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n452_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT118), .B1(new_n708_), .B2(KEYINPUT56), .ZN(new_n709_));
  INV_X1    g508(.A(new_n434_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n711_));
  OAI22_X1  g510(.A1(new_n706_), .A2(KEYINPUT55), .B1(new_n711_), .B2(new_n435_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT55), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n441_), .A2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT56), .B(new_n451_), .C1(new_n712_), .C2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT119), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n433_), .A2(new_n434_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n443_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n441_), .A2(new_n713_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n707_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT119), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n720_), .A2(new_n721_), .A3(KEYINPUT56), .A4(new_n451_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n451_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT118), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT56), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n723_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n709_), .A2(new_n716_), .A3(new_n722_), .A4(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n493_), .A2(new_n453_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n702_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT57), .B1(new_n730_), .B2(new_n596_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT57), .ZN(new_n732_));
  AOI211_X1 g531(.A(KEYINPUT118), .B(KEYINPUT56), .C1(new_n720_), .C2(new_n451_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n724_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n716_), .A2(new_n722_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n728_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n732_), .B(new_n557_), .C1(new_n737_), .C2(new_n702_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n731_), .A2(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n697_), .A2(new_n453_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n715_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT56), .B1(new_n720_), .B2(new_n451_), .ZN(new_n742_));
  OAI211_X1 g541(.A(KEYINPUT58), .B(new_n740_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT121), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n723_), .A2(new_n725_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n715_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT121), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n746_), .A2(new_n747_), .A3(KEYINPUT58), .A4(new_n740_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n740_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT58), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  AND4_X1   g550(.A1(new_n535_), .A2(new_n744_), .A3(new_n748_), .A4(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n739_), .A2(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT122), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n752_), .B1(new_n731_), .B2(new_n738_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n548_), .B1(new_n757_), .B2(KEYINPUT122), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n694_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  NOR4_X1   g558(.A1(new_n604_), .A2(new_n257_), .A3(new_n577_), .A4(new_n287_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT123), .Z(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT124), .B1(new_n759_), .B2(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n691_), .A2(new_n693_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n739_), .A2(KEYINPUT122), .A3(new_n753_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n548_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n757_), .A2(KEYINPUT122), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT124), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n761_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n763_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(G113gat), .B1(new_n772_), .B2(new_n493_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n756_), .A2(new_n758_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n762_), .B1(new_n774_), .B2(new_n764_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT59), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT125), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT125), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(KEYINPUT59), .C1(new_n759_), .C2(new_n762_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n764_), .B1(new_n549_), .B2(new_n757_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT126), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT59), .B1(new_n761_), .B2(new_n781_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n780_), .B(new_n782_), .C1(new_n781_), .C2(new_n761_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n777_), .A2(new_n779_), .A3(new_n783_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n493_), .A2(G113gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n773_), .B1(new_n784_), .B2(new_n785_), .ZN(G1340gat));
  NAND4_X1  g585(.A1(new_n777_), .A2(new_n457_), .A3(new_n779_), .A4(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(G120gat), .ZN(new_n788_));
  INV_X1    g587(.A(G120gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n633_), .B2(KEYINPUT60), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n772_), .B(new_n790_), .C1(KEYINPUT60), .C2(new_n789_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n788_), .A2(new_n791_), .ZN(G1341gat));
  AOI21_X1  g591(.A(G127gat), .B1(new_n772_), .B2(new_n549_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n548_), .A2(G127gat), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n793_), .B1(new_n784_), .B2(new_n794_), .ZN(G1342gat));
  AOI21_X1  g594(.A(G134gat), .B1(new_n772_), .B2(new_n596_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n535_), .A2(G134gat), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n784_), .B2(new_n797_), .ZN(G1343gat));
  NOR2_X1   g597(.A1(new_n759_), .A2(new_n383_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n604_), .A2(new_n257_), .A3(new_n368_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n493_), .A3(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g601(.A1(new_n799_), .A2(new_n457_), .A3(new_n800_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g603(.A1(new_n799_), .A2(new_n549_), .A3(new_n800_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(KEYINPUT61), .B(G155gat), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1346gat));
  AND4_X1   g606(.A1(G162gat), .A2(new_n799_), .A3(new_n535_), .A4(new_n800_), .ZN(new_n808_));
  INV_X1    g607(.A(G162gat), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n799_), .A2(new_n596_), .A3(new_n800_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n808_), .B1(new_n809_), .B2(new_n810_), .ZN(G1347gat));
  NAND3_X1  g610(.A1(new_n604_), .A2(new_n368_), .A3(new_n288_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n780_), .A2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(G169gat), .B1(new_n814_), .B2(new_n494_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT62), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n816_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n814_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(new_n493_), .A3(new_n272_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(new_n818_), .A3(new_n820_), .ZN(G1348gat));
  AOI21_X1  g620(.A(G176gat), .B1(new_n819_), .B2(new_n457_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n812_), .A2(new_n273_), .A3(new_n633_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n769_), .B2(new_n823_), .ZN(G1349gat));
  NOR3_X1   g623(.A1(new_n814_), .A2(new_n259_), .A3(new_n766_), .ZN(new_n825_));
  INV_X1    g624(.A(G183gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n769_), .A2(new_n549_), .A3(new_n813_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(G1350gat));
  OAI21_X1  g627(.A(G190gat), .B1(new_n814_), .B2(new_n584_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n596_), .A2(new_n260_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n814_), .B2(new_n830_), .ZN(G1351gat));
  NOR3_X1   g630(.A1(new_n564_), .A2(new_n258_), .A3(new_n368_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n769_), .A2(new_n493_), .A3(new_n287_), .A4(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(G197gat), .ZN(new_n834_));
  OR3_X1    g633(.A1(new_n833_), .A2(KEYINPUT127), .A3(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT127), .B1(new_n833_), .B2(new_n834_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n834_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(G1352gat));
  AND3_X1   g637(.A1(new_n769_), .A2(new_n287_), .A3(new_n832_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n457_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g640(.A(KEYINPUT63), .B(G211gat), .C1(new_n839_), .C2(new_n548_), .ZN(new_n842_));
  XOR2_X1   g641(.A(KEYINPUT63), .B(G211gat), .Z(new_n843_));
  AND3_X1   g642(.A1(new_n839_), .A2(new_n548_), .A3(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1354gat));
  AOI21_X1  g644(.A(G218gat), .B1(new_n839_), .B2(new_n596_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n535_), .A2(G218gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n839_), .B2(new_n847_), .ZN(G1355gat));
endmodule


