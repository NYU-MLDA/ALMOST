//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT10), .B(G99gat), .Z(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G106gat), .Z(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G85gat), .B(G92gat), .Z(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n207_));
  INV_X1    g006(.A(G85gat), .ZN(new_n208_));
  INV_X1    g007(.A(G92gat), .ZN(new_n209_));
  OR3_X1    g008(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT9), .ZN(new_n210_));
  AND3_X1   g009(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n205_), .A2(new_n207_), .A3(new_n210_), .A4(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT8), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT66), .B1(new_n211_), .B2(new_n212_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT66), .ZN(new_n220_));
  NAND3_X1  g019(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n223_));
  NOR2_X1   g022(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n224_));
  OAI22_X1  g023(.A1(new_n223_), .A2(new_n224_), .B1(G99gat), .B2(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n226_));
  INV_X1    g025(.A(G99gat), .ZN(new_n227_));
  INV_X1    g026(.A(G106gat), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n216_), .A2(new_n222_), .A3(new_n225_), .A4(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n215_), .B1(new_n230_), .B2(new_n206_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n206_), .A2(new_n215_), .ZN(new_n232_));
  OR2_X1    g031(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n233_), .A2(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n229_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n232_), .B1(new_n236_), .B2(new_n213_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n214_), .B1(new_n231_), .B2(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G57gat), .B(G64gat), .Z(new_n239_));
  INV_X1    g038(.A(KEYINPUT11), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G57gat), .B(G64gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT11), .ZN(new_n243_));
  XOR2_X1   g042(.A(G71gat), .B(G78gat), .Z(new_n244_));
  NAND3_X1  g043(.A1(new_n241_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n243_), .A2(new_n244_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n238_), .A2(new_n248_), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n247_), .B(new_n214_), .C1(new_n231_), .C2(new_n237_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n202_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n238_), .A2(KEYINPUT67), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n253_), .B(new_n214_), .C1(new_n231_), .C2(new_n237_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n248_), .A2(KEYINPUT12), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n250_), .A2(KEYINPUT12), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n255_), .A2(new_n257_), .B1(new_n249_), .B2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n251_), .B1(new_n259_), .B2(new_n202_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G176gat), .B(G204gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G120gat), .B(G148gat), .ZN(new_n264_));
  XOR2_X1   g063(.A(new_n263_), .B(new_n264_), .Z(new_n265_));
  XNOR2_X1  g064(.A(new_n260_), .B(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n266_), .B(KEYINPUT13), .Z(new_n267_));
  XNOR2_X1  g066(.A(G113gat), .B(G141gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G169gat), .B(G197gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(KEYINPUT72), .B(G8gat), .Z(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(G1gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(KEYINPUT14), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT73), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G15gat), .B(G22gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G1gat), .B(G8gat), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n274_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G29gat), .B(G36gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G43gat), .B(G50gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n284_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n279_), .A2(new_n280_), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G229gat), .A2(G233gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT81), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n285_), .A2(new_n289_), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n284_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n279_), .A2(new_n294_), .A3(new_n280_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n290_), .B1(new_n285_), .B2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n270_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n296_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n270_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n292_), .A3(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n297_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G183gat), .B(G211gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G127gat), .B(G155gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n308_), .B(KEYINPUT76), .Z(new_n309_));
  AND2_X1   g108(.A1(new_n279_), .A2(new_n280_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G231gat), .A2(G233gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n247_), .B(new_n311_), .Z(new_n312_));
  AND2_X1   g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n310_), .A2(new_n312_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n309_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n281_), .B(new_n312_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT77), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n306_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT17), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT78), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n315_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n321_), .B1(new_n315_), .B2(new_n320_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n267_), .A2(new_n301_), .A3(new_n324_), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n325_), .A2(KEYINPUT106), .ZN(new_n326_));
  INV_X1    g125(.A(G155gat), .ZN(new_n327_));
  INV_X1    g126(.A(G162gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(G141gat), .ZN(new_n330_));
  INV_X1    g129(.A(G148gat), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n329_), .A2(KEYINPUT1), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G155gat), .B(G162gat), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n332_), .B(new_n333_), .C1(KEYINPUT1), .C2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT89), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n330_), .A2(new_n331_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(KEYINPUT90), .A2(KEYINPUT3), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n333_), .A2(KEYINPUT2), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT2), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(G141gat), .A3(G148gat), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n341_), .A2(new_n343_), .B1(KEYINPUT90), .B2(KEYINPUT3), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT91), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT92), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n334_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT91), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n340_), .A2(new_n349_), .A3(new_n344_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n334_), .A2(new_n347_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n346_), .A2(new_n348_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n337_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G127gat), .B(G134gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G113gat), .B(G120gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT88), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n354_), .A2(new_n355_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n357_), .B(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n353_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G225gat), .A2(G233gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n358_), .A2(new_n356_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n337_), .A2(new_n352_), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n361_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G1gat), .B(G29gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(new_n208_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT0), .B(G57gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n359_), .B1(new_n337_), .B2(new_n352_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n371_), .A2(KEYINPUT4), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n361_), .A2(new_n364_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n372_), .B1(new_n373_), .B2(KEYINPUT4), .ZN(new_n374_));
  XOR2_X1   g173(.A(new_n362_), .B(KEYINPUT100), .Z(new_n375_));
  OAI211_X1 g174(.A(new_n365_), .B(new_n370_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT33), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT101), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XOR2_X1   g182(.A(G211gat), .B(G218gat), .Z(new_n384_));
  INV_X1    g183(.A(KEYINPUT94), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G211gat), .B(G218gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT94), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(KEYINPUT95), .A3(new_n388_), .ZN(new_n389_));
  XOR2_X1   g188(.A(G197gat), .B(G204gat), .Z(new_n390_));
  AND3_X1   g189(.A1(new_n389_), .A2(KEYINPUT21), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n390_), .B1(new_n389_), .B2(KEYINPUT21), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n387_), .B(new_n385_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT21), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n391_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT23), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n397_), .A2(G183gat), .A3(G190gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT83), .ZN(new_n399_));
  INV_X1    g198(.A(G183gat), .ZN(new_n400_));
  INV_X1    g199(.A(G190gat), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT23), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n401_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT22), .B(G169gat), .ZN(new_n407_));
  INV_X1    g206(.A(G176gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(new_n406_), .A3(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT26), .B(G190gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT25), .B(G183gat), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n411_), .A2(new_n412_), .B1(new_n402_), .B2(new_n398_), .ZN(new_n413_));
  NOR3_X1   g212(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n414_), .B1(new_n416_), .B2(new_n406_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n413_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n410_), .A2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n396_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n389_), .A2(KEYINPUT21), .ZN(new_n421_));
  INV_X1    g220(.A(new_n390_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n393_), .A2(new_n394_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n389_), .A2(KEYINPUT21), .A3(new_n390_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT25), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n427_), .B1(new_n428_), .B2(G183gat), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n411_), .B(new_n429_), .C1(new_n412_), .C2(new_n427_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n403_), .A2(new_n417_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n402_), .A2(new_n398_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(new_n404_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT85), .ZN(new_n434_));
  NOR3_X1   g233(.A1(new_n434_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n435_));
  OAI21_X1  g234(.A(G169gat), .B1(new_n435_), .B2(G176gat), .ZN(new_n436_));
  INV_X1    g235(.A(G169gat), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n437_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n438_), .B1(new_n407_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n434_), .A2(new_n408_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n433_), .B(new_n436_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n431_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT20), .B1(new_n426_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n383_), .B1(new_n420_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n396_), .A2(new_n419_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n426_), .A2(new_n444_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n383_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n447_), .A2(KEYINPUT20), .A3(new_n448_), .A4(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n446_), .A2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G64gat), .B(G92gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G8gat), .B(G36gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n451_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n446_), .A2(new_n456_), .A3(new_n450_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n362_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n337_), .A2(new_n352_), .A3(new_n363_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT4), .B1(new_n462_), .B2(new_n371_), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n371_), .A2(KEYINPUT4), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n461_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n373_), .A2(new_n375_), .ZN(new_n466_));
  NOR3_X1   g265(.A1(new_n465_), .A2(new_n370_), .A3(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n460_), .A2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n375_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n365_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(KEYINPUT33), .A3(new_n370_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n376_), .A2(KEYINPUT101), .A3(new_n377_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n380_), .A2(new_n468_), .A3(new_n472_), .A4(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n369_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n376_), .ZN(new_n476_));
  AND4_X1   g275(.A1(KEYINPUT20), .A2(new_n447_), .A3(new_n383_), .A4(new_n448_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n478_), .B1(new_n396_), .B2(new_n443_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n426_), .A2(new_n410_), .A3(new_n418_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n383_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n477_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n457_), .A2(KEYINPUT32), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n451_), .A2(new_n483_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n476_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n474_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n443_), .A2(KEYINPUT30), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT30), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n431_), .A2(new_n489_), .A3(new_n442_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G227gat), .A2(G233gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT86), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G15gat), .B(G43gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G71gat), .B(G99gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  OR3_X1    g296(.A1(new_n491_), .A2(KEYINPUT87), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n490_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n489_), .B1(new_n431_), .B2(new_n442_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT87), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT87), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n488_), .A2(new_n502_), .A3(new_n490_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n503_), .A3(new_n497_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n359_), .B(KEYINPUT31), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n498_), .A2(new_n504_), .A3(new_n506_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT29), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(new_n337_), .B2(new_n352_), .ZN(new_n513_));
  OAI211_X1 g312(.A(G228gat), .B(G233gat), .C1(new_n513_), .C2(new_n426_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n426_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G228gat), .A2(G233gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G22gat), .B(G50gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n521_), .B1(new_n353_), .B2(KEYINPUT29), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G78gat), .B(G106gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n523_), .B(KEYINPUT96), .Z(new_n524_));
  OR2_X1    g323(.A1(new_n524_), .A2(KEYINPUT97), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n337_), .A2(new_n352_), .A3(new_n512_), .A4(new_n520_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n522_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n524_), .B1(new_n522_), .B2(new_n526_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n514_), .B(new_n517_), .C1(new_n528_), .C2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n517_), .A2(new_n514_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n522_), .A2(new_n526_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n524_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n531_), .A2(new_n527_), .A3(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n511_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT102), .B1(new_n482_), .B2(new_n457_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT102), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n540_), .B(new_n456_), .C1(new_n477_), .C2(new_n481_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n539_), .A2(KEYINPUT27), .A3(new_n458_), .A4(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT103), .B(KEYINPUT27), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n446_), .A2(new_n456_), .A3(new_n450_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n456_), .B1(new_n446_), .B2(new_n450_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n543_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT104), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n460_), .A2(KEYINPUT104), .A3(new_n543_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n542_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n530_), .A2(new_n535_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n530_), .A2(new_n535_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n476_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n487_), .A2(new_n538_), .B1(new_n551_), .B2(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n287_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G232gat), .A2(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT35), .ZN(new_n562_));
  OR2_X1    g361(.A1(new_n561_), .A2(KEYINPUT35), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n238_), .A2(new_n294_), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n558_), .A2(new_n562_), .A3(new_n563_), .A4(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n564_), .ZN(new_n566_));
  OAI211_X1 g365(.A(KEYINPUT35), .B(new_n561_), .C1(new_n566_), .C2(new_n557_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G190gat), .B(G218gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G134gat), .B(G162gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n569_), .B(new_n570_), .Z(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n572_), .A2(KEYINPUT36), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n568_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(KEYINPUT36), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n568_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT107), .Z(new_n578_));
  NOR2_X1   g377(.A1(new_n556_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n325_), .A2(KEYINPUT106), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n326_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n476_), .ZN(new_n582_));
  OAI21_X1  g381(.A(G1gat), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT79), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n584_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n315_), .A2(new_n320_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT78), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n315_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(KEYINPUT79), .A3(new_n588_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n585_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT37), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(new_n576_), .B2(KEYINPUT71), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n577_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n574_), .B(new_n576_), .C1(KEYINPUT71), .C2(new_n591_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n590_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n267_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT80), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n556_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n301_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n595_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n585_), .A2(new_n589_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n267_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n601_), .B1(new_n605_), .B2(KEYINPUT80), .ZN(new_n606_));
  INV_X1    g405(.A(G1gat), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n600_), .A2(new_n606_), .A3(new_n607_), .A4(new_n476_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n608_), .A2(KEYINPUT105), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT38), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(KEYINPUT105), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n610_), .B1(new_n609_), .B2(new_n611_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n583_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT108), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OAI211_X1 g415(.A(KEYINPUT108), .B(new_n583_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1324gat));
  OAI21_X1  g417(.A(G8gat), .B1(new_n581_), .B2(new_n551_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n619_), .A2(KEYINPUT39), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(KEYINPUT39), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n600_), .A2(new_n606_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n551_), .A2(new_n271_), .ZN(new_n623_));
  AOI22_X1  g422(.A1(new_n620_), .A2(new_n621_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n624_), .B(new_n625_), .Z(G1325gat));
  INV_X1    g425(.A(G15gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n622_), .A2(new_n627_), .A3(new_n510_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT110), .Z(new_n629_));
  OAI21_X1  g428(.A(G15gat), .B1(new_n581_), .B2(new_n511_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT41), .Z(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(G1326gat));
  INV_X1    g431(.A(G22gat), .ZN(new_n633_));
  INV_X1    g432(.A(new_n536_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n622_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n581_), .A2(new_n536_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT42), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n636_), .A2(new_n637_), .A3(G22gat), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n637_), .B1(new_n636_), .B2(G22gat), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n635_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT111), .ZN(G1327gat));
  NOR2_X1   g441(.A1(new_n556_), .A2(new_n577_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n597_), .A2(new_n590_), .A3(new_n601_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT114), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n643_), .A2(KEYINPUT114), .A3(new_n644_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n476_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n652_), .A2(KEYINPUT113), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(KEYINPUT113), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT43), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n537_), .B1(new_n474_), .B2(new_n486_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n554_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n582_), .B1(new_n658_), .B2(new_n552_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n550_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n656_), .B(new_n602_), .C1(new_n657_), .C2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT112), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n476_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n376_), .A2(new_n377_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n664_), .A2(new_n460_), .A3(new_n467_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n376_), .A2(KEYINPUT101), .A3(new_n377_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT101), .B1(new_n376_), .B2(new_n377_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n663_), .B1(new_n665_), .B2(new_n668_), .ZN(new_n669_));
  OAI22_X1  g468(.A1(new_n669_), .A2(new_n537_), .B1(new_n550_), .B2(new_n659_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT112), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n670_), .A2(new_n671_), .A3(new_n656_), .A4(new_n602_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT43), .B1(new_n556_), .B2(new_n595_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n662_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  AOI211_X1 g473(.A(new_n653_), .B(new_n655_), .C1(new_n674_), .C2(new_n644_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n674_), .A2(KEYINPUT113), .A3(new_n652_), .A4(new_n644_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(new_n582_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n651_), .B1(new_n679_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g479(.A(G36gat), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n647_), .A2(new_n681_), .A3(new_n550_), .A4(new_n648_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT45), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n678_), .A2(new_n551_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n684_), .B2(new_n681_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(KEYINPUT46), .B(new_n683_), .C1(new_n684_), .C2(new_n681_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1329gat));
  OAI211_X1 g488(.A(G43gat), .B(new_n510_), .C1(new_n675_), .C2(new_n677_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT115), .ZN(new_n691_));
  INV_X1    g490(.A(G43gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n692_), .B1(new_n649_), .B2(new_n511_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n653_), .B1(new_n674_), .B2(new_n644_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n654_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n676_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT115), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n696_), .A2(new_n697_), .A3(G43gat), .A4(new_n510_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n691_), .A2(new_n693_), .A3(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT47), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n691_), .A2(new_n698_), .A3(new_n701_), .A4(new_n693_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1330gat));
  AOI21_X1  g502(.A(G50gat), .B1(new_n650_), .B2(new_n634_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n678_), .A2(new_n536_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(G50gat), .ZN(G1331gat));
  NAND4_X1  g505(.A1(new_n579_), .A2(new_n597_), .A3(new_n601_), .A4(new_n590_), .ZN(new_n707_));
  INV_X1    g506(.A(G57gat), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n582_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n596_), .A2(new_n267_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT116), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n556_), .A2(new_n301_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT117), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n711_), .A2(KEYINPUT117), .A3(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n708_), .B1(new_n717_), .B2(new_n582_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT118), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n718_), .A2(new_n719_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n709_), .B1(new_n720_), .B2(new_n721_), .ZN(G1332gat));
  OAI21_X1  g521(.A(G64gat), .B1(new_n707_), .B2(new_n551_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT48), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n551_), .A2(G64gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n717_), .B2(new_n725_), .ZN(G1333gat));
  OAI21_X1  g525(.A(G71gat), .B1(new_n707_), .B2(new_n511_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT49), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n511_), .A2(G71gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n717_), .B2(new_n729_), .ZN(G1334gat));
  OAI21_X1  g529(.A(G78gat), .B1(new_n707_), .B2(new_n536_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT50), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n536_), .A2(G78gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n717_), .B2(new_n733_), .ZN(G1335gat));
  NOR3_X1   g533(.A1(new_n590_), .A2(new_n267_), .A3(new_n301_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n643_), .A2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n208_), .B1(new_n736_), .B2(new_n582_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT119), .Z(new_n738_));
  XNOR2_X1  g537(.A(new_n735_), .B(KEYINPUT120), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n674_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT121), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n741_), .A2(new_n582_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n738_), .B1(new_n742_), .B2(G85gat), .ZN(G1336gat));
  OAI21_X1  g542(.A(G92gat), .B1(new_n741_), .B2(new_n551_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n736_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n745_), .A2(new_n209_), .A3(new_n550_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1337gat));
  OAI21_X1  g546(.A(G99gat), .B1(new_n740_), .B2(new_n511_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(new_n203_), .A3(new_n510_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g550(.A1(new_n745_), .A2(new_n204_), .A3(new_n634_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G106gat), .B1(new_n740_), .B2(new_n536_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(KEYINPUT52), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(KEYINPUT52), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n752_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g556(.A1(new_n604_), .A2(KEYINPUT54), .A3(new_n267_), .A4(new_n601_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n590_), .A2(new_n267_), .A3(new_n601_), .A4(new_n595_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n758_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT58), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n258_), .A2(new_n249_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n256_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT122), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n255_), .A2(new_n257_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT122), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n258_), .A2(new_n249_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n767_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n202_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n766_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(KEYINPUT123), .ZN(new_n773_));
  AND4_X1   g572(.A1(KEYINPUT55), .A2(new_n767_), .A3(new_n202_), .A4(new_n769_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT55), .B1(new_n259_), .B2(new_n202_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT123), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n766_), .A2(new_n770_), .A3(new_n777_), .A4(new_n771_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n773_), .A2(new_n776_), .A3(new_n778_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n265_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT56), .B1(new_n779_), .B2(new_n265_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT124), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n285_), .A2(new_n295_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n291_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n291_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n285_), .A2(new_n289_), .A3(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n270_), .A3(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n300_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n265_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n260_), .A2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n789_), .A2(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n779_), .A2(new_n782_), .A3(KEYINPUT56), .A4(new_n265_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n763_), .B1(new_n783_), .B2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n779_), .A2(new_n265_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n265_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(KEYINPUT124), .A3(new_n800_), .ZN(new_n801_));
  NAND4_X1  g600(.A1(new_n801_), .A2(KEYINPUT58), .A3(new_n794_), .A4(new_n793_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n796_), .A2(new_n602_), .A3(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n792_), .B1(new_n297_), .B2(new_n300_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n789_), .A2(new_n266_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n804_), .B1(new_n809_), .B2(new_n577_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n577_), .ZN(new_n811_));
  AOI211_X1 g610(.A(KEYINPUT57), .B(new_n811_), .C1(new_n806_), .C2(new_n808_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n803_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n324_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n762_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n550_), .A2(new_n582_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n552_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(G113gat), .B1(new_n818_), .B2(new_n301_), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT59), .B1(new_n815_), .B2(new_n817_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n817_), .A2(KEYINPUT59), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n301_), .A2(new_n791_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n577_), .B1(new_n823_), .B2(new_n807_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT57), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n809_), .A2(new_n804_), .A3(new_n577_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n590_), .B1(new_n827_), .B2(new_n803_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n821_), .B1(new_n828_), .B2(new_n762_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n820_), .A2(new_n829_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n301_), .A2(G113gat), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n819_), .B1(new_n830_), .B2(new_n831_), .ZN(G1340gat));
  INV_X1    g631(.A(new_n817_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT60), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n267_), .B2(G120gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n324_), .B1(new_n827_), .B2(new_n803_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n833_), .B(new_n835_), .C1(new_n836_), .C2(new_n762_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n820_), .A2(new_n597_), .A3(new_n829_), .A4(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G120gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n818_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT125), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT125), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n839_), .A2(new_n843_), .A3(new_n840_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1341gat));
  AOI21_X1  g644(.A(G127gat), .B1(new_n818_), .B2(new_n590_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n324_), .A2(G127gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n830_), .B2(new_n847_), .ZN(G1342gat));
  AOI21_X1  g647(.A(G134gat), .B1(new_n818_), .B2(new_n578_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n602_), .A2(G134gat), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n830_), .B2(new_n850_), .ZN(G1343gat));
  NOR2_X1   g650(.A1(new_n815_), .A2(new_n554_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n816_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n853_), .A2(new_n601_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(new_n330_), .ZN(G1344gat));
  NOR2_X1   g654(.A1(new_n853_), .A2(new_n267_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(new_n331_), .ZN(G1345gat));
  OAI21_X1  g656(.A(G155gat), .B1(new_n853_), .B2(new_n603_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n852_), .A2(new_n327_), .A3(new_n590_), .A4(new_n816_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n858_), .A2(new_n861_), .A3(new_n859_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1346gat));
  NOR3_X1   g664(.A1(new_n853_), .A2(new_n328_), .A3(new_n595_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n853_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n578_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n866_), .B1(new_n328_), .B2(new_n868_), .ZN(G1347gat));
  NAND2_X1  g668(.A1(new_n813_), .A2(new_n603_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n870_), .A2(new_n761_), .A3(new_n758_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n551_), .A2(new_n476_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n553_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n871_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n437_), .B1(new_n875_), .B2(new_n301_), .ZN(new_n876_));
  AND4_X1   g675(.A1(new_n301_), .A2(new_n871_), .A3(new_n407_), .A4(new_n874_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT62), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(KEYINPUT62), .B2(new_n876_), .ZN(G1348gat));
  AOI21_X1  g678(.A(G176gat), .B1(new_n875_), .B2(new_n597_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n815_), .A2(new_n408_), .A3(new_n267_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n874_), .B2(new_n881_), .ZN(G1349gat));
  NOR2_X1   g681(.A1(new_n814_), .A2(new_n412_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n590_), .B(new_n874_), .C1(new_n836_), .C2(new_n762_), .ZN(new_n884_));
  AOI22_X1  g683(.A1(new_n875_), .A2(new_n883_), .B1(new_n884_), .B2(new_n400_), .ZN(G1350gat));
  NAND3_X1  g684(.A1(new_n875_), .A2(new_n578_), .A3(new_n411_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n875_), .A2(new_n602_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n887_), .B2(new_n401_), .ZN(G1351gat));
  OAI211_X1 g687(.A(new_n658_), .B(new_n872_), .C1(new_n836_), .C2(new_n762_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n301_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g691(.A1(new_n890_), .A2(new_n597_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g693(.A1(new_n889_), .A2(new_n814_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT127), .ZN(new_n896_));
  NAND2_X1  g695(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n895_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n896_), .B1(new_n895_), .B2(new_n897_), .ZN(new_n900_));
  OAI22_X1  g699(.A1(new_n899_), .A2(new_n900_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n901_));
  INV_X1    g700(.A(new_n900_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n902_), .A2(new_n903_), .A3(new_n898_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n904_), .ZN(G1354gat));
  AND3_X1   g704(.A1(new_n890_), .A2(G218gat), .A3(new_n602_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G218gat), .B1(new_n890_), .B2(new_n578_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(new_n907_), .ZN(G1355gat));
endmodule


