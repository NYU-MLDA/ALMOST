//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n939_;
  INV_X1    g000(.A(G204gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(new_n202_), .A2(G197gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(KEYINPUT80), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT80), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G204gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n203_), .B1(new_n207_), .B2(G197gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT21), .B1(new_n208_), .B2(KEYINPUT83), .ZN(new_n209_));
  XOR2_X1   g008(.A(G211gat), .B(G218gat), .Z(new_n210_));
  INV_X1    g009(.A(new_n203_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT80), .B(G204gat), .ZN(new_n212_));
  INV_X1    g011(.A(G197gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n211_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT83), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n210_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n209_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n218_));
  INV_X1    g017(.A(G183gat), .ZN(new_n219_));
  INV_X1    g018(.A(G190gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n221_), .B(new_n222_), .C1(G183gat), .C2(G190gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT22), .B(G169gat), .Z(new_n225_));
  OAI211_X1 g024(.A(new_n223_), .B(new_n224_), .C1(G176gat), .C2(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n221_), .A2(new_n222_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT25), .B(G183gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  OR2_X1    g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n231_), .A2(KEYINPUT24), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(KEYINPUT24), .A3(new_n224_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n227_), .A2(new_n230_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n226_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(G197gat), .B1(new_n204_), .B2(new_n206_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT21), .B1(new_n213_), .B2(new_n202_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT81), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT81), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT21), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n241_), .B1(G197gat), .B2(G204gat), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n240_), .B(new_n242_), .C1(new_n212_), .C2(G197gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n210_), .B1(new_n208_), .B2(new_n241_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT82), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n246_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n217_), .B(new_n236_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n209_), .A2(new_n216_), .ZN(new_n250_));
  AND2_X1   g049(.A1(new_n239_), .A2(new_n243_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n210_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n252_), .B1(new_n214_), .B2(KEYINPUT21), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT82), .B1(new_n251_), .B2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n250_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT26), .B1(new_n220_), .B2(KEYINPUT75), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT26), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G190gat), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n229_), .B(new_n257_), .C1(KEYINPUT75), .C2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n260_), .A2(new_n227_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(new_n226_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n249_), .B(KEYINPUT20), .C1(new_n256_), .C2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G226gat), .A2(G233gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT19), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n217_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n235_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n217_), .B(new_n263_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n270_), .A2(KEYINPUT20), .A3(new_n266_), .A4(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G8gat), .B(G36gat), .ZN(new_n274_));
  INV_X1    g073(.A(G92gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT18), .B(G64gat), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n276_), .B(new_n277_), .Z(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n273_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n268_), .A2(new_n272_), .A3(new_n278_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(KEYINPUT86), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT27), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT86), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n273_), .A2(new_n284_), .A3(new_n279_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  AND4_X1   g085(.A1(KEYINPUT20), .A2(new_n270_), .A3(new_n267_), .A4(new_n271_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT93), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n226_), .A2(new_n288_), .A3(new_n234_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n217_), .B(new_n289_), .C1(new_n247_), .C2(new_n248_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n236_), .A2(new_n288_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT20), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT94), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n269_), .A2(new_n262_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT94), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n295_), .B(KEYINPUT20), .C1(new_n290_), .C2(new_n291_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n293_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n287_), .B1(new_n297_), .B2(new_n266_), .ZN(new_n298_));
  OAI211_X1 g097(.A(KEYINPUT27), .B(new_n280_), .C1(new_n298_), .C2(new_n279_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n286_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT96), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G78gat), .B(G106gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT84), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT79), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT1), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n306_), .B1(G155gat), .B2(G162gat), .ZN(new_n307_));
  NOR2_X1   g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n305_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(G155gat), .A3(G162gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n308_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT1), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n311_), .A2(new_n313_), .A3(KEYINPUT77), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n309_), .A2(new_n310_), .A3(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(G141gat), .B(G148gat), .Z(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(G141gat), .ZN(new_n318_));
  INV_X1    g117(.A(G148gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(new_n319_), .A3(KEYINPUT78), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT3), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT3), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n322_), .A2(new_n318_), .A3(new_n319_), .A4(KEYINPUT78), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT2), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n324_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n321_), .A2(new_n323_), .A3(new_n325_), .A4(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n327_), .A2(new_n312_), .A3(new_n311_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n317_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT29), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n269_), .A2(new_n304_), .A3(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n304_), .B1(new_n269_), .B2(new_n330_), .ZN(new_n332_));
  INV_X1    g131(.A(G228gat), .ZN(new_n333_));
  INV_X1    g132(.A(G233gat), .ZN(new_n334_));
  OAI22_X1  g133(.A1(new_n331_), .A2(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n269_), .A2(new_n330_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT79), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n333_), .A2(new_n334_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n269_), .A2(new_n304_), .A3(new_n330_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n303_), .B1(new_n335_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n329_), .A2(KEYINPUT29), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n343_), .B(KEYINPUT28), .Z(new_n344_));
  XNOR2_X1  g143(.A(G22gat), .B(G50gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT85), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n335_), .A2(new_n340_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n302_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n347_), .B1(new_n335_), .B2(new_n340_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n342_), .B(new_n346_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n351_));
  XOR2_X1   g150(.A(KEYINPUT88), .B(KEYINPUT0), .Z(new_n352_));
  XNOR2_X1  g151(.A(G1gat), .B(G29gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G57gat), .B(G85gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT87), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G127gat), .B(G134gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G113gat), .B(G120gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n329_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n317_), .A2(new_n328_), .A3(new_n363_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(KEYINPUT4), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n363_), .B1(new_n317_), .B2(new_n328_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n360_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n317_), .A2(new_n328_), .A3(new_n363_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n360_), .B1(new_n372_), .B2(new_n368_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n357_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n363_), .B(KEYINPUT31), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G227gat), .A2(G233gat), .ZN(new_n377_));
  INV_X1    g176(.A(G15gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(G43gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G71gat), .B(G99gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n383_), .B1(new_n261_), .B2(new_n226_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT76), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n261_), .A2(new_n226_), .A3(new_n383_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n386_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n382_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n387_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT76), .B1(new_n392_), .B2(new_n384_), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n380_), .B(new_n381_), .Z(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n376_), .B1(new_n391_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n394_), .B1(new_n393_), .B2(new_n388_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n390_), .A2(new_n382_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n376_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n397_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n371_), .A2(new_n374_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n356_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT95), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(KEYINPUT95), .A3(new_n356_), .ZN(new_n406_));
  AND4_X1   g205(.A1(new_n375_), .A2(new_n401_), .A3(new_n405_), .A4(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n346_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n335_), .A2(new_n303_), .A3(new_n340_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n408_), .B1(new_n409_), .B2(new_n341_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n351_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT96), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n286_), .A2(new_n299_), .A3(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n301_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT97), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT97), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n301_), .A2(new_n411_), .A3(new_n416_), .A4(new_n413_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n367_), .A2(new_n360_), .A3(new_n370_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT91), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n372_), .A2(new_n368_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n357_), .B1(new_n421_), .B2(new_n359_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n367_), .A2(KEYINPUT91), .A3(new_n360_), .A4(new_n370_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n420_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NOR3_X1   g223(.A1(new_n372_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n370_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n359_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n356_), .B1(new_n427_), .B2(new_n373_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT90), .B1(new_n428_), .B2(KEYINPUT33), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT33), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n375_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n424_), .B1(new_n429_), .B2(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(KEYINPUT33), .B(new_n357_), .C1(new_n371_), .C2(new_n374_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT89), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n281_), .A2(KEYINPUT86), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n278_), .B1(new_n268_), .B2(new_n272_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n285_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n433_), .B(new_n436_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT92), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n405_), .A2(new_n375_), .A3(new_n406_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n279_), .A2(KEYINPUT32), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n273_), .A2(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n443_), .B(new_n445_), .C1(new_n298_), .C2(new_n444_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n282_), .A2(new_n285_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT92), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(new_n436_), .A4(new_n433_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n442_), .A2(new_n446_), .A3(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n351_), .A2(new_n410_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n443_), .B1(new_n351_), .B2(new_n410_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n300_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n450_), .A2(new_n452_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n415_), .B(new_n417_), .C1(new_n455_), .C2(new_n401_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G230gat), .A2(G233gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G85gat), .B(G92gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT9), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT9), .ZN(new_n461_));
  INV_X1    g260(.A(G85gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n461_), .B1(new_n462_), .B2(new_n275_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n460_), .A2(KEYINPUT64), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G99gat), .A2(G106gat), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT10), .B(G99gat), .ZN(new_n470_));
  OR2_X1    g269(.A1(new_n470_), .A2(G106gat), .ZN(new_n471_));
  OR4_X1    g270(.A1(KEYINPUT64), .A2(new_n461_), .A3(new_n462_), .A4(new_n275_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n464_), .A2(new_n469_), .A3(new_n471_), .A4(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT8), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT7), .ZN(new_n475_));
  INV_X1    g274(.A(G99gat), .ZN(new_n476_));
  INV_X1    g275(.A(G106gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n478_), .A2(new_n467_), .A3(new_n468_), .A4(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n459_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n474_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n480_), .A2(new_n474_), .A3(new_n481_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n473_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G57gat), .B(G64gat), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n485_), .A2(KEYINPUT11), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT65), .B(G71gat), .Z(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(G78gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(KEYINPUT11), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT65), .B(G71gat), .ZN(new_n490_));
  INV_X1    g289(.A(G78gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n486_), .A2(new_n488_), .A3(new_n489_), .A4(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n489_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n490_), .A2(new_n491_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n490_), .A2(new_n491_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n493_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n484_), .A2(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n498_), .B(new_n473_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(KEYINPUT12), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT12), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n484_), .A2(new_n499_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n458_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n457_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  XOR2_X1   g307(.A(G176gat), .B(G204gat), .Z(new_n509_));
  XNOR2_X1  g308(.A(G120gat), .B(G148gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n506_), .A2(new_n508_), .A3(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n513_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n516_));
  AND2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n517_), .A2(KEYINPUT13), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(KEYINPUT13), .A3(new_n516_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(G1gat), .B(G8gat), .Z(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT74), .ZN(new_n525_));
  INV_X1    g324(.A(G1gat), .ZN(new_n526_));
  INV_X1    g325(.A(G8gat), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT14), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n524_), .A2(new_n525_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n525_), .B1(new_n524_), .B2(new_n528_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n523_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n531_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(new_n522_), .A3(new_n529_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(G29gat), .ZN(new_n536_));
  INV_X1    g335(.A(G36gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G29gat), .A2(G36gat), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(G50gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(G50gat), .A3(new_n539_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT68), .B(G43gat), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n544_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n535_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n547_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT15), .B1(new_n551_), .B2(new_n545_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553_));
  NOR3_X1   g352(.A1(new_n546_), .A2(new_n547_), .A3(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n549_), .B(new_n550_), .C1(new_n555_), .C2(new_n535_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n550_), .ZN(new_n557_));
  AOI211_X1 g356(.A(new_n547_), .B(new_n546_), .C1(new_n532_), .C2(new_n534_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n535_), .A2(new_n548_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AND3_X1   g363(.A1(new_n556_), .A2(new_n560_), .A3(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n564_), .B1(new_n556_), .B2(new_n560_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n521_), .A2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(KEYINPUT69), .B(KEYINPUT70), .Z(new_n569_));
  XNOR2_X1  g368(.A(G190gat), .B(G218gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G134gat), .B(G162gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT36), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT71), .Z(new_n576_));
  OR2_X1    g375(.A1(new_n576_), .A2(KEYINPUT72), .ZN(new_n577_));
  INV_X1    g376(.A(new_n484_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n548_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G232gat), .A2(G233gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT34), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT67), .B(KEYINPUT35), .ZN(new_n582_));
  OAI221_X1 g381(.A(new_n579_), .B1(new_n581_), .B2(new_n582_), .C1(new_n578_), .C2(new_n555_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n582_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n583_), .A2(new_n585_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n576_), .A2(KEYINPUT72), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n577_), .A2(new_n586_), .A3(new_n587_), .A4(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n586_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n573_), .A2(new_n574_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n575_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT73), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(KEYINPUT37), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT37), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n589_), .B(new_n592_), .C1(new_n594_), .C2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n498_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(new_n535_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(G211gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(KEYINPUT16), .B(G183gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(KEYINPUT17), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n603_), .A2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n607_), .A2(KEYINPUT17), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n610_), .B1(new_n603_), .B2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n600_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n456_), .A2(new_n568_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT98), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n526_), .A3(new_n443_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT38), .ZN(new_n620_));
  NOR3_X1   g419(.A1(new_n521_), .A2(new_n567_), .A3(new_n614_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n450_), .A2(new_n452_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n454_), .A2(new_n453_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n401_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n415_), .A2(new_n417_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n622_), .B(new_n593_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n622_), .B1(new_n456_), .B2(new_n593_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n621_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n443_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G1gat), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n620_), .A2(new_n632_), .ZN(G1324gat));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n301_), .A2(new_n413_), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n635_), .B(new_n621_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n636_), .A2(new_n637_), .A3(G8gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n637_), .B1(new_n636_), .B2(G8gat), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n634_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(G8gat), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT101), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n636_), .A2(new_n637_), .A3(G8gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(KEYINPUT39), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n616_), .B(KEYINPUT98), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n635_), .A2(new_n527_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n645_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n618_), .A2(KEYINPUT100), .A3(new_n527_), .A4(new_n635_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n640_), .A2(new_n644_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT40), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n640_), .A2(new_n644_), .A3(KEYINPUT40), .A4(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1325gat));
  AND2_X1   g454(.A1(new_n456_), .A2(new_n568_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n656_), .A2(new_n378_), .A3(new_n401_), .A4(new_n615_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n401_), .B(new_n621_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n658_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT41), .B1(new_n658_), .B2(G15gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n657_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT102), .Z(G1326gat));
  XNOR2_X1  g461(.A(new_n451_), .B(KEYINPUT103), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n630_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n664_), .A2(new_n665_), .A3(G22gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n664_), .B2(G22gat), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n663_), .A2(G22gat), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT104), .ZN(new_n669_));
  OAI22_X1  g468(.A1(new_n666_), .A2(new_n667_), .B1(new_n616_), .B2(new_n669_), .ZN(G1327gat));
  OAI21_X1  g469(.A(new_n600_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT43), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n673_), .B(new_n600_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n568_), .A3(new_n614_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n675_), .A2(KEYINPUT44), .A3(new_n568_), .A4(new_n614_), .ZN(new_n679_));
  AND3_X1   g478(.A1(new_n678_), .A2(new_n443_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n614_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n593_), .A2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n656_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n443_), .A2(new_n536_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT105), .ZN(new_n685_));
  OAI22_X1  g484(.A1(new_n680_), .A2(new_n536_), .B1(new_n683_), .B2(new_n685_), .ZN(G1328gat));
  NAND3_X1  g485(.A1(new_n678_), .A2(new_n635_), .A3(new_n679_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(G36gat), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n656_), .A2(new_n537_), .A3(new_n635_), .A4(new_n682_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT45), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT46), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n688_), .A2(KEYINPUT46), .A3(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1329gat));
  NAND4_X1  g494(.A1(new_n678_), .A2(G43gat), .A3(new_n401_), .A4(new_n679_), .ZN(new_n696_));
  INV_X1    g495(.A(G43gat), .ZN(new_n697_));
  INV_X1    g496(.A(new_n401_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n683_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g500(.A1(new_n678_), .A2(G50gat), .A3(new_n451_), .A4(new_n679_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n541_), .B1(new_n683_), .B2(new_n663_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1331gat));
  INV_X1    g503(.A(new_n456_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n556_), .A2(new_n560_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n563_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n556_), .A2(new_n560_), .A3(new_n564_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT106), .B1(new_n705_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT106), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n456_), .A2(new_n711_), .A3(new_n567_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n710_), .A2(new_n521_), .A3(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n615_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n714_), .A2(new_n631_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(G57gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n614_), .A2(new_n709_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n521_), .A2(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n593_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT99), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n718_), .B1(new_n720_), .B2(new_n627_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(KEYINPUT107), .B(G57gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n443_), .A3(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n723_), .A2(KEYINPUT108), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(KEYINPUT108), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n716_), .A2(new_n724_), .A3(new_n725_), .ZN(G1332gat));
  NAND2_X1  g525(.A1(new_n721_), .A2(new_n635_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(new_n728_), .A3(G64gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G64gat), .ZN(new_n730_));
  INV_X1    g529(.A(new_n635_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n731_), .A2(G64gat), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT109), .Z(new_n733_));
  OAI22_X1  g532(.A1(new_n729_), .A2(new_n730_), .B1(new_n714_), .B2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT110), .ZN(G1333gat));
  INV_X1    g534(.A(KEYINPUT49), .ZN(new_n736_));
  INV_X1    g535(.A(new_n718_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n401_), .B(new_n737_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(G71gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G71gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n736_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(G71gat), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT111), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n738_), .A2(new_n739_), .A3(G71gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(KEYINPUT49), .A3(new_n745_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n698_), .A2(G71gat), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT112), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n713_), .A2(new_n615_), .A3(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n742_), .A2(new_n746_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT113), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n742_), .A2(new_n746_), .A3(new_n752_), .A4(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1334gat));
  INV_X1    g553(.A(new_n663_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n721_), .A2(new_n755_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(G78gat), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G78gat), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n755_), .A2(new_n491_), .ZN(new_n760_));
  OAI22_X1  g559(.A1(new_n758_), .A2(new_n759_), .B1(new_n714_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n761_), .B(new_n762_), .ZN(G1335gat));
  NOR2_X1   g562(.A1(new_n681_), .A2(new_n709_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n674_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n673_), .B1(new_n456_), .B2(new_n600_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n521_), .B(new_n764_), .C1(new_n765_), .C2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT116), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n675_), .A2(KEYINPUT116), .A3(new_n521_), .A4(new_n764_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n443_), .A2(G85gat), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT117), .Z(new_n772_));
  NAND3_X1  g571(.A1(new_n769_), .A2(new_n770_), .A3(new_n772_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n710_), .A2(new_n521_), .A3(new_n682_), .A4(new_n712_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n462_), .B1(new_n774_), .B2(new_n631_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1336gat));
  NAND4_X1  g575(.A1(new_n769_), .A2(G92gat), .A3(new_n770_), .A4(new_n635_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n275_), .B1(new_n774_), .B2(new_n731_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1337gat));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n780_), .A2(KEYINPUT51), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n769_), .A2(new_n401_), .A3(new_n770_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(G99gat), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(KEYINPUT51), .ZN(new_n784_));
  NOR3_X1   g583(.A1(new_n774_), .A2(new_n470_), .A3(new_n698_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AND4_X1   g585(.A1(new_n781_), .A2(new_n783_), .A3(new_n784_), .A4(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n785_), .B1(new_n782_), .B2(G99gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n781_), .B1(new_n788_), .B2(new_n784_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1338gat));
  NAND4_X1  g589(.A1(new_n675_), .A2(new_n451_), .A3(new_n521_), .A4(new_n764_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n791_), .A2(new_n792_), .A3(G106gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n791_), .B2(G106gat), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n451_), .A2(new_n477_), .ZN(new_n795_));
  OAI22_X1  g594(.A1(new_n793_), .A2(new_n794_), .B1(new_n774_), .B2(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g596(.A(KEYINPUT56), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n505_), .A2(KEYINPUT55), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n800_), .B(new_n458_), .C1(new_n502_), .C2(new_n504_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n502_), .A2(new_n458_), .A3(new_n504_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n799_), .A2(new_n801_), .A3(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n798_), .B1(new_n804_), .B2(new_n514_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n506_), .A2(new_n800_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n505_), .A2(KEYINPUT55), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n802_), .A3(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(KEYINPUT56), .A3(new_n513_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT120), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n805_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT120), .B(new_n798_), .C1(new_n804_), .C2(new_n514_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n557_), .B(new_n549_), .C1(new_n555_), .C2(new_n535_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n550_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n563_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n708_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n812_), .A2(new_n817_), .A3(new_n515_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT58), .B1(new_n811_), .B2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT56), .B1(new_n808_), .B2(new_n513_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n816_), .B1(new_n820_), .B2(KEYINPUT120), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n805_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .A4(new_n515_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n819_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n600_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT121), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n505_), .A2(new_n507_), .A3(new_n513_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n567_), .B2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n709_), .A2(new_n515_), .A3(KEYINPUT119), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(new_n805_), .B2(new_n809_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n517_), .A2(new_n816_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n593_), .B(new_n828_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n827_), .A2(KEYINPUT121), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n593_), .B(new_n837_), .C1(new_n834_), .C2(new_n835_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n826_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n614_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n599_), .A2(new_n520_), .A3(new_n717_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(KEYINPUT54), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n451_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n635_), .A2(new_n631_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n401_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G113gat), .B1(new_n848_), .B2(new_n709_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT122), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(KEYINPUT59), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n825_), .A2(new_n600_), .B1(new_n836_), .B2(new_n838_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n681_), .B1(new_n852_), .B2(new_n840_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT54), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n843_), .B(new_n854_), .ZN(new_n855_));
  OAI211_X1 g654(.A(new_n452_), .B(new_n846_), .C1(new_n853_), .C2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n851_), .B1(new_n856_), .B2(new_n698_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n845_), .A2(new_n401_), .A3(new_n846_), .A4(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT123), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n857_), .A2(new_n859_), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n862_), .A2(new_n567_), .A3(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n849_), .B1(new_n866_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g666(.A(G120gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n520_), .B2(KEYINPUT60), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n848_), .B(new_n869_), .C1(KEYINPUT60), .C2(new_n868_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n520_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n868_), .B2(new_n871_), .ZN(G1341gat));
  AOI21_X1  g671(.A(G127gat), .B1(new_n848_), .B2(new_n681_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n862_), .A2(new_n865_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n681_), .A2(G127gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(G1342gat));
  NAND4_X1  g675(.A1(new_n861_), .A2(G134gat), .A3(new_n600_), .A4(new_n864_), .ZN(new_n877_));
  INV_X1    g676(.A(G134gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n847_), .B2(new_n593_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT124), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n877_), .A2(new_n879_), .A3(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(G1343gat));
  NOR2_X1   g683(.A1(new_n853_), .A2(new_n855_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n401_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n886_), .A2(new_n451_), .A3(new_n846_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n567_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(new_n318_), .ZN(G1344gat));
  NOR2_X1   g688(.A1(new_n887_), .A2(new_n520_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(new_n319_), .ZN(G1345gat));
  NOR2_X1   g690(.A1(new_n887_), .A2(new_n614_), .ZN(new_n892_));
  XOR2_X1   g691(.A(KEYINPUT61), .B(G155gat), .Z(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1346gat));
  INV_X1    g693(.A(G162gat), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n887_), .A2(new_n895_), .A3(new_n599_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n887_), .A2(new_n593_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n895_), .B2(new_n897_), .ZN(G1347gat));
  NAND2_X1  g697(.A1(new_n635_), .A2(new_n407_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n885_), .A2(new_n755_), .A3(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n709_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n900_), .A2(KEYINPUT125), .A3(new_n709_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(G169gat), .A3(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n906_), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n907_), .B(new_n908_), .C1(new_n225_), .C2(new_n901_), .ZN(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n900_), .B2(new_n521_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n521_), .A2(G176gat), .ZN(new_n911_));
  INV_X1    g710(.A(new_n845_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n899_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n910_), .B1(new_n911_), .B2(new_n913_), .ZN(G1349gat));
  NAND3_X1  g713(.A1(new_n635_), .A2(new_n407_), .A3(new_n681_), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n912_), .A2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n885_), .A2(new_n755_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n915_), .A2(new_n229_), .ZN(new_n918_));
  AOI22_X1  g717(.A1(new_n916_), .A2(new_n219_), .B1(new_n917_), .B2(new_n918_), .ZN(G1350gat));
  INV_X1    g718(.A(new_n900_), .ZN(new_n920_));
  OAI21_X1  g719(.A(G190gat), .B1(new_n920_), .B2(new_n599_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n589_), .A2(new_n592_), .A3(new_n228_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n920_), .B2(new_n922_), .ZN(G1351gat));
  NAND3_X1  g722(.A1(new_n886_), .A2(new_n453_), .A3(new_n635_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n567_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n213_), .ZN(G1352gat));
  AND3_X1   g725(.A1(new_n886_), .A2(new_n453_), .A3(new_n635_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n521_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(G204gat), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n929_), .B1(new_n212_), .B2(new_n928_), .ZN(G1353gat));
  NAND2_X1  g729(.A1(new_n927_), .A2(new_n681_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  AND2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n931_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n934_), .B1(new_n931_), .B2(new_n932_), .ZN(G1354gat));
  NAND3_X1  g734(.A1(new_n927_), .A2(G218gat), .A3(new_n600_), .ZN(new_n936_));
  INV_X1    g735(.A(G218gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n937_), .B1(new_n924_), .B2(new_n593_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n936_), .A2(new_n938_), .ZN(new_n939_));
  XOR2_X1   g738(.A(new_n939_), .B(KEYINPUT127), .Z(G1355gat));
endmodule


