//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 0 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n617_,
    new_n618_, new_n619_, new_n621_, new_n622_, new_n623_, new_n624_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n843_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n871_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT97), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT19), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT23), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT83), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT84), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n207_), .A2(KEYINPUT83), .A3(KEYINPUT23), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n211_), .A2(KEYINPUT84), .A3(G183gat), .A4(G190gat), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n210_), .A2(new_n214_), .A3(new_n215_), .A4(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n206_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT22), .B(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G169gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(new_n221_), .ZN(new_n225_));
  OR2_X1    g024(.A1(new_n225_), .A2(KEYINPUT24), .ZN(new_n226_));
  NOR2_X1   g025(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n227_));
  AND2_X1   g026(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n228_));
  AND2_X1   g027(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n230_));
  OAI22_X1  g029(.A1(new_n227_), .A2(new_n228_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n225_), .A2(KEYINPUT24), .A3(new_n205_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n208_), .A2(new_n212_), .ZN(new_n233_));
  AND4_X1   g032(.A1(new_n226_), .A2(new_n231_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n223_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT103), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G197gat), .B(G204gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT21), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT95), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G211gat), .B(G218gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n241_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G197gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(G204gat), .ZN(new_n247_));
  INV_X1    g046(.A(G204gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n248_), .A2(G197gat), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n242_), .B(KEYINPUT21), .C1(new_n247_), .C2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n239_), .A2(new_n240_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(new_n243_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n245_), .A2(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n234_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT103), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n238_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n253_), .A2(KEYINPUT96), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n226_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(new_n217_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT86), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT22), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n260_), .B(G169gat), .C1(new_n261_), .C2(KEYINPUT85), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT85), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n263_), .B(KEYINPUT22), .C1(new_n224_), .C2(KEYINPUT86), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT85), .B1(new_n261_), .B2(G169gat), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n262_), .A2(new_n264_), .A3(new_n221_), .A4(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n233_), .A2(new_n218_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n267_), .A3(new_n205_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n259_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n245_), .A2(new_n252_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT96), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n257_), .A2(new_n269_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT20), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n204_), .B1(new_n256_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT104), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n269_), .B1(new_n257_), .B2(new_n272_), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT20), .B1(new_n254_), .B2(new_n253_), .ZN(new_n278_));
  OR3_X1    g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n204_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT104), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n280_), .B(new_n204_), .C1(new_n256_), .C2(new_n274_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n276_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G8gat), .B(G36gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G64gat), .B(G92gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n285_), .B(new_n286_), .Z(new_n287_));
  NAND2_X1  g086(.A1(new_n282_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT106), .ZN(new_n289_));
  INV_X1    g088(.A(new_n287_), .ZN(new_n290_));
  AND4_X1   g089(.A1(KEYINPUT98), .A2(new_n223_), .A3(new_n253_), .A4(new_n235_), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT98), .B1(new_n254_), .B2(new_n253_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT20), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n270_), .B(KEYINPUT96), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n295_), .B2(new_n269_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n204_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n204_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n277_), .A2(new_n278_), .A3(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n290_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT106), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n282_), .A2(new_n301_), .A3(new_n287_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n289_), .A2(new_n300_), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT27), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT98), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n305_), .B1(new_n236_), .B2(new_n270_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n254_), .A2(KEYINPUT98), .A3(new_n253_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n298_), .B1(new_n308_), .B2(new_n274_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n299_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(new_n287_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n300_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT27), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n304_), .A2(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G78gat), .B(G106gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT92), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT28), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT88), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n321_), .B1(G155gat), .B2(G162gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G155gat), .A2(G162gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n323_), .A2(KEYINPUT88), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT1), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G155gat), .ZN(new_n326_));
  INV_X1    g125(.A(G162gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n323_), .A2(KEYINPUT88), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n321_), .A2(G155gat), .A3(G162gat), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT1), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n325_), .A2(new_n328_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT89), .ZN(new_n334_));
  XOR2_X1   g133(.A(G141gat), .B(G148gat), .Z(new_n335_));
  AND3_X1   g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n334_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT91), .ZN(new_n338_));
  AND2_X1   g137(.A1(KEYINPUT90), .A2(KEYINPUT3), .ZN(new_n339_));
  NOR2_X1   g138(.A1(KEYINPUT90), .A2(KEYINPUT3), .ZN(new_n340_));
  OAI22_X1  g139(.A1(new_n339_), .A2(new_n340_), .B1(G141gat), .B2(G148gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(KEYINPUT90), .A2(KEYINPUT3), .ZN(new_n342_));
  INV_X1    g141(.A(G141gat), .ZN(new_n343_));
  INV_X1    g142(.A(G148gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT2), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n341_), .A2(new_n345_), .A3(new_n347_), .A4(new_n348_), .ZN(new_n349_));
  AOI22_X1  g148(.A1(new_n329_), .A2(new_n330_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n338_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n349_), .A2(new_n338_), .A3(new_n350_), .ZN(new_n352_));
  OAI22_X1  g151(.A1(new_n336_), .A2(new_n337_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n353_), .A2(KEYINPUT29), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G22gat), .B(G50gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n353_), .A2(KEYINPUT29), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n295_), .ZN(new_n358_));
  AND2_X1   g157(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(G233gat), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n361_), .B(KEYINPUT94), .Z(new_n362_));
  NAND2_X1  g161(.A1(new_n358_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n362_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n357_), .A2(new_n270_), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n356_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n356_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n320_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n354_), .B(new_n355_), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n365_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n372_), .A2(new_n366_), .A3(new_n319_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n369_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G127gat), .B(G134gat), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n375_), .A2(G113gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(G113gat), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n376_), .A2(G120gat), .A3(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(G120gat), .B1(new_n376_), .B2(new_n377_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n353_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n349_), .A2(new_n350_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT91), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n349_), .A2(new_n338_), .A3(new_n350_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n386_), .B(new_n380_), .C1(new_n337_), .C2(new_n336_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n382_), .A2(KEYINPUT100), .A3(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n336_), .A2(new_n337_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT100), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n389_), .A2(new_n390_), .A3(new_n386_), .A4(new_n380_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(KEYINPUT4), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393_));
  XOR2_X1   g192(.A(new_n393_), .B(KEYINPUT101), .Z(new_n394_));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n382_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n392_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n394_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n388_), .A2(new_n398_), .A3(new_n391_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT0), .B(G57gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(G85gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(G1gat), .B(G29gat), .Z(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n400_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n397_), .A2(new_n404_), .A3(new_n399_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT87), .B(KEYINPUT30), .ZN(new_n410_));
  XOR2_X1   g209(.A(new_n380_), .B(new_n410_), .Z(new_n411_));
  XNOR2_X1  g210(.A(G71gat), .B(G99gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G15gat), .B(G43gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT31), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G227gat), .A2(G233gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n415_), .B(new_n416_), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(new_n269_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n413_), .B(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n409_), .A2(new_n419_), .ZN(new_n420_));
  NOR3_X1   g219(.A1(new_n316_), .A2(new_n374_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT33), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n406_), .A2(KEYINPUT102), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT102), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n404_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n424_), .B1(new_n425_), .B2(KEYINPUT33), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(KEYINPUT33), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n392_), .A2(new_n396_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n405_), .B1(new_n428_), .B2(new_n398_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n388_), .A2(new_n391_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n394_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n312_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n423_), .A2(new_n426_), .A3(new_n427_), .A4(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n282_), .A2(KEYINPUT32), .A3(new_n290_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n290_), .A2(KEYINPUT32), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n408_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n433_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n374_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT105), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n304_), .A2(new_n315_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n374_), .A2(new_n409_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n438_), .A2(KEYINPUT105), .A3(new_n439_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n442_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n419_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n421_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(G120gat), .B(G148gat), .Z(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G176gat), .B(G204gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n458_), .A2(KEYINPUT73), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT77), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT69), .B(G71gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(G78gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G57gat), .B(G64gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(KEYINPUT11), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n463_), .B(KEYINPUT11), .Z(new_n466_));
  OAI21_X1  g265(.A(new_n465_), .B1(new_n462_), .B2(new_n466_), .ZN(new_n467_));
  XOR2_X1   g266(.A(KEYINPUT70), .B(KEYINPUT71), .Z(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n467_), .B(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT65), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n471_), .B1(G85gat), .B2(G92gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT9), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n473_), .B1(G85gat), .B2(G92gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT6), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G106gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(KEYINPUT10), .B(G99gat), .Z(new_n479_));
  AOI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n474_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT8), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(G99gat), .A2(G106gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT7), .ZN(new_n486_));
  INV_X1    g285(.A(new_n483_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n476_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n484_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G85gat), .B(G92gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT66), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n482_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n482_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n493_), .B1(new_n486_), .B2(new_n476_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n481_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT12), .B1(new_n470_), .B2(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n470_), .A2(new_n495_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G230gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT64), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n481_), .A2(KEYINPUT72), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT72), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n503_), .B1(new_n474_), .B2(new_n480_), .ZN(new_n504_));
  OAI22_X1  g303(.A1(new_n502_), .A2(new_n504_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n470_), .A2(new_n505_), .A3(KEYINPUT12), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n498_), .A2(new_n501_), .A3(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n470_), .A2(new_n495_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n500_), .B1(new_n508_), .B2(new_n497_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n460_), .B(new_n510_), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n511_), .A2(KEYINPUT13), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(KEYINPUT13), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G29gat), .B(G36gat), .ZN(new_n516_));
  INV_X1    g315(.A(G43gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(G50gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT15), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G15gat), .B(G22gat), .ZN(new_n522_));
  INV_X1    g321(.A(G1gat), .ZN(new_n523_));
  INV_X1    g322(.A(G8gat), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT14), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G1gat), .B(G8gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n521_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT82), .Z(new_n531_));
  INV_X1    g330(.A(new_n520_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n529_), .B(new_n531_), .C1(new_n528_), .C2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n520_), .B(new_n528_), .Z(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(G229gat), .A3(G233gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G113gat), .B(G141gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n224_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(new_n246_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n533_), .A2(new_n535_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n515_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n450_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT34), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT35), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n521_), .A2(new_n505_), .ZN(new_n551_));
  AOI211_X1 g350(.A(new_n549_), .B(new_n548_), .C1(new_n551_), .C2(KEYINPUT78), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n532_), .B2(new_n495_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n552_), .A2(new_n553_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n550_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT79), .B(G190gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(G218gat), .ZN(new_n559_));
  XOR2_X1   g358(.A(G134gat), .B(G162gat), .Z(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n556_), .A2(new_n557_), .A3(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n552_), .B(new_n553_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n557_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n561_), .A2(new_n557_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n563_), .A2(new_n564_), .A3(new_n565_), .A4(new_n550_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n567_), .B(KEYINPUT37), .Z(new_n568_));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n528_), .B(new_n569_), .Z(new_n570_));
  XNOR2_X1  g369(.A(new_n470_), .B(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G183gat), .B(G211gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(G155gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT81), .B(G127gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n575_), .B(new_n576_), .Z(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT17), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n571_), .A2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n577_), .B(KEYINPUT17), .Z(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(new_n580_), .B2(new_n571_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n568_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n545_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT107), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n545_), .A2(KEYINPUT107), .A3(new_n583_), .ZN(new_n587_));
  AOI21_X1  g386(.A(G1gat), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n408_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT108), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT108), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n588_), .A2(new_n591_), .A3(new_n408_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT38), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n567_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(new_n582_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n545_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(G1gat), .B1(new_n598_), .B2(new_n409_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n590_), .A2(KEYINPUT38), .A3(new_n592_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n595_), .A2(new_n599_), .A3(new_n600_), .ZN(G1324gat));
  INV_X1    g400(.A(KEYINPUT109), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n598_), .B2(new_n443_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n545_), .A2(KEYINPUT109), .A3(new_n597_), .A4(new_n316_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(G8gat), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT39), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n603_), .A2(new_n607_), .A3(G8gat), .A4(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n586_), .A2(new_n587_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n524_), .A3(new_n316_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT40), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n609_), .A2(KEYINPUT40), .A3(new_n611_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1325gat));
  OAI21_X1  g415(.A(G15gat), .B1(new_n598_), .B2(new_n449_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT41), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n584_), .A2(G15gat), .A3(new_n449_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(G1326gat));
  XOR2_X1   g419(.A(new_n374_), .B(KEYINPUT110), .Z(new_n621_));
  OAI21_X1  g420(.A(G22gat), .B1(new_n598_), .B2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT42), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n621_), .A2(G22gat), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n623_), .B1(new_n584_), .B2(new_n624_), .ZN(G1327gat));
  NAND3_X1  g424(.A1(new_n515_), .A2(new_n582_), .A3(new_n543_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n450_), .A2(new_n567_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(G29gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n628_), .A3(new_n408_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n568_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT43), .B1(new_n450_), .B2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n316_), .A2(new_n374_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n420_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT105), .B1(new_n438_), .B2(new_n439_), .ZN(new_n635_));
  AOI211_X1 g434(.A(new_n441_), .B(new_n374_), .C1(new_n433_), .C2(new_n437_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n444_), .B1(new_n304_), .B2(new_n315_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n634_), .B1(new_n638_), .B2(new_n419_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(new_n640_), .A3(new_n568_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n631_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n626_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT111), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(KEYINPUT44), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n642_), .A2(new_n643_), .A3(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n646_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n648_), .A2(new_n409_), .A3(new_n649_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n629_), .B1(new_n650_), .B2(new_n628_), .ZN(G1328gat));
  NOR3_X1   g450(.A1(new_n450_), .A2(KEYINPUT43), .A3(new_n630_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n640_), .B1(new_n639_), .B2(new_n568_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n643_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n645_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n316_), .A3(new_n647_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(G36gat), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT113), .ZN(new_n658_));
  INV_X1    g457(.A(G36gat), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n443_), .A2(KEYINPUT112), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n443_), .A2(KEYINPUT112), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n627_), .A2(new_n658_), .A3(new_n659_), .A4(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n639_), .A2(new_n659_), .A3(new_n596_), .A4(new_n643_), .ZN(new_n665_));
  OAI21_X1  g464(.A(KEYINPUT113), .B1(new_n665_), .B2(new_n662_), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n664_), .A2(new_n666_), .A3(KEYINPUT45), .ZN(new_n667_));
  AOI21_X1  g466(.A(KEYINPUT45), .B1(new_n664_), .B2(new_n666_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n657_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT114), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT46), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT46), .ZN(new_n673_));
  AOI211_X1 g472(.A(KEYINPUT114), .B(new_n673_), .C1(new_n657_), .C2(new_n669_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n672_), .A2(new_n674_), .ZN(G1329gat));
  NAND4_X1  g474(.A1(new_n655_), .A2(G43gat), .A3(new_n419_), .A4(new_n647_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n627_), .A2(new_n419_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(KEYINPUT115), .A2(G43gat), .ZN(new_n678_));
  OR2_X1    g477(.A1(KEYINPUT115), .A2(G43gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n676_), .A2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g481(.A(new_n621_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n627_), .A2(new_n519_), .A3(new_n683_), .ZN(new_n684_));
  NOR3_X1   g483(.A1(new_n648_), .A2(new_n439_), .A3(new_n649_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(new_n519_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT116), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1331gat));
  INV_X1    g487(.A(G57gat), .ZN(new_n689_));
  INV_X1    g488(.A(new_n543_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n514_), .A2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n450_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n583_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n689_), .B1(new_n693_), .B2(new_n409_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT117), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n692_), .A2(new_n597_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n409_), .A2(new_n689_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n695_), .B1(new_n696_), .B2(new_n697_), .ZN(G1332gat));
  INV_X1    g497(.A(G64gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n696_), .B2(new_n663_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT48), .Z(new_n701_));
  INV_X1    g500(.A(new_n693_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n699_), .A3(new_n663_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1333gat));
  INV_X1    g503(.A(new_n696_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G71gat), .B1(new_n705_), .B2(new_n449_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT118), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT49), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n706_), .A2(KEYINPUT118), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n706_), .A2(KEYINPUT118), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(KEYINPUT49), .A3(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n702_), .A2(new_n419_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n709_), .B(new_n712_), .C1(G71gat), .C2(new_n713_), .ZN(G1334gat));
  INV_X1    g513(.A(G78gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n696_), .B2(new_n683_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT50), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n702_), .A2(new_n715_), .A3(new_n683_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1335gat));
  NAND3_X1  g518(.A1(new_n514_), .A2(new_n582_), .A3(new_n690_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n639_), .A2(new_n596_), .A3(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(G85gat), .B1(new_n723_), .B2(new_n408_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n720_), .B1(new_n631_), .B2(new_n641_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n725_), .A2(new_n408_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n726_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g526(.A(G92gat), .B1(new_n723_), .B2(new_n316_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n663_), .A2(G92gat), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n725_), .B2(new_n729_), .ZN(G1337gat));
  NAND2_X1  g529(.A1(new_n725_), .A2(new_n419_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n419_), .A2(new_n479_), .ZN(new_n732_));
  AOI22_X1  g531(.A1(new_n731_), .A2(G99gat), .B1(new_n723_), .B2(new_n732_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g533(.A(KEYINPUT52), .ZN(new_n735_));
  AOI211_X1 g534(.A(KEYINPUT119), .B(new_n478_), .C1(new_n725_), .C2(new_n374_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT119), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n642_), .A2(new_n374_), .A3(new_n721_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(G106gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n736_), .B2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n723_), .A2(new_n478_), .A3(new_n374_), .ZN(new_n741_));
  AOI211_X1 g540(.A(new_n439_), .B(new_n720_), .C1(new_n631_), .C2(new_n641_), .ZN(new_n742_));
  OAI21_X1  g541(.A(KEYINPUT119), .B1(new_n742_), .B2(new_n478_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n738_), .A2(new_n737_), .A3(G106gat), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(KEYINPUT52), .A3(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n740_), .A2(new_n741_), .A3(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT53), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT53), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n740_), .A2(new_n745_), .A3(new_n748_), .A4(new_n741_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1339gat));
  AOI21_X1  g549(.A(new_n501_), .B1(new_n498_), .B2(new_n506_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT55), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n507_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n498_), .A2(KEYINPUT55), .A3(new_n501_), .A4(new_n506_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n457_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT56), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n507_), .A2(new_n509_), .A3(new_n458_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n458_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT56), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n757_), .A2(new_n543_), .A3(new_n758_), .A4(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n511_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n534_), .A2(new_n531_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n529_), .B1(new_n528_), .B2(new_n532_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n539_), .B(new_n764_), .C1(new_n765_), .C2(new_n531_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n542_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT120), .Z(new_n768_));
  NAND2_X1  g567(.A1(new_n763_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n762_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT57), .B1(new_n770_), .B2(new_n567_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT57), .ZN(new_n772_));
  AOI211_X1 g571(.A(new_n772_), .B(new_n596_), .C1(new_n762_), .C2(new_n769_), .ZN(new_n773_));
  OAI21_X1  g572(.A(KEYINPUT121), .B1(new_n771_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT121), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n596_), .B1(new_n762_), .B2(new_n769_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(KEYINPUT57), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n774_), .A2(new_n777_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n757_), .A2(new_n768_), .A3(new_n758_), .A4(new_n761_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT122), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n568_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT123), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n779_), .A2(new_n783_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT123), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n568_), .B(new_n788_), .C1(new_n782_), .C2(new_n784_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n786_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n581_), .B1(new_n778_), .B2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n583_), .A2(new_n690_), .A3(new_n515_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT54), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n791_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n632_), .A2(new_n408_), .A3(new_n419_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(G113gat), .B1(new_n797_), .B2(new_n543_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n792_), .B(KEYINPUT54), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n771_), .A2(new_n773_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n790_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n799_), .B1(new_n801_), .B2(new_n581_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT59), .ZN(new_n803_));
  INV_X1    g602(.A(new_n796_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n802_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n797_), .B2(new_n803_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n806_), .A2(new_n690_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n798_), .B1(new_n807_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g607(.A(G120gat), .B1(new_n806_), .B2(new_n515_), .ZN(new_n809_));
  INV_X1    g608(.A(G120gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n515_), .B2(KEYINPUT60), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT124), .B1(new_n810_), .B2(KEYINPUT60), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT124), .ZN(new_n814_));
  OAI211_X1 g613(.A(new_n797_), .B(new_n813_), .C1(new_n814_), .C2(new_n811_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n809_), .A2(new_n815_), .ZN(G1341gat));
  AOI21_X1  g615(.A(G127gat), .B1(new_n797_), .B2(new_n581_), .ZN(new_n817_));
  INV_X1    g616(.A(G127gat), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n806_), .A2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n817_), .B1(new_n819_), .B2(new_n581_), .ZN(G1342gat));
  INV_X1    g619(.A(G134gat), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n774_), .A2(new_n777_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n789_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n759_), .B(KEYINPUT56), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n824_), .A2(KEYINPUT122), .A3(new_n768_), .A4(new_n758_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(new_n781_), .A3(new_n783_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n788_), .B1(new_n826_), .B2(new_n568_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n823_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n822_), .B1(new_n828_), .B2(new_n787_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n799_), .B1(new_n829_), .B2(new_n581_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n804_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n821_), .B1(new_n831_), .B2(new_n567_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT125), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT125), .B(new_n821_), .C1(new_n831_), .C2(new_n567_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n630_), .A2(new_n821_), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n805_), .B(new_n836_), .C1(new_n797_), .C2(new_n803_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n834_), .A2(new_n835_), .A3(new_n837_), .ZN(G1343gat));
  NOR2_X1   g637(.A1(new_n439_), .A2(new_n409_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n830_), .A2(new_n449_), .A3(new_n662_), .A4(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n690_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(new_n343_), .ZN(G1344gat));
  NOR2_X1   g641(.A1(new_n840_), .A2(new_n515_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n843_), .B(new_n344_), .ZN(G1345gat));
  NOR2_X1   g643(.A1(new_n840_), .A2(new_n582_), .ZN(new_n845_));
  XOR2_X1   g644(.A(KEYINPUT61), .B(G155gat), .Z(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(G1346gat));
  NOR3_X1   g646(.A1(new_n840_), .A2(new_n327_), .A3(new_n630_), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n840_), .A2(new_n567_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n327_), .B2(new_n849_), .ZN(G1347gat));
  NAND2_X1  g649(.A1(new_n663_), .A2(new_n633_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n683_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n802_), .A2(new_n543_), .A3(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT126), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT62), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n853_), .A2(G169gat), .A3(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n854_), .A2(KEYINPUT62), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n802_), .A2(new_n852_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n859_), .A2(new_n220_), .A3(new_n543_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n857_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n853_), .A2(G169gat), .A3(new_n861_), .A4(new_n855_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n858_), .A2(new_n860_), .A3(new_n862_), .ZN(G1348gat));
  AOI21_X1  g662(.A(G176gat), .B1(new_n859_), .B2(new_n514_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n795_), .A2(new_n374_), .A3(new_n851_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n515_), .A2(new_n221_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(G1349gat));
  AOI21_X1  g666(.A(G183gat), .B1(new_n865_), .B2(new_n581_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n582_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n859_), .B2(new_n869_), .ZN(G1350gat));
  NAND2_X1  g669(.A1(new_n859_), .A2(new_n568_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G190gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n859_), .B1(new_n230_), .B2(new_n229_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n567_), .B2(new_n873_), .ZN(G1351gat));
  OAI211_X1 g673(.A(new_n449_), .B(new_n445_), .C1(new_n791_), .C2(new_n794_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n662_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n543_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n514_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g679(.A1(new_n830_), .A2(new_n449_), .A3(new_n445_), .A4(new_n663_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT127), .ZN(new_n882_));
  XOR2_X1   g681(.A(KEYINPUT63), .B(G211gat), .Z(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NOR4_X1   g683(.A1(new_n881_), .A2(new_n882_), .A3(new_n582_), .A4(new_n884_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n875_), .A2(new_n582_), .A3(new_n662_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n883_), .ZN(new_n887_));
  OR2_X1    g686(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(KEYINPUT127), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n885_), .B1(new_n887_), .B2(new_n889_), .ZN(G1354gat));
  AOI21_X1  g689(.A(G218gat), .B1(new_n876_), .B2(new_n596_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n881_), .A2(new_n630_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(G218gat), .B2(new_n892_), .ZN(G1355gat));
endmodule


