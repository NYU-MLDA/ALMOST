//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207_));
  INV_X1    g006(.A(G1gat), .ZN(new_n208_));
  INV_X1    g007(.A(G8gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G1gat), .B(G8gat), .ZN(new_n212_));
  XOR2_X1   g011(.A(new_n211_), .B(new_n212_), .Z(new_n213_));
  OR2_X1    g012(.A1(G29gat), .A2(G36gat), .ZN(new_n214_));
  INV_X1    g013(.A(G43gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G29gat), .A2(G36gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G50gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n215_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n214_), .A2(new_n216_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G43gat), .ZN(new_n223_));
  AOI21_X1  g022(.A(G50gat), .B1(new_n223_), .B2(new_n217_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT77), .B1(new_n221_), .B2(new_n224_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n219_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT77), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n223_), .A2(G50gat), .A3(new_n217_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT15), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n225_), .A2(KEYINPUT15), .A3(new_n229_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n213_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n221_), .A2(new_n224_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n213_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NOR3_X1   g038(.A1(new_n234_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n213_), .A2(new_n237_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(new_n235_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n206_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT82), .ZN(new_n245_));
  INV_X1    g044(.A(new_n213_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n233_), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT15), .B1(new_n225_), .B2(new_n229_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n249_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n206_), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n250_), .B(new_n251_), .C1(new_n235_), .C2(new_n242_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n244_), .A2(new_n245_), .A3(new_n252_), .ZN(new_n253_));
  OAI211_X1 g052(.A(KEYINPUT82), .B(new_n206_), .C1(new_n240_), .C2(new_n243_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G190gat), .B(G218gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(G134gat), .ZN(new_n257_));
  INV_X1    g056(.A(G162gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(KEYINPUT36), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT7), .ZN(new_n262_));
  INV_X1    g061(.A(G99gat), .ZN(new_n263_));
  INV_X1    g062(.A(G106gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G99gat), .A2(G106gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT6), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n265_), .A2(new_n268_), .A3(new_n269_), .A4(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT66), .ZN(new_n272_));
  AND3_X1   g071(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(new_n270_), .A4(new_n265_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G85gat), .B(G92gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT67), .B(KEYINPUT8), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n272_), .A2(new_n277_), .A3(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n271_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT8), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT71), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G85gat), .A2(G92gat), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n268_), .B(new_n269_), .C1(KEYINPUT9), .C2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n288_), .B1(KEYINPUT9), .B2(new_n282_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT10), .B(G99gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n290_), .B(KEYINPUT65), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n291_), .B2(G106gat), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n285_), .A2(new_n286_), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n286_), .B1(new_n285_), .B2(new_n292_), .ZN(new_n294_));
  OAI22_X1  g093(.A1(new_n247_), .A2(new_n248_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT68), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n285_), .A2(new_n296_), .A3(new_n292_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n296_), .B1(new_n285_), .B2(new_n292_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n237_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G232gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT75), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT34), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT35), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n295_), .A2(new_n299_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT76), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n302_), .A2(new_n303_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n295_), .A2(new_n308_), .A3(new_n299_), .A4(new_n304_), .ZN(new_n309_));
  AND3_X1   g108(.A1(new_n306_), .A2(new_n307_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n307_), .B1(new_n306_), .B2(new_n309_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n261_), .B1(new_n312_), .B2(KEYINPUT78), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n312_), .A2(KEYINPUT36), .A3(new_n260_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT78), .ZN(new_n315_));
  OAI221_X1 g114(.A(new_n315_), .B1(KEYINPUT36), .B2(new_n260_), .C1(new_n310_), .C2(new_n311_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT37), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G127gat), .B(G155gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G183gat), .B(G211gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT80), .B1(new_n323_), .B2(KEYINPUT17), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(new_n213_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G231gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(G57gat), .ZN(new_n328_));
  INV_X1    g127(.A(G64gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G57gat), .A2(G64gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT69), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n330_), .A2(KEYINPUT69), .A3(new_n331_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT11), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G71gat), .B(G78gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT11), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n334_), .A2(new_n340_), .A3(new_n335_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n336_), .A2(KEYINPUT11), .A3(new_n338_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n327_), .B(new_n345_), .ZN(new_n346_));
  OR2_X1    g145(.A1(new_n323_), .A2(KEYINPUT17), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT37), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n313_), .A2(new_n314_), .A3(new_n349_), .A4(new_n316_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n318_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n352_));
  OR2_X1    g151(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n344_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n285_), .A2(new_n292_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT68), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n285_), .A2(new_n296_), .A3(new_n292_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(new_n345_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT70), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n354_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G230gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT64), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n297_), .A2(new_n298_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(KEYINPUT70), .A3(new_n345_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n360_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT12), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n358_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n362_), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n342_), .A2(KEYINPUT12), .A3(new_n343_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n369_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n367_), .A2(new_n368_), .A3(new_n370_), .A4(new_n354_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G120gat), .B(G148gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(G204gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT5), .ZN(new_n374_));
  INV_X1    g173(.A(G176gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n365_), .A2(new_n371_), .A3(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT72), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT72), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n365_), .A2(new_n371_), .A3(new_n379_), .A4(new_n376_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT73), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n365_), .A2(new_n371_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n376_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n381_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n382_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n352_), .B(new_n353_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n381_), .A2(new_n385_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT73), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n381_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n390_), .A2(KEYINPUT74), .A3(KEYINPUT13), .A4(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n388_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n351_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n255_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT99), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT83), .B(G190gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT26), .ZN(new_n399_));
  INV_X1    g198(.A(G190gat), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n400_), .A2(KEYINPUT26), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT25), .B(G183gat), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n399_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT84), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n203_), .A2(new_n375_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G169gat), .A2(G176gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(KEYINPUT24), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT85), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT24), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(new_n203_), .A3(new_n375_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G183gat), .A2(G190gat), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT23), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n411_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT84), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n399_), .A2(new_n418_), .A3(new_n401_), .A4(new_n402_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n404_), .A2(new_n409_), .A3(new_n417_), .A4(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(G197gat), .B(G204gat), .Z(new_n421_));
  XNOR2_X1  g220(.A(G211gat), .B(G218gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT89), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n421_), .A2(KEYINPUT21), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G197gat), .B(G204gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT21), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n422_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n424_), .A2(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n425_), .A2(new_n426_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n422_), .B(new_n427_), .C1(new_n430_), .C2(new_n423_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n406_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT22), .B(G169gat), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n433_), .B1(new_n434_), .B2(new_n375_), .ZN(new_n435_));
  INV_X1    g234(.A(G183gat), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n398_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n414_), .A2(new_n415_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n435_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n420_), .A2(new_n432_), .A3(new_n439_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n414_), .B(new_n415_), .C1(G183gat), .C2(G190gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n435_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n400_), .A2(KEYINPUT26), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n402_), .A2(new_n401_), .A3(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n445_), .A2(new_n407_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT92), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT91), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n416_), .A2(new_n448_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n411_), .A2(new_n414_), .A3(KEYINPUT91), .A4(new_n415_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n446_), .A2(new_n447_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n449_), .A2(new_n407_), .A3(new_n445_), .A4(new_n450_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT92), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n443_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n440_), .B(KEYINPUT20), .C1(new_n454_), .C2(new_n432_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G226gat), .A2(G233gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT19), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n420_), .A2(new_n439_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n432_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n454_), .A2(new_n432_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n457_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT18), .B(G64gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(G92gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G8gat), .B(G36gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n467_), .B(new_n468_), .Z(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(KEYINPUT32), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n458_), .A2(new_n465_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT90), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n432_), .B(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(new_n442_), .A3(new_n452_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n464_), .B1(new_n474_), .B2(new_n462_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n455_), .A2(new_n457_), .ZN(new_n476_));
  OAI211_X1 g275(.A(KEYINPUT32), .B(new_n469_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT0), .B(G57gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(G85gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(G1gat), .B(G29gat), .Z(new_n480_));
  XOR2_X1   g279(.A(new_n479_), .B(new_n480_), .Z(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT96), .ZN(new_n483_));
  OR2_X1    g282(.A1(G155gat), .A2(G162gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT1), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G155gat), .A2(G162gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G141gat), .A2(G148gat), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(G141gat), .A2(G148gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n487_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT87), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT87), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n487_), .A2(new_n490_), .A3(new_n494_), .A4(new_n491_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n489_), .B(KEYINPUT2), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(KEYINPUT3), .ZN(new_n497_));
  OR3_X1    g296(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n484_), .A2(new_n486_), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n493_), .A2(new_n495_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(G127gat), .A2(G134gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(G113gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G127gat), .A2(G134gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(G127gat), .A2(G134gat), .ZN(new_n507_));
  OAI21_X1  g306(.A(G113gat), .B1(new_n507_), .B2(new_n502_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n506_), .A2(new_n508_), .A3(G120gat), .ZN(new_n509_));
  AOI21_X1  g308(.A(G120gat), .B1(new_n506_), .B2(new_n508_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT93), .B1(new_n501_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n493_), .A2(new_n495_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n499_), .A2(new_n500_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n511_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT94), .ZN(new_n519_));
  AND4_X1   g318(.A1(new_n519_), .A2(new_n511_), .A3(new_n513_), .A4(new_n514_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n519_), .B1(new_n501_), .B2(new_n511_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n512_), .B(new_n518_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G225gat), .A2(G233gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n483_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n521_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n501_), .A2(new_n519_), .A3(new_n511_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n518_), .A2(new_n512_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n528_), .A2(new_n529_), .A3(KEYINPUT96), .A4(new_n523_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n523_), .B(KEYINPUT95), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT4), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n535_));
  AOI21_X1  g334(.A(KEYINPUT4), .B1(new_n515_), .B2(new_n516_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n533_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n482_), .B1(new_n531_), .B2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n536_), .B1(new_n522_), .B2(KEYINPUT4), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n525_), .B(new_n530_), .C1(new_n539_), .C2(new_n532_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n540_), .A2(new_n481_), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n471_), .B(new_n477_), .C1(new_n538_), .C2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT97), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(KEYINPUT33), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(new_n540_), .B2(new_n481_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n544_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n531_), .A2(new_n537_), .A3(new_n482_), .A4(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n458_), .A2(new_n469_), .A3(new_n465_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n469_), .B1(new_n458_), .B2(new_n465_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  OAI221_X1 g349(.A(new_n481_), .B1(new_n532_), .B2(new_n522_), .C1(new_n539_), .C2(new_n524_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n545_), .A2(new_n547_), .A3(new_n550_), .A4(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n542_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G78gat), .B(G106gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n554_), .B(KEYINPUT88), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n515_), .A2(KEYINPUT29), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G228gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n432_), .B(KEYINPUT90), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n515_), .A2(KEYINPUT29), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n558_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n558_), .A3(new_n461_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n557_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n557_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n560_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n473_), .A2(new_n566_), .ZN(new_n567_));
  OAI211_X1 g366(.A(new_n565_), .B(new_n562_), .C1(new_n567_), .C2(new_n558_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n556_), .B1(new_n564_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G22gat), .B(G50gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT28), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n564_), .A2(new_n568_), .A3(new_n556_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n572_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n564_), .A2(new_n568_), .A3(new_n556_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n575_), .B1(new_n576_), .B2(new_n569_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n531_), .A2(new_n537_), .A3(new_n482_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n540_), .A2(new_n481_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n574_), .B2(new_n577_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n469_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n584_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n458_), .A2(new_n465_), .A3(new_n469_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(KEYINPUT27), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT98), .B1(new_n550_), .B2(KEYINPUT27), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT27), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n590_), .B(new_n591_), .C1(new_n548_), .C2(new_n549_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n588_), .B1(new_n589_), .B2(new_n592_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n553_), .A2(new_n579_), .B1(new_n583_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G71gat), .B(G99gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n511_), .B(new_n595_), .Z(new_n596_));
  NAND2_X1  g395(.A1(G227gat), .A2(G233gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT86), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT30), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n596_), .B(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(G15gat), .B(G43gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT31), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n460_), .B(new_n602_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n600_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n603_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n397_), .B1(new_n594_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n606_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n583_), .A2(new_n593_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n578_), .B1(new_n542_), .B2(new_n552_), .ZN(new_n610_));
  OAI211_X1 g409(.A(KEYINPUT99), .B(new_n608_), .C1(new_n609_), .C2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n593_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(new_n578_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n582_), .A2(new_n608_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n607_), .A2(new_n611_), .A3(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT81), .B1(new_n351_), .B2(new_n393_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n396_), .A2(new_n616_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT100), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n208_), .A3(new_n582_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT38), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n348_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n317_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n255_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n388_), .A2(new_n392_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n616_), .A2(new_n625_), .A3(new_n626_), .A4(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n582_), .ZN(new_n629_));
  OAI21_X1  g428(.A(G1gat), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n621_), .A2(new_n622_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n623_), .A2(new_n630_), .A3(new_n631_), .ZN(G1324gat));
  NAND3_X1  g431(.A1(new_n620_), .A2(new_n209_), .A3(new_n612_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G8gat), .B1(new_n628_), .B2(new_n593_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT39), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g436(.A(G15gat), .B1(new_n628_), .B2(new_n608_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT41), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n618_), .A2(G15gat), .A3(new_n608_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n639_), .A2(new_n640_), .ZN(G1326gat));
  OAI21_X1  g440(.A(G22gat), .B1(new_n628_), .B2(new_n579_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT42), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n579_), .A2(G22gat), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT101), .Z(new_n645_));
  OAI21_X1  g444(.A(new_n643_), .B1(new_n618_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT102), .ZN(G1327gat));
  AND2_X1   g446(.A1(new_n616_), .A2(new_n317_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n393_), .A2(new_n348_), .A3(new_n255_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(G29gat), .B1(new_n650_), .B2(new_n582_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT43), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n318_), .A2(new_n350_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n616_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n654_), .B2(KEYINPUT104), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n656_));
  AOI211_X1 g455(.A(new_n656_), .B(KEYINPUT43), .C1(new_n616_), .C2(new_n653_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n649_), .B(KEYINPUT103), .Z(new_n659_));
  AND3_X1   g458(.A1(new_n658_), .A2(KEYINPUT44), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT44), .B1(new_n658_), .B2(new_n659_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(new_n629_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n651_), .B1(new_n664_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g464(.A(G36gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n662_), .B2(new_n612_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT46), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n650_), .A2(new_n666_), .A3(new_n612_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT45), .Z(new_n670_));
  OR3_X1    g469(.A1(new_n667_), .A2(new_n668_), .A3(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n668_), .B1(new_n667_), .B2(new_n670_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1329gat));
  AOI21_X1  g472(.A(G43gat), .B1(new_n650_), .B2(new_n606_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT105), .Z(new_n675_));
  NAND2_X1  g474(.A1(new_n606_), .A2(G43gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n675_), .B1(new_n663_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g477(.A(G50gat), .B1(new_n650_), .B2(new_n578_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n579_), .A2(new_n219_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n662_), .B2(new_n680_), .ZN(G1331gat));
  AND3_X1   g480(.A1(new_n616_), .A2(new_n255_), .A3(new_n393_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n351_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G57gat), .B1(new_n685_), .B2(new_n582_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT106), .ZN(new_n687_));
  OAI21_X1  g486(.A(G57gat), .B1(new_n629_), .B2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n682_), .A2(new_n625_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(KEYINPUT106), .B2(new_n328_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n686_), .B1(new_n688_), .B2(new_n690_), .ZN(G1332gat));
  OAI21_X1  g490(.A(G64gat), .B1(new_n689_), .B2(new_n593_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT48), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n685_), .A2(new_n329_), .A3(new_n612_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1333gat));
  OAI21_X1  g494(.A(G71gat), .B1(new_n689_), .B2(new_n608_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT49), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n608_), .A2(G71gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n697_), .B1(new_n684_), .B2(new_n698_), .ZN(G1334gat));
  OAI21_X1  g498(.A(G78gat), .B1(new_n689_), .B2(new_n579_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT50), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n579_), .A2(G78gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n684_), .B2(new_n702_), .ZN(G1335gat));
  NOR3_X1   g502(.A1(new_n627_), .A2(new_n348_), .A3(new_n626_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n648_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(G85gat), .B1(new_n706_), .B2(new_n582_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n658_), .A2(new_n704_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(new_n582_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n709_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g509(.A(G92gat), .B1(new_n706_), .B2(new_n612_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n612_), .A2(G92gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n708_), .B2(new_n712_), .ZN(G1337gat));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n658_), .A2(new_n606_), .A3(new_n704_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G99gat), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n705_), .A2(new_n608_), .A3(new_n291_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n714_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n718_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n716_), .A2(KEYINPUT107), .A3(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n719_), .A2(KEYINPUT108), .A3(KEYINPUT51), .A4(new_n721_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n719_), .A2(KEYINPUT51), .A3(new_n721_), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n717_), .A2(KEYINPUT51), .A3(new_n718_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT108), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n723_), .B2(new_n726_), .ZN(G1338gat));
  NAND2_X1  g526(.A1(new_n654_), .A2(KEYINPUT104), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT43), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n654_), .A2(KEYINPUT104), .A3(new_n652_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n729_), .A2(new_n578_), .A3(new_n730_), .A4(new_n704_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT109), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n658_), .A2(KEYINPUT109), .A3(new_n578_), .A4(new_n704_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n734_), .A3(G106gat), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT52), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT52), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n733_), .A2(new_n734_), .A3(new_n737_), .A4(G106gat), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n706_), .A2(new_n264_), .A3(new_n578_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT53), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(new_n743_), .A3(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1339gat));
  INV_X1    g544(.A(KEYINPUT54), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n394_), .B2(new_n255_), .ZN(new_n747_));
  NOR4_X1   g546(.A1(new_n351_), .A2(new_n393_), .A3(KEYINPUT54), .A4(new_n626_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n255_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT12), .B1(new_n363_), .B2(new_n345_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n370_), .A2(new_n354_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(KEYINPUT55), .A4(new_n368_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT110), .B1(new_n371_), .B2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n362_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n371_), .A2(new_n756_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n755_), .A2(new_n757_), .A3(new_n758_), .A4(new_n759_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n760_), .A2(KEYINPUT56), .A3(new_n384_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT56), .B1(new_n760_), .B2(new_n384_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n750_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT111), .ZN(new_n764_));
  INV_X1    g563(.A(new_n252_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n206_), .B1(new_n242_), .B2(new_n236_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT112), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT113), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(new_n234_), .B2(new_n239_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n249_), .A2(KEYINPUT113), .A3(new_n238_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n236_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n765_), .B1(new_n767_), .B2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n772_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT111), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n750_), .B(new_n774_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n764_), .A2(new_n773_), .A3(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n317_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT57), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT114), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n776_), .A2(KEYINPUT57), .A3(new_n777_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n381_), .A2(new_n772_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT115), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT115), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n381_), .A2(new_n772_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n761_), .A2(new_n762_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT58), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT58), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n790_), .A2(new_n653_), .A3(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n782_), .A2(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(KEYINPUT57), .B1(new_n776_), .B2(new_n777_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT114), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n781_), .A2(new_n794_), .A3(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n749_), .B1(new_n798_), .B2(new_n624_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n613_), .A2(new_n582_), .A3(new_n606_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(G113gat), .B1(new_n801_), .B2(new_n626_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n782_), .A2(new_n793_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n624_), .B1(new_n803_), .B2(new_n795_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT116), .ZN(new_n805_));
  INV_X1    g604(.A(new_n749_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n624_), .C1(new_n803_), .C2(new_n795_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n805_), .A2(new_n806_), .A3(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810_));
  INV_X1    g609(.A(new_n800_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n809_), .A2(new_n810_), .A3(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT59), .B1(new_n799_), .B2(new_n800_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n814_), .A2(G113gat), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n802_), .B1(new_n815_), .B2(new_n626_), .ZN(G1340gat));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(new_n817_), .A3(new_n393_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n812_), .A2(new_n813_), .A3(new_n393_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT117), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(G120gat), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(G120gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n627_), .B2(KEYINPUT60), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n801_), .B(new_n823_), .C1(KEYINPUT60), .C2(new_n822_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n821_), .A2(new_n824_), .ZN(G1341gat));
  NAND3_X1  g624(.A1(new_n812_), .A2(new_n813_), .A3(new_n348_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(G127gat), .ZN(new_n827_));
  INV_X1    g626(.A(G127gat), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n801_), .A2(new_n828_), .A3(new_n348_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT118), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n827_), .A2(new_n832_), .A3(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1342gat));
  AOI21_X1  g633(.A(G134gat), .B1(new_n801_), .B2(new_n317_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n653_), .ZN(new_n836_));
  XOR2_X1   g635(.A(KEYINPUT119), .B(G134gat), .Z(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n835_), .B1(new_n814_), .B2(new_n838_), .ZN(G1343gat));
  NOR3_X1   g638(.A1(new_n799_), .A2(new_n629_), .A3(new_n606_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n612_), .A2(new_n579_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n626_), .A3(new_n841_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT120), .B(G141gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1344gat));
  NAND3_X1  g643(.A1(new_n840_), .A2(new_n393_), .A3(new_n841_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g645(.A1(new_n840_), .A2(new_n841_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(new_n624_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT61), .B(G155gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(KEYINPUT121), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n848_), .B(new_n850_), .ZN(G1346gat));
  NOR3_X1   g650(.A1(new_n847_), .A2(new_n258_), .A3(new_n836_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n840_), .A2(new_n317_), .A3(new_n841_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n852_), .B1(new_n258_), .B2(new_n853_), .ZN(G1347gat));
  AND4_X1   g653(.A1(new_n579_), .A2(new_n809_), .A3(new_n612_), .A4(new_n614_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n626_), .A2(new_n434_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT123), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n612_), .A2(new_n614_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n255_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n809_), .A2(new_n579_), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n203_), .B1(new_n862_), .B2(KEYINPUT62), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(KEYINPUT62), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n861_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n858_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT124), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT124), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n858_), .B(new_n869_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1348gat));
  AOI21_X1  g670(.A(G176gat), .B1(new_n855_), .B2(new_n393_), .ZN(new_n872_));
  NOR4_X1   g671(.A1(new_n799_), .A2(new_n578_), .A3(new_n627_), .A4(new_n859_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(G176gat), .B2(new_n873_), .ZN(G1349gat));
  NOR2_X1   g673(.A1(new_n799_), .A2(new_n859_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(new_n579_), .A3(new_n348_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT125), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n624_), .A2(new_n402_), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n877_), .A2(new_n436_), .B1(new_n855_), .B2(new_n878_), .ZN(G1350gat));
  NAND4_X1  g678(.A1(new_n855_), .A2(new_n401_), .A3(new_n444_), .A4(new_n317_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT126), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n855_), .A2(new_n653_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(G190gat), .ZN(new_n883_));
  AOI211_X1 g682(.A(KEYINPUT126), .B(new_n400_), .C1(new_n855_), .C2(new_n653_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n880_), .B1(new_n883_), .B2(new_n884_), .ZN(G1351gat));
  INV_X1    g684(.A(new_n583_), .ZN(new_n886_));
  NOR4_X1   g685(.A1(new_n799_), .A2(new_n593_), .A3(new_n606_), .A4(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n626_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n393_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n887_), .A2(new_n348_), .A3(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n893_), .B(new_n894_), .Z(G1354gat));
  INV_X1    g694(.A(G218gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n887_), .A2(new_n896_), .A3(new_n317_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n896_), .B1(new_n887_), .B2(new_n653_), .ZN(new_n899_));
  OAI21_X1  g698(.A(KEYINPUT127), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n899_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT127), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n901_), .A2(new_n902_), .A3(new_n897_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n900_), .A2(new_n903_), .ZN(G1355gat));
endmodule


