//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT19), .ZN(new_n209_));
  INV_X1    g008(.A(G218gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G211gat), .ZN(new_n211_));
  INV_X1    g010(.A(G211gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G218gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT21), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G197gat), .B(G204gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT88), .ZN(new_n218_));
  INV_X1    g017(.A(G197gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n218_), .B1(new_n219_), .B2(G204gat), .ZN(new_n220_));
  INV_X1    g019(.A(G204gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n221_), .A2(KEYINPUT88), .A3(G197gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n219_), .A2(G204gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n220_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(KEYINPUT21), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n216_), .A2(new_n215_), .ZN(new_n226_));
  AOI22_X1  g025(.A1(new_n217_), .A2(new_n225_), .B1(new_n214_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT75), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(KEYINPUT75), .A2(G169gat), .A3(G176gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(G183gat), .A3(G190gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G183gat), .A2(G190gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT23), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n240_), .A2(KEYINPUT76), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT76), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n242_), .B1(new_n239_), .B2(KEYINPUT23), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n238_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n244_));
  NOR3_X1   g043(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT25), .B(G183gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT26), .B(G190gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n245_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n236_), .A2(new_n244_), .A3(new_n248_), .ZN(new_n249_));
  AND2_X1   g048(.A1(KEYINPUT77), .A2(G176gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(KEYINPUT77), .A2(G176gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT22), .B(G169gat), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n252_), .A2(new_n253_), .A3(KEYINPUT78), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT78), .B1(new_n252_), .B2(new_n253_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n233_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n240_), .A2(new_n238_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(G183gat), .A2(G190gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT79), .B1(new_n257_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT79), .ZN(new_n261_));
  AOI211_X1 g060(.A(new_n261_), .B(new_n258_), .C1(new_n240_), .C2(new_n238_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n227_), .B(new_n249_), .C1(new_n256_), .C2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT94), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(new_n265_), .A3(KEYINPUT20), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n244_), .A2(new_n259_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n232_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n235_), .A2(new_n228_), .B1(new_n240_), .B2(new_n238_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n267_), .A2(new_n268_), .B1(new_n248_), .B2(new_n269_), .ZN(new_n270_));
  OR2_X1    g069(.A1(new_n270_), .A2(new_n227_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n265_), .B1(new_n264_), .B2(KEYINPUT20), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n209_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT20), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n275_), .B1(new_n270_), .B2(new_n227_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n209_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n249_), .B1(new_n256_), .B2(new_n263_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n217_), .A2(new_n225_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n226_), .A2(new_n214_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n276_), .A2(new_n277_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n207_), .B1(new_n274_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n273_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n287_), .A2(new_n271_), .A3(new_n266_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n283_), .B1(new_n288_), .B2(new_n209_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n207_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n286_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n274_), .A2(new_n207_), .A3(new_n284_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n293_), .A2(new_n292_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n288_), .A2(new_n209_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n277_), .B1(new_n276_), .B2(new_n282_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n206_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n291_), .A2(new_n292_), .B1(new_n294_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G225gat), .A2(G233gat), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT96), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G127gat), .B(G134gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G113gat), .B(G120gat), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n301_), .A2(new_n302_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G141gat), .B(G148gat), .Z(new_n306_));
  INV_X1    g105(.A(G155gat), .ZN(new_n307_));
  INV_X1    g106(.A(G162gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(new_n308_), .A3(KEYINPUT84), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT84), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n310_), .B1(G155gat), .B2(G162gat), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT1), .B1(new_n307_), .B2(new_n308_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(G155gat), .A3(G162gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n306_), .B1(new_n312_), .B2(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318_));
  NOR2_X1   g117(.A1(KEYINPUT85), .A2(KEYINPUT3), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n324_));
  OAI22_X1  g123(.A1(KEYINPUT85), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n320_), .A2(new_n323_), .A3(new_n324_), .A4(new_n325_), .ZN(new_n326_));
  AOI22_X1  g125(.A1(new_n309_), .A2(new_n311_), .B1(G155gat), .B2(G162gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  AND4_X1   g127(.A1(new_n300_), .A2(new_n305_), .A3(new_n317_), .A4(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n309_), .A2(new_n311_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(new_n313_), .A3(new_n315_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n331_), .A2(new_n306_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n305_), .B1(new_n332_), .B2(new_n300_), .ZN(new_n333_));
  OAI21_X1  g132(.A(KEYINPUT4), .B1(new_n329_), .B2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n317_), .A2(new_n328_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n305_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n299_), .B1(new_n334_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n299_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n329_), .A2(new_n333_), .A3(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G1gat), .B(G29gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(G85gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT0), .B(G57gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  OR3_X1    g143(.A1(new_n338_), .A2(new_n340_), .A3(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n344_), .B1(new_n338_), .B2(new_n340_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n298_), .A2(new_n348_), .ZN(new_n349_));
  XOR2_X1   g148(.A(G22gat), .B(G50gat), .Z(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT29), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n332_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n353_), .B1(new_n332_), .B2(new_n352_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n351_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n353_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(new_n335_), .B2(KEYINPUT29), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(new_n350_), .A3(new_n354_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n364_));
  OAI21_X1  g163(.A(G228gat), .B1(new_n363_), .B2(new_n364_), .ZN(new_n365_));
  OAI211_X1 g164(.A(new_n281_), .B(new_n365_), .C1(new_n352_), .C2(new_n332_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT90), .ZN(new_n367_));
  XOR2_X1   g166(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n368_));
  OAI21_X1  g167(.A(new_n281_), .B1(new_n332_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n365_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n367_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n368_), .B1(new_n317_), .B2(new_n328_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n367_), .B(new_n370_), .C1(new_n372_), .C2(new_n227_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n366_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G78gat), .B(G106gat), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n361_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n366_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n370_), .B1(new_n372_), .B2(new_n227_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT90), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n378_), .B1(new_n380_), .B2(new_n373_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT92), .ZN(new_n382_));
  INV_X1    g181(.A(new_n376_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n383_), .B(new_n366_), .C1(new_n371_), .C2(new_n374_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT92), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n377_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n361_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n375_), .A2(new_n376_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n388_), .B1(new_n389_), .B2(new_n385_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n387_), .B1(new_n390_), .B2(KEYINPUT91), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT91), .ZN(new_n392_));
  AOI211_X1 g191(.A(new_n392_), .B(new_n388_), .C1(new_n389_), .C2(new_n385_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT93), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n381_), .A2(new_n383_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n385_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n361_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n392_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n390_), .A2(KEYINPUT91), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT93), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .A4(new_n387_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n394_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT80), .B(KEYINPUT30), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n278_), .B(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT83), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G15gat), .B(G43gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT81), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G227gat), .A2(G233gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(KEYINPUT82), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n408_), .B(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G71gat), .B(G99gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n406_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n404_), .A2(new_n405_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n413_), .B1(new_n406_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n305_), .B(KEYINPUT31), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n414_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NOR3_X1   g222(.A1(new_n349_), .A2(new_n402_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT97), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT33), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n425_), .B1(new_n346_), .B2(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(KEYINPUT33), .B(new_n344_), .C1(new_n338_), .C2(new_n340_), .ZN(new_n428_));
  OAI22_X1  g227(.A1(new_n335_), .A2(KEYINPUT96), .B1(new_n303_), .B2(new_n304_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n332_), .A2(new_n300_), .A3(new_n305_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n299_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT98), .B1(new_n431_), .B2(new_n344_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n339_), .B1(new_n329_), .B2(new_n333_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n344_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT98), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n334_), .A2(new_n299_), .A3(new_n337_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n432_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n428_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n427_), .A2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n293_), .A2(new_n285_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n346_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n207_), .A2(KEYINPUT32), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n289_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n295_), .A2(new_n296_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n347_), .B(new_n445_), .C1(new_n446_), .C2(new_n444_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n394_), .A2(new_n443_), .A3(new_n401_), .A4(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n423_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n298_), .A2(new_n348_), .B1(new_n394_), .B2(new_n401_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT99), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n349_), .A2(new_n402_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT99), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n452_), .A2(new_n453_), .A3(new_n448_), .A4(new_n423_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n424_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT69), .B(G15gat), .ZN(new_n456_));
  INV_X1    g255(.A(G22gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT14), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT70), .B(G8gat), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n459_), .B1(new_n460_), .B2(G1gat), .ZN(new_n461_));
  OR3_X1    g260(.A1(new_n458_), .A2(KEYINPUT71), .A3(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT71), .B1(new_n458_), .B2(new_n461_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G1gat), .B(G8gat), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n462_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G29gat), .B(G36gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT68), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G43gat), .B(G50gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n473_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n467_), .A2(new_n468_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G229gat), .A2(G233gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n467_), .A2(new_n468_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n473_), .B(KEYINPUT15), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n478_), .B(KEYINPUT74), .Z(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n484_), .B1(new_n469_), .B2(new_n473_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n477_), .A2(new_n479_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G113gat), .B(G141gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G169gat), .B(G197gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n487_), .B(new_n488_), .Z(new_n489_));
  XNOR2_X1  g288(.A(new_n486_), .B(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G120gat), .B(G148gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT5), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G176gat), .B(G204gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G230gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G57gat), .B(G64gat), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(KEYINPUT11), .ZN(new_n500_));
  XOR2_X1   g299(.A(G71gat), .B(G78gat), .Z(new_n501_));
  NAND3_X1  g300(.A1(new_n499_), .A2(new_n500_), .A3(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n500_), .A2(new_n501_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G85gat), .B(G92gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(G99gat), .ZN(new_n507_));
  INV_X1    g306(.A(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT7), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT66), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n509_), .B(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G99gat), .A2(G106gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n513_), .B(KEYINPUT6), .Z(new_n514_));
  OAI21_X1  g313(.A(new_n506_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT8), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT65), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n505_), .A2(KEYINPUT9), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT9), .ZN(new_n519_));
  INV_X1    g318(.A(G85gat), .ZN(new_n520_));
  INV_X1    g319(.A(G92gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT64), .ZN(new_n524_));
  XOR2_X1   g323(.A(KEYINPUT10), .B(G99gat), .Z(new_n525_));
  AOI21_X1  g324(.A(new_n514_), .B1(new_n508_), .B2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n517_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n523_), .A2(KEYINPUT64), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT64), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n529_), .B1(new_n518_), .B2(new_n522_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n526_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(KEYINPUT65), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n504_), .B(new_n516_), .C1(new_n527_), .C2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT12), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n531_), .B(KEYINPUT65), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n504_), .B1(new_n535_), .B2(new_n516_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n516_), .B1(new_n527_), .B2(new_n532_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT12), .ZN(new_n539_));
  INV_X1    g338(.A(new_n504_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n497_), .B1(new_n537_), .B2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n538_), .A2(new_n540_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n497_), .B1(new_n544_), .B2(new_n533_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n496_), .B1(new_n543_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n497_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n544_), .A2(KEYINPUT12), .A3(new_n533_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n549_), .B2(new_n541_), .ZN(new_n550_));
  NOR3_X1   g349(.A1(new_n550_), .A2(new_n545_), .A3(new_n495_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT13), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT13), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(new_n547_), .B2(new_n551_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G127gat), .B(G155gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT16), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G183gat), .B(G211gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT72), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n504_), .B(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n480_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n563_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n469_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n564_), .A2(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n560_), .B1(new_n567_), .B2(KEYINPUT17), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n560_), .A2(KEYINPUT17), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n567_), .A2(KEYINPUT73), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n568_), .B(new_n569_), .C1(KEYINPUT73), .C2(new_n567_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT37), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n481_), .A2(new_n538_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  OAI22_X1  g379(.A1(new_n538_), .A2(new_n475_), .B1(KEYINPUT35), .B2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n576_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n587_), .A2(KEYINPUT36), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT35), .B(new_n580_), .C1(new_n576_), .C2(new_n581_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n584_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n584_), .A2(new_n589_), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n587_), .B(KEYINPUT36), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n575_), .B(new_n590_), .C1(new_n591_), .C2(new_n593_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n584_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n593_), .B1(new_n584_), .B2(new_n589_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT37), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n574_), .B1(new_n594_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR4_X1   g398(.A1(new_n455_), .A2(new_n491_), .A3(new_n556_), .A4(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(G1gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n347_), .B(KEYINPUT100), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n600_), .A2(new_n601_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT38), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OR3_X1    g405(.A1(new_n595_), .A2(new_n596_), .A3(KEYINPUT102), .ZN(new_n607_));
  OAI21_X1  g406(.A(KEYINPUT102), .B1(new_n595_), .B2(new_n596_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n455_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n556_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(KEYINPUT101), .A3(new_n490_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n556_), .B2(new_n491_), .ZN(new_n613_));
  AND4_X1   g412(.A1(new_n572_), .A2(new_n611_), .A3(new_n573_), .A4(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n609_), .A2(new_n614_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n601_), .B1(new_n615_), .B2(new_n347_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n604_), .A2(new_n605_), .ZN(new_n617_));
  OR3_X1    g416(.A1(new_n606_), .A2(new_n616_), .A3(new_n617_), .ZN(G1324gat));
  INV_X1    g417(.A(new_n298_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n609_), .A2(new_n614_), .A3(new_n619_), .ZN(new_n620_));
  AND3_X1   g419(.A1(new_n620_), .A2(KEYINPUT39), .A3(G8gat), .ZN(new_n621_));
  AOI21_X1  g420(.A(KEYINPUT39), .B1(new_n620_), .B2(G8gat), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n460_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n600_), .A2(new_n619_), .A3(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT103), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n623_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n627_), .B1(new_n623_), .B2(new_n626_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1325gat));
  NAND2_X1  g429(.A1(new_n615_), .A2(new_n422_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT105), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n632_), .A3(G15gat), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n632_), .B1(new_n631_), .B2(G15gat), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT41), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n635_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT41), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(new_n633_), .ZN(new_n639_));
  INV_X1    g438(.A(G15gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n600_), .A2(new_n640_), .A3(new_n422_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT106), .Z(new_n642_));
  NAND3_X1  g441(.A1(new_n636_), .A2(new_n639_), .A3(new_n642_), .ZN(G1326gat));
  XOR2_X1   g442(.A(new_n402_), .B(KEYINPUT107), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n600_), .A2(new_n457_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n615_), .A2(new_n644_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(G22gat), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(KEYINPUT42), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(KEYINPUT42), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(G1327gat));
  NAND3_X1  g449(.A1(new_n607_), .A2(new_n574_), .A3(new_n608_), .ZN(new_n651_));
  NOR4_X1   g450(.A1(new_n455_), .A2(new_n491_), .A3(new_n556_), .A4(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(G29gat), .B1(new_n652_), .B2(new_n347_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n611_), .A2(new_n574_), .A3(new_n613_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n451_), .A2(new_n454_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n424_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n594_), .A2(new_n597_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n657_), .A2(new_n658_), .A3(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT43), .B1(new_n455_), .B2(new_n659_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n654_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT44), .ZN(new_n664_));
  AND3_X1   g463(.A1(new_n664_), .A2(G29gat), .A3(new_n603_), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n663_), .A2(KEYINPUT44), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n653_), .B1(new_n665_), .B2(new_n666_), .ZN(G1328gat));
  AOI21_X1  g466(.A(new_n298_), .B1(new_n663_), .B2(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(G36gat), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT108), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n298_), .A2(G36gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n652_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n651_), .A2(new_n556_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n657_), .A2(new_n490_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n672_), .ZN(new_n676_));
  OAI21_X1  g475(.A(KEYINPUT108), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n673_), .A2(new_n677_), .A3(KEYINPUT45), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n673_), .A2(new_n677_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT45), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n670_), .A2(KEYINPUT46), .A3(new_n678_), .A4(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT46), .ZN(new_n683_));
  INV_X1    g482(.A(G36gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n684_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n681_), .A2(new_n678_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n682_), .A2(new_n687_), .ZN(G1329gat));
  INV_X1    g487(.A(G43gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n689_), .B1(new_n675_), .B2(new_n423_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n664_), .A2(G43gat), .A3(new_n422_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n663_), .A2(KEYINPUT44), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n690_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT47), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT47), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n695_), .B(new_n690_), .C1(new_n691_), .C2(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(G1330gat));
  AOI21_X1  g496(.A(G50gat), .B1(new_n652_), .B2(new_n644_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n664_), .A2(G50gat), .A3(new_n402_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n666_), .ZN(G1331gat));
  NAND2_X1  g499(.A1(new_n607_), .A2(new_n608_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n657_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n556_), .A2(new_n491_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n702_), .A2(new_n574_), .A3(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(G57gat), .A3(new_n347_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n705_), .A2(new_n706_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n455_), .A2(new_n490_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n599_), .A2(new_n610_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(G57gat), .B1(new_n712_), .B2(new_n603_), .ZN(new_n713_));
  NOR3_X1   g512(.A1(new_n707_), .A2(new_n708_), .A3(new_n713_), .ZN(G1332gat));
  INV_X1    g513(.A(G64gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n704_), .B2(new_n619_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT48), .Z(new_n717_));
  NAND2_X1  g516(.A1(new_n619_), .A2(new_n715_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT110), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n711_), .B2(new_n719_), .ZN(G1333gat));
  INV_X1    g519(.A(G71gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n721_), .B1(new_n704_), .B2(new_n422_), .ZN(new_n722_));
  XOR2_X1   g521(.A(new_n722_), .B(KEYINPUT49), .Z(new_n723_));
  NAND2_X1  g522(.A1(new_n422_), .A2(new_n721_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT111), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n723_), .B1(new_n711_), .B2(new_n725_), .ZN(G1334gat));
  INV_X1    g525(.A(G78gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n704_), .B2(new_n644_), .ZN(new_n728_));
  XOR2_X1   g527(.A(new_n728_), .B(KEYINPUT50), .Z(new_n729_));
  NAND3_X1  g528(.A1(new_n712_), .A2(new_n727_), .A3(new_n644_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1335gat));
  INV_X1    g530(.A(new_n574_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n703_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n658_), .B1(new_n657_), .B2(new_n660_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n455_), .A2(KEYINPUT43), .A3(new_n659_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n733_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT113), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  OAI211_X1 g537(.A(KEYINPUT113), .B(new_n733_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n347_), .A2(G85gat), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT114), .ZN(new_n742_));
  NOR4_X1   g541(.A1(new_n455_), .A2(new_n490_), .A3(new_n610_), .A4(new_n651_), .ZN(new_n743_));
  AOI21_X1  g542(.A(G85gat), .B1(new_n743_), .B2(new_n603_), .ZN(new_n744_));
  OR2_X1    g543(.A1(new_n744_), .A2(KEYINPUT112), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(KEYINPUT112), .ZN(new_n746_));
  AOI22_X1  g545(.A1(new_n740_), .A2(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(G1336gat));
  NAND3_X1  g546(.A1(new_n743_), .A2(new_n521_), .A3(new_n619_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n298_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(new_n521_), .ZN(G1337gat));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n422_), .A2(new_n525_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n743_), .B2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n423_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(new_n507_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT51), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(new_n753_), .C1(new_n754_), .C2(new_n507_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1338gat));
  NAND3_X1  g558(.A1(new_n743_), .A2(new_n508_), .A3(new_n402_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n402_), .B(new_n733_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(new_n762_), .A3(G106gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(G106gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT53), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n760_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1339gat));
  INV_X1    g568(.A(G113gat), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n598_), .A2(new_n491_), .A3(new_n553_), .A4(new_n555_), .ZN(new_n771_));
  XOR2_X1   g570(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n771_), .A2(KEYINPUT117), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n771_), .A2(KEYINPUT117), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n771_), .B2(KEYINPUT117), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n774_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n486_), .A2(new_n489_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n489_), .B1(new_n477_), .B2(new_n483_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n482_), .A2(new_n474_), .A3(new_n484_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n784_), .A2(new_n551_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n537_), .A2(new_n497_), .A3(new_n542_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n543_), .A2(KEYINPUT55), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n550_), .A2(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n786_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n790_), .A2(new_n791_), .A3(new_n496_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n786_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n550_), .A2(new_n788_), .ZN(new_n794_));
  AOI211_X1 g593(.A(KEYINPUT55), .B(new_n548_), .C1(new_n549_), .C2(new_n541_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n793_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT56), .B1(new_n796_), .B2(new_n495_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n785_), .B1(new_n792_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT58), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n659_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(KEYINPUT58), .B(new_n785_), .C1(new_n792_), .C2(new_n797_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n543_), .A2(new_n546_), .A3(new_n496_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n490_), .A2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n791_), .B1(new_n790_), .B2(new_n496_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n796_), .A2(KEYINPUT56), .A3(new_n495_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n804_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(KEYINPUT118), .B1(new_n552_), .B2(new_n784_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n784_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n809_), .B(new_n810_), .C1(new_n547_), .C2(new_n551_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n701_), .B1(new_n807_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT57), .B(new_n701_), .C1(new_n807_), .C2(new_n812_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n802_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n574_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n779_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n402_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n619_), .A2(new_n423_), .A3(new_n602_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n770_), .B1(new_n822_), .B2(new_n491_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT119), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n825_), .B(new_n770_), .C1(new_n822_), .C2(new_n491_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(KEYINPUT59), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n822_), .A2(new_n828_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .A4(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n491_), .A2(new_n770_), .ZN(new_n833_));
  AOI22_X1  g632(.A1(new_n824_), .A2(new_n826_), .B1(new_n832_), .B2(new_n833_), .ZN(G1340gat));
  INV_X1    g633(.A(new_n822_), .ZN(new_n835_));
  INV_X1    g634(.A(G120gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n610_), .B2(KEYINPUT60), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n835_), .B(new_n837_), .C1(KEYINPUT60), .C2(new_n836_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n610_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n836_), .ZN(G1341gat));
  INV_X1    g639(.A(G127gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n835_), .A2(new_n841_), .A3(new_n732_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n574_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n841_), .ZN(G1342gat));
  INV_X1    g643(.A(G134gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n822_), .B2(new_n701_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT121), .B(new_n845_), .C1(new_n822_), .C2(new_n701_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n659_), .A2(new_n845_), .ZN(new_n850_));
  AOI22_X1  g649(.A1(new_n848_), .A2(new_n849_), .B1(new_n832_), .B2(new_n850_), .ZN(G1343gat));
  NOR3_X1   g650(.A1(new_n619_), .A2(new_n422_), .A3(new_n602_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n801_), .A2(new_n800_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n732_), .B1(new_n853_), .B2(new_n816_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n402_), .B(new_n852_), .C1(new_n854_), .C2(new_n778_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n855_), .A2(new_n491_), .ZN(new_n856_));
  XOR2_X1   g655(.A(new_n856_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g656(.A1(new_n855_), .A2(new_n610_), .ZN(new_n858_));
  XOR2_X1   g657(.A(new_n858_), .B(G148gat), .Z(G1345gat));
  INV_X1    g658(.A(KEYINPUT122), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n855_), .B2(new_n574_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n820_), .B1(new_n779_), .B2(new_n818_), .ZN(new_n862_));
  NAND4_X1  g661(.A1(new_n862_), .A2(KEYINPUT122), .A3(new_n732_), .A4(new_n852_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n861_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1346gat));
  NOR3_X1   g666(.A1(new_n855_), .A2(new_n308_), .A3(new_n659_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n308_), .B1(new_n855_), .B2(new_n701_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  OAI211_X1 g670(.A(KEYINPUT123), .B(new_n308_), .C1(new_n855_), .C2(new_n701_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n868_), .B1(new_n871_), .B2(new_n872_), .ZN(G1347gat));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n874_));
  NOR3_X1   g673(.A1(new_n603_), .A2(new_n423_), .A3(new_n298_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n644_), .A2(new_n876_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n490_), .B(new_n877_), .C1(new_n854_), .C2(new_n778_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n874_), .B1(new_n878_), .B2(G169gat), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n878_), .A2(new_n874_), .A3(G169gat), .ZN(new_n881_));
  XOR2_X1   g680(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n880_), .A2(new_n881_), .A3(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n878_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n879_), .A2(new_n882_), .B1(new_n253_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n886_), .ZN(G1348gat));
  AOI21_X1  g686(.A(new_n778_), .B1(new_n574_), .B2(new_n817_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n877_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n556_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n888_), .A2(new_n402_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n875_), .A2(new_n556_), .A3(G176gat), .ZN(new_n893_));
  AOI22_X1  g692(.A1(new_n891_), .A2(new_n252_), .B1(new_n892_), .B2(new_n893_), .ZN(G1349gat));
  INV_X1    g693(.A(new_n890_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n895_), .A2(new_n246_), .A3(new_n574_), .ZN(new_n896_));
  INV_X1    g695(.A(G183gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n892_), .A2(new_n732_), .A3(new_n875_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n896_), .B1(new_n897_), .B2(new_n898_), .ZN(G1350gat));
  OAI21_X1  g698(.A(G190gat), .B1(new_n895_), .B2(new_n659_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n607_), .A2(new_n247_), .A3(new_n608_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n895_), .B2(new_n901_), .ZN(G1351gat));
  NOR3_X1   g701(.A1(new_n298_), .A2(new_n422_), .A3(new_n347_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n862_), .A2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n904_), .A2(new_n491_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(new_n219_), .ZN(G1352gat));
  INV_X1    g705(.A(new_n904_), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n907_), .B(new_n556_), .C1(KEYINPUT126), .C2(new_n221_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n904_), .A2(new_n610_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT126), .B(G204gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n909_), .B2(new_n910_), .ZN(G1353gat));
  XOR2_X1   g710(.A(KEYINPUT63), .B(G211gat), .Z(new_n912_));
  NAND3_X1  g711(.A1(new_n907_), .A2(new_n732_), .A3(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n914_), .B1(new_n904_), .B2(new_n574_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n913_), .A2(new_n915_), .ZN(G1354gat));
  OAI21_X1  g715(.A(G218gat), .B1(new_n904_), .B2(new_n659_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n607_), .A2(new_n210_), .A3(new_n608_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n904_), .B2(new_n918_), .ZN(G1355gat));
endmodule


