//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n841_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n851_, new_n852_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT15), .Z(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n205_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G229gat), .A2(G233gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(new_n213_), .B2(new_n204_), .ZN(new_n217_));
  XOR2_X1   g016(.A(new_n212_), .B(new_n204_), .Z(new_n218_));
  AOI22_X1  g017(.A1(new_n214_), .A2(new_n217_), .B1(new_n218_), .B2(new_n216_), .ZN(new_n219_));
  XOR2_X1   g018(.A(G113gat), .B(G141gat), .Z(new_n220_));
  XNOR2_X1  g019(.A(G169gat), .B(G197gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n219_), .A2(new_n222_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G155gat), .B(G162gat), .Z(new_n226_));
  INV_X1    g025(.A(KEYINPUT1), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G141gat), .A2(G148gat), .ZN(new_n229_));
  INV_X1    g028(.A(G141gat), .ZN(new_n230_));
  INV_X1    g029(.A(G148gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n228_), .A2(new_n229_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n229_), .A2(KEYINPUT79), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n236_), .B(new_n237_), .C1(new_n238_), .C2(KEYINPUT2), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n238_), .A2(KEYINPUT2), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n226_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n234_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT80), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT29), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT28), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT81), .ZN(new_n249_));
  XOR2_X1   g048(.A(G22gat), .B(G50gat), .Z(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT81), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n248_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n250_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT21), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT84), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G211gat), .B(G218gat), .ZN(new_n259_));
  AOI211_X1 g058(.A(new_n256_), .B(new_n257_), .C1(new_n258_), .C2(new_n259_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT83), .B(KEYINPUT21), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(new_n262_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n257_), .A2(KEYINPUT82), .ZN(new_n264_));
  INV_X1    g063(.A(G197gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(G204gat), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT21), .B1(new_n266_), .B2(KEYINPUT82), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n263_), .B(new_n259_), .C1(new_n264_), .C2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n261_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n245_), .B1(new_n234_), .B2(new_n241_), .ZN(new_n271_));
  OAI211_X1 g070(.A(G228gat), .B(G233gat), .C1(new_n270_), .C2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT85), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n270_), .B1(G228gat), .B2(G233gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(new_n245_), .B2(new_n244_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G78gat), .B(G106gat), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n278_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n251_), .A2(new_n255_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(KEYINPUT87), .ZN(new_n282_));
  OR3_X1    g081(.A1(new_n277_), .A2(KEYINPUT87), .A3(new_n278_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n282_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n251_), .A2(new_n255_), .ZN(new_n285_));
  OAI22_X1  g084(.A1(new_n281_), .A2(KEYINPUT86), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n281_), .A2(KEYINPUT86), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G1gat), .B(G29gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(G85gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT0), .B(G57gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n290_), .B(new_n291_), .Z(new_n292_));
  XNOR2_X1  g091(.A(G127gat), .B(G134gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT77), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G113gat), .B(G120gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n244_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n296_), .A2(new_n242_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  MUX2_X1   g099(.A(new_n298_), .B(new_n300_), .S(KEYINPUT4), .Z(new_n301_));
  AND2_X1   g100(.A1(G225gat), .A2(G233gat), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n300_), .A2(new_n302_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n292_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n304_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n292_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT92), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT92), .B1(new_n305_), .B2(new_n308_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT26), .B(G190gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT73), .B1(new_n316_), .B2(G183gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT25), .B(G183gat), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n315_), .B(new_n317_), .C1(new_n318_), .C2(KEYINPUT73), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT74), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT23), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n321_), .B1(G183gat), .B2(G190gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n323_), .A2(KEYINPUT23), .ZN(new_n324_));
  INV_X1    g123(.A(G169gat), .ZN(new_n325_));
  INV_X1    g124(.A(G176gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  OAI22_X1  g126(.A1(new_n322_), .A2(new_n324_), .B1(KEYINPUT24), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT24), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n328_), .B1(new_n327_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n320_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT22), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n326_), .B1(new_n334_), .B2(KEYINPUT75), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n335_), .A2(G169gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n323_), .A2(new_n321_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n337_), .B(new_n338_), .C1(G183gat), .C2(G190gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(G169gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n336_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n333_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G227gat), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(G71gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(G99gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n342_), .B(new_n347_), .Z(new_n348_));
  XOR2_X1   g147(.A(KEYINPUT78), .B(KEYINPUT31), .Z(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G15gat), .B(G43gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n351_), .B(KEYINPUT76), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT30), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n296_), .B(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(new_n350_), .B(new_n354_), .Z(new_n355_));
  NOR2_X1   g154(.A1(new_n314_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n342_), .A2(new_n269_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n357_), .A2(KEYINPUT20), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G226gat), .A2(G233gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT19), .ZN(new_n360_));
  XOR2_X1   g159(.A(KEYINPUT22), .B(G169gat), .Z(new_n361_));
  OAI211_X1 g160(.A(new_n339_), .B(new_n329_), .C1(G176gat), .C2(new_n361_), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n328_), .B(KEYINPUT89), .Z(new_n363_));
  AOI22_X1  g162(.A1(new_n330_), .A2(KEYINPUT88), .B1(new_n325_), .B2(new_n326_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n364_), .B1(KEYINPUT88), .B2(new_n330_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n318_), .A2(new_n315_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n362_), .B1(new_n363_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n360_), .B1(new_n369_), .B2(new_n270_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n358_), .A2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n371_), .A2(KEYINPUT90), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(KEYINPUT90), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n269_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n375_), .B(KEYINPUT20), .C1(new_n342_), .C2(new_n269_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n360_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT18), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  NAND3_X1  g180(.A1(new_n374_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT93), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AOI22_X1  g183(.A1(new_n372_), .A2(new_n373_), .B1(new_n360_), .B2(new_n376_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(KEYINPUT93), .A3(new_n381_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT27), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n376_), .A2(new_n360_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n358_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT91), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n269_), .B1(new_n369_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n368_), .A2(KEYINPUT91), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n390_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n360_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n389_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n381_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n388_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n387_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT94), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT94), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n387_), .A2(new_n401_), .A3(new_n398_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n385_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n397_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT27), .B1(new_n405_), .B2(new_n382_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT95), .B1(new_n403_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT95), .ZN(new_n409_));
  AOI211_X1 g208(.A(new_n409_), .B(new_n406_), .C1(new_n400_), .C2(new_n402_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n288_), .B(new_n356_), .C1(new_n408_), .C2(new_n410_), .ZN(new_n411_));
  AND2_X1   g210(.A1(new_n381_), .A2(KEYINPUT32), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n396_), .A2(new_n412_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n309_), .B(new_n413_), .C1(new_n404_), .C2(new_n412_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT33), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n305_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n292_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n416_), .A2(new_n382_), .A3(new_n405_), .A4(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n305_), .A2(new_n415_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n414_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n288_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n402_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n401_), .B1(new_n387_), .B2(new_n398_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n407_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n313_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n422_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n355_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n225_), .B1(new_n411_), .B2(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G85gat), .B(G92gat), .Z(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT9), .ZN(new_n431_));
  XOR2_X1   g230(.A(KEYINPUT10), .B(G99gat), .Z(new_n432_));
  INV_X1    g231(.A(G106gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G99gat), .A2(G106gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT6), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(G99gat), .A3(G106gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT65), .B(G92gat), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT9), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(G85gat), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n431_), .A2(new_n434_), .A3(new_n439_), .A4(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n346_), .A2(new_n433_), .A3(KEYINPUT67), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT67), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n445_), .B1(G99gat), .B2(G106gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT7), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n444_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT68), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT66), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  OAI211_X1 g252(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n453_), .A2(new_n454_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n444_), .A2(new_n446_), .A3(KEYINPUT68), .A4(new_n447_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n450_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT8), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n457_), .A2(new_n458_), .A3(new_n430_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n457_), .B2(new_n430_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n443_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G57gat), .B(G64gat), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n462_), .A2(KEYINPUT11), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(KEYINPUT11), .ZN(new_n464_));
  XOR2_X1   g263(.A(G71gat), .B(G78gat), .Z(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n464_), .A2(new_n465_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n461_), .A2(new_n469_), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n468_), .B(new_n443_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(KEYINPUT12), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT12), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n461_), .A2(new_n473_), .A3(new_n469_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G230gat), .A2(G233gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT64), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT69), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n470_), .A2(new_n471_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n477_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT69), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n483_), .A3(new_n477_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n479_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G120gat), .B(G148gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT5), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G176gat), .B(G204gat), .ZN(new_n488_));
  XOR2_X1   g287(.A(new_n487_), .B(new_n488_), .Z(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n479_), .A2(new_n482_), .A3(new_n484_), .A4(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n494_), .A2(KEYINPUT13), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(KEYINPUT13), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n498_), .A2(KEYINPUT70), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(KEYINPUT70), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G190gat), .B(G218gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G134gat), .B(G162gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n505_), .B(KEYINPUT36), .Z(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n461_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n508_), .A2(new_n205_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G232gat), .A2(G233gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT35), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n508_), .A2(new_n204_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n509_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n512_), .A2(new_n513_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n517_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n507_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n505_), .A2(KEYINPUT36), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n518_), .A2(new_n522_), .A3(new_n519_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(KEYINPUT72), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n525_), .A3(KEYINPUT37), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT37), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n521_), .B(new_n523_), .C1(KEYINPUT72), .C2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n213_), .B(new_n468_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G231gat), .A2(G233gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535_));
  XOR2_X1   g334(.A(G127gat), .B(G155gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT16), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  OR3_X1    g338(.A1(new_n534_), .A2(new_n535_), .A3(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(KEYINPUT17), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n534_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n530_), .A2(new_n543_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n429_), .A2(new_n502_), .A3(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n545_), .A2(new_n207_), .A3(new_n314_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT38), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n524_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n411_), .B2(new_n428_), .ZN(new_n550_));
  NOR3_X1   g349(.A1(new_n497_), .A2(new_n225_), .A3(new_n543_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(G1gat), .B1(new_n553_), .B2(new_n313_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n546_), .A2(new_n547_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n548_), .A2(new_n554_), .A3(new_n555_), .ZN(G1324gat));
  XNOR2_X1  g355(.A(KEYINPUT97), .B(KEYINPUT40), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n408_), .A2(new_n410_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n552_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(G8gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT96), .B(KEYINPUT39), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n561_), .B(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n545_), .A2(new_n208_), .A3(new_n559_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n557_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n561_), .A2(new_n563_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n562_), .B1(new_n560_), .B2(G8gat), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n565_), .B(new_n557_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n566_), .A2(new_n570_), .ZN(G1325gat));
  INV_X1    g370(.A(G15gat), .ZN(new_n572_));
  INV_X1    g371(.A(new_n355_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n545_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n574_), .B(KEYINPUT98), .Z(new_n575_));
  OAI21_X1  g374(.A(G15gat), .B1(new_n553_), .B2(new_n355_), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n576_), .A2(KEYINPUT41), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(KEYINPUT41), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n575_), .A2(new_n577_), .A3(new_n578_), .ZN(G1326gat));
  INV_X1    g378(.A(G22gat), .ZN(new_n580_));
  INV_X1    g379(.A(new_n288_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n552_), .B2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT42), .Z(new_n583_));
  NAND3_X1  g382(.A1(new_n545_), .A2(new_n580_), .A3(new_n581_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(G1327gat));
  INV_X1    g384(.A(new_n543_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n524_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n497_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n429_), .A2(new_n589_), .ZN(new_n590_));
  OR3_X1    g389(.A1(new_n590_), .A2(G29gat), .A3(new_n313_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n225_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n498_), .A2(new_n592_), .A3(new_n543_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT99), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT43), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n411_), .A2(new_n428_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n595_), .B1(new_n596_), .B2(new_n530_), .ZN(new_n597_));
  AOI211_X1 g396(.A(KEYINPUT43), .B(new_n529_), .C1(new_n411_), .C2(new_n428_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n594_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT44), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  OAI211_X1 g400(.A(KEYINPUT44), .B(new_n594_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n314_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(G29gat), .B1(new_n603_), .B2(new_n604_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n591_), .B1(new_n605_), .B2(new_n606_), .ZN(G1328gat));
  NAND3_X1  g406(.A1(new_n601_), .A2(new_n559_), .A3(new_n602_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(G36gat), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n590_), .A2(G36gat), .A3(new_n558_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT101), .B(KEYINPUT45), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n609_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT46), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n609_), .A2(KEYINPUT46), .A3(new_n612_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(G1329gat));
  INV_X1    g416(.A(new_n590_), .ZN(new_n618_));
  AOI21_X1  g417(.A(G43gat), .B1(new_n618_), .B2(new_n573_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT102), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n601_), .A2(G43gat), .A3(new_n573_), .A4(new_n602_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT47), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT47), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n620_), .A2(new_n624_), .A3(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(G1330gat));
  AOI21_X1  g425(.A(G50gat), .B1(new_n618_), .B2(new_n581_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n601_), .A2(new_n602_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n581_), .A2(G50gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n627_), .B1(new_n628_), .B2(new_n629_), .ZN(G1331gat));
  NAND2_X1  g429(.A1(new_n596_), .A2(new_n225_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n544_), .A2(new_n497_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT103), .Z(new_n633_));
  NOR2_X1   g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(G57gat), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(new_n635_), .A3(new_n314_), .ZN(new_n636_));
  AND4_X1   g435(.A1(new_n225_), .A2(new_n550_), .A3(new_n501_), .A4(new_n586_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(new_n314_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n636_), .B1(new_n638_), .B2(new_n635_), .ZN(G1332gat));
  INV_X1    g438(.A(G64gat), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n637_), .B2(new_n559_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(KEYINPUT104), .B(KEYINPUT48), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n641_), .B(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n634_), .A2(new_n640_), .A3(new_n559_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1333gat));
  AOI21_X1  g444(.A(new_n344_), .B1(new_n637_), .B2(new_n573_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT49), .Z(new_n647_));
  NOR2_X1   g446(.A1(new_n355_), .A2(G71gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT105), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n634_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(G1334gat));
  INV_X1    g450(.A(G78gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n652_), .B1(new_n637_), .B2(new_n581_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT50), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n634_), .A2(new_n652_), .A3(new_n581_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1335gat));
  NAND2_X1  g455(.A1(new_n596_), .A2(new_n530_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT43), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT107), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n596_), .A2(new_n595_), .A3(new_n530_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n658_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT107), .B1(new_n597_), .B2(new_n598_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n497_), .A2(new_n225_), .A3(new_n543_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT108), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n661_), .A2(new_n662_), .A3(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G85gat), .B1(new_n665_), .B2(new_n313_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n592_), .B1(new_n411_), .B2(new_n428_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n501_), .A2(new_n587_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n667_), .A2(new_n669_), .A3(KEYINPUT106), .ZN(new_n670_));
  AOI21_X1  g469(.A(KEYINPUT106), .B1(new_n667_), .B2(new_n669_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n313_), .A2(G85gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n666_), .B1(new_n672_), .B2(new_n673_), .ZN(G1336gat));
  INV_X1    g473(.A(new_n665_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n559_), .A2(new_n440_), .ZN(new_n676_));
  INV_X1    g475(.A(G92gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n559_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n678_));
  AOI22_X1  g477(.A1(new_n675_), .A2(new_n676_), .B1(new_n677_), .B2(new_n678_), .ZN(G1337gat));
  OAI21_X1  g478(.A(G99gat), .B1(new_n665_), .B2(new_n355_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n573_), .A2(new_n432_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n681_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT109), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT109), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n684_), .B(new_n681_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n680_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT51), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT51), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n680_), .A2(new_n686_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1338gat));
  OAI211_X1 g490(.A(new_n581_), .B(new_n664_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT52), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(G106gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n692_), .B2(G106gat), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n581_), .A2(new_n433_), .ZN(new_n696_));
  OAI22_X1  g495(.A1(new_n694_), .A2(new_n695_), .B1(new_n672_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g497(.A(KEYINPUT118), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT115), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n313_), .A2(new_n355_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n558_), .A2(new_n700_), .A3(new_n288_), .A4(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n288_), .B(new_n701_), .C1(new_n408_), .C2(new_n410_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(KEYINPUT115), .ZN(new_n704_));
  XNOR2_X1  g503(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n702_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n492_), .A2(new_n592_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n475_), .A2(KEYINPUT110), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n472_), .A2(new_n709_), .A3(new_n474_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n708_), .A2(new_n481_), .A3(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT111), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT55), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n479_), .A2(new_n713_), .A3(new_n484_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n475_), .A2(KEYINPUT55), .A3(new_n477_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT112), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n475_), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(new_n477_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n708_), .A2(new_n720_), .A3(new_n710_), .A4(new_n481_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n712_), .A2(new_n714_), .A3(new_n719_), .A4(new_n721_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n722_), .A2(KEYINPUT56), .A3(new_n489_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT56), .B1(new_n722_), .B2(new_n489_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n707_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n218_), .A2(new_n215_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n215_), .B1(new_n213_), .B2(new_n204_), .ZN(new_n727_));
  AOI211_X1 g526(.A(new_n222_), .B(new_n726_), .C1(new_n214_), .C2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n728_), .A2(new_n223_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT113), .B1(new_n493_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT113), .ZN(new_n731_));
  INV_X1    g530(.A(new_n729_), .ZN(new_n732_));
  AOI211_X1 g531(.A(new_n731_), .B(new_n732_), .C1(new_n490_), .C2(new_n492_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n730_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n725_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n735_), .A2(KEYINPUT57), .A3(new_n524_), .ZN(new_n736_));
  AOI21_X1  g535(.A(KEYINPUT57), .B1(new_n735_), .B2(new_n524_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT58), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n492_), .A2(new_n729_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n722_), .A2(new_n489_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT56), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n722_), .A2(KEYINPUT56), .A3(new_n489_), .ZN(new_n743_));
  AOI211_X1 g542(.A(new_n738_), .B(new_n739_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n739_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n745_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n529_), .B1(new_n746_), .B2(new_n738_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT114), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n530_), .B1(new_n750_), .B2(KEYINPUT58), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT114), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n737_), .B1(new_n749_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT117), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n736_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n737_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n744_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n751_), .B2(KEYINPUT114), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n747_), .A2(new_n748_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n756_), .B(new_n754_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n543_), .B1(new_n755_), .B2(new_n761_), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n498_), .A2(new_n225_), .A3(new_n586_), .A4(new_n529_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT54), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n706_), .B1(new_n762_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT59), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n756_), .B(new_n736_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n768_), .B2(new_n586_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n703_), .B(new_n700_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n699_), .B1(new_n765_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT54), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n763_), .B(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n543_), .B2(new_n767_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n702_), .A2(new_n704_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT59), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n756_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT117), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(new_n736_), .A3(new_n760_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n774_), .B1(new_n780_), .B2(new_n543_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n777_), .B(KEYINPUT118), .C1(new_n781_), .C2(new_n706_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n592_), .A2(KEYINPUT119), .A3(G113gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(KEYINPUT119), .B2(G113gat), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n772_), .A2(new_n782_), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(G113gat), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n775_), .A2(new_n776_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n786_), .B1(new_n788_), .B2(new_n225_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT120), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT120), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n785_), .A2(new_n792_), .A3(new_n789_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n791_), .A2(new_n793_), .ZN(G1340gat));
  INV_X1    g593(.A(G120gat), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n498_), .B2(KEYINPUT60), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n787_), .B(new_n796_), .C1(KEYINPUT60), .C2(new_n795_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n777_), .B(new_n501_), .C1(new_n781_), .C2(new_n706_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n797_), .B1(new_n799_), .B2(new_n795_), .ZN(G1341gat));
  NAND3_X1  g599(.A1(new_n772_), .A2(new_n586_), .A3(new_n782_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(G127gat), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n543_), .A2(G127gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n788_), .B2(new_n803_), .ZN(G1342gat));
  XOR2_X1   g603(.A(KEYINPUT121), .B(G134gat), .Z(new_n805_));
  AND4_X1   g604(.A1(new_n530_), .A2(new_n772_), .A3(new_n782_), .A4(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(G134gat), .B1(new_n787_), .B2(new_n549_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(G1343gat));
  NOR4_X1   g607(.A1(new_n559_), .A2(new_n288_), .A3(new_n313_), .A4(new_n573_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT122), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n769_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n769_), .B2(new_n809_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n225_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(KEYINPUT123), .B(G141gat), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(G1344gat));
  NOR2_X1   g615(.A1(new_n813_), .A2(new_n502_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(new_n231_), .ZN(G1345gat));
  INV_X1    g617(.A(new_n813_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n586_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT61), .B(G155gat), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(G1346gat));
  OR3_X1    g621(.A1(new_n813_), .A2(G162gat), .A3(new_n524_), .ZN(new_n823_));
  OAI21_X1  g622(.A(G162gat), .B1(new_n813_), .B2(new_n529_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(G1347gat));
  NAND2_X1  g624(.A1(new_n762_), .A2(new_n764_), .ZN(new_n826_));
  NOR4_X1   g625(.A1(new_n558_), .A2(new_n581_), .A3(new_n314_), .A4(new_n355_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n592_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(G169gat), .B1(new_n828_), .B2(new_n225_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT62), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n831_), .B(new_n834_), .C1(new_n361_), .C2(new_n830_), .ZN(G1348gat));
  NAND2_X1  g634(.A1(new_n769_), .A2(new_n827_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n836_), .A2(new_n326_), .A3(new_n502_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT124), .ZN(new_n838_));
  AOI21_X1  g637(.A(G176gat), .B1(new_n829_), .B2(new_n497_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1349gat));
  NOR2_X1   g639(.A1(new_n543_), .A2(new_n318_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT125), .B1(new_n828_), .B2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n836_), .A2(new_n543_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(G183gat), .B2(new_n844_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n828_), .A2(KEYINPUT125), .A3(new_n842_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1350gat));
  OAI21_X1  g646(.A(G190gat), .B1(new_n828_), .B2(new_n529_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n549_), .A2(new_n315_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n828_), .B2(new_n849_), .ZN(G1351gat));
  NOR4_X1   g649(.A1(new_n775_), .A2(new_n558_), .A3(new_n573_), .A4(new_n426_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n592_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n501_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g654(.A(new_n543_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n851_), .A2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT126), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(KEYINPUT127), .B2(new_n859_), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(KEYINPUT127), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n857_), .B2(new_n861_), .ZN(G1354gat));
  INV_X1    g661(.A(G218gat), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n851_), .A2(new_n863_), .A3(new_n549_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n851_), .A2(new_n530_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n865_), .B2(new_n863_), .ZN(G1355gat));
endmodule


