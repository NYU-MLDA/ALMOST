//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT25), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT25), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT26), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT26), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(G190gat), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n209_), .A2(new_n211_), .A3(new_n213_), .A4(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(KEYINPUT24), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT24), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n207_), .A2(new_n216_), .A3(new_n220_), .A4(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT22), .B(G169gat), .ZN(new_n224_));
  INV_X1    g023(.A(G176gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n205_), .B(new_n206_), .C1(G183gat), .C2(G190gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(new_n219_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT21), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G197gat), .A2(G204gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(G197gat), .A2(G204gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n229_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OR2_X1    g032(.A1(G197gat), .A2(G204gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n234_), .A2(KEYINPUT21), .A3(new_n230_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G211gat), .B(G218gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n233_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(G211gat), .B(G218gat), .Z(new_n238_));
  NAND4_X1  g037(.A1(new_n238_), .A2(KEYINPUT21), .A3(new_n234_), .A4(new_n230_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n223_), .A2(new_n228_), .A3(new_n237_), .A4(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT100), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n240_), .A2(new_n241_), .A3(KEYINPUT20), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n241_), .B1(new_n240_), .B2(KEYINPUT20), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n239_), .A2(new_n237_), .ZN(new_n244_));
  AOI21_X1  g043(.A(G176gat), .B1(KEYINPUT82), .B2(KEYINPUT22), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(G169gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(new_n227_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n222_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n219_), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n249_), .A2(new_n217_), .A3(new_n221_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n209_), .A2(new_n211_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n213_), .A2(new_n215_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(KEYINPUT81), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT81), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n216_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n251_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n244_), .B1(new_n247_), .B2(new_n257_), .ZN(new_n258_));
  NOR3_X1   g057(.A1(new_n242_), .A2(new_n243_), .A3(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G226gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT101), .B1(new_n259_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n243_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT20), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n249_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n251_), .A2(new_n216_), .B1(new_n227_), .B2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n266_), .B1(new_n268_), .B2(new_n244_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n241_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n258_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n265_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT101), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n262_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT94), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n275_), .B1(new_n268_), .B2(new_n244_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n223_), .A2(new_n228_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n239_), .A2(new_n237_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(KEYINPUT94), .A3(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n244_), .A2(new_n257_), .A3(new_n247_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n276_), .A2(KEYINPUT20), .A3(new_n279_), .A4(new_n280_), .ZN(new_n281_));
  OR2_X1    g080(.A1(new_n281_), .A2(new_n262_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n264_), .A2(new_n274_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT102), .ZN(new_n284_));
  XOR2_X1   g083(.A(G8gat), .B(G36gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT18), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G64gat), .B(G92gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n283_), .A2(new_n284_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n257_), .A2(new_n247_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n262_), .B1(new_n291_), .B2(new_n278_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n281_), .A2(new_n262_), .B1(new_n269_), .B2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT102), .B1(new_n293_), .B2(new_n288_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n294_), .B1(new_n283_), .B2(new_n289_), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT27), .B1(new_n290_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n281_), .A2(new_n262_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n292_), .A2(new_n269_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n288_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT95), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n293_), .A2(KEYINPUT95), .A3(new_n288_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n298_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(new_n289_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n301_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n305_));
  OR2_X1    g104(.A1(new_n305_), .A2(KEYINPUT27), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n296_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT90), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT89), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT2), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT2), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(G141gat), .A3(G148gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT87), .B(KEYINPUT3), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n319_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT88), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  OAI211_X1 g125(.A(KEYINPUT88), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n314_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT3), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT87), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT87), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT3), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n334_), .A2(new_n321_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n326_), .A2(new_n327_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(KEYINPUT89), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n313_), .B1(new_n329_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n322_), .A2(new_n315_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n312_), .A2(KEYINPUT1), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT86), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n312_), .A2(KEYINPUT1), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n342_), .A2(new_n310_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n339_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n309_), .B1(new_n338_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n313_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n334_), .A2(new_n321_), .ZN(new_n347_));
  AND4_X1   g146(.A1(KEYINPUT89), .A2(new_n347_), .A3(new_n336_), .A4(new_n319_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT89), .B1(new_n335_), .B2(new_n336_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n346_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n344_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(KEYINPUT90), .A3(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n345_), .A2(new_n352_), .A3(KEYINPUT29), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n244_), .B1(G228gat), .B2(G233gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n356_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n357_));
  OAI211_X1 g156(.A(G228gat), .B(G233gat), .C1(new_n357_), .C2(new_n244_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G78gat), .B(G106gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(KEYINPUT90), .B1(new_n350_), .B2(new_n351_), .ZN(new_n362_));
  NOR3_X1   g161(.A1(new_n338_), .A2(new_n309_), .A3(new_n344_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n356_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT28), .ZN(new_n365_));
  XOR2_X1   g164(.A(G22gat), .B(G50gat), .Z(new_n366_));
  NAND2_X1  g165(.A1(new_n345_), .A2(new_n352_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT28), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n367_), .A2(new_n368_), .A3(new_n356_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(new_n366_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n366_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n368_), .B1(new_n367_), .B2(new_n356_), .ZN(new_n372_));
  AOI211_X1 g171(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n345_), .C2(new_n352_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n371_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n361_), .A2(new_n370_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n360_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(KEYINPUT91), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n355_), .A2(new_n358_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n378_), .B1(new_n355_), .B2(new_n358_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n374_), .A2(new_n370_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT92), .ZN(new_n383_));
  AND3_X1   g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n383_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n375_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n308_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G113gat), .B(G120gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G127gat), .B(G134gat), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(KEYINPUT83), .ZN(new_n391_));
  INV_X1    g190(.A(G134gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G127gat), .ZN(new_n393_));
  INV_X1    g192(.A(G127gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(G134gat), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n393_), .A2(new_n395_), .A3(KEYINPUT83), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n389_), .B1(new_n391_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n393_), .A2(new_n395_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT83), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n390_), .A2(KEYINPUT83), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n400_), .A2(new_n401_), .A3(new_n388_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n397_), .A2(KEYINPUT84), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT84), .B1(new_n397_), .B2(new_n402_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n345_), .A2(new_n352_), .A3(new_n405_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n350_), .A2(new_n402_), .A3(new_n397_), .A4(new_n351_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G225gat), .A2(G233gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G1gat), .B(G29gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(G85gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(KEYINPUT0), .B(G57gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n345_), .A2(new_n352_), .A3(new_n416_), .A4(new_n405_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT97), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n406_), .A2(new_n407_), .A3(KEYINPUT4), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n408_), .B(KEYINPUT96), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n415_), .B1(new_n418_), .B2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT97), .ZN(new_n423_));
  AND2_X1   g222(.A1(new_n417_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n417_), .A2(new_n423_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n419_), .B(new_n420_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n426_), .A2(new_n409_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n422_), .B1(new_n427_), .B2(new_n413_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G227gat), .A2(G233gat), .ZN(new_n429_));
  INV_X1    g228(.A(G15gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT30), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n291_), .B(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(G71gat), .B(G99gat), .Z(new_n434_));
  XNOR2_X1  g233(.A(new_n434_), .B(G43gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n433_), .B(new_n435_), .ZN(new_n436_));
  OR3_X1    g235(.A1(new_n403_), .A2(new_n404_), .A3(KEYINPUT31), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT31), .B1(new_n403_), .B2(new_n404_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n439_), .A2(KEYINPUT85), .ZN(new_n440_));
  OR2_X1    g239(.A1(new_n436_), .A2(new_n440_), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n439_), .A2(KEYINPUT85), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n436_), .B1(new_n442_), .B2(new_n440_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n441_), .A2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n428_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n387_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n381_), .A2(new_n382_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT92), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n428_), .B1(new_n450_), .B2(new_n375_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n359_), .B(new_n376_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n452_), .A2(new_n382_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n454_));
  OAI211_X1 g253(.A(new_n419_), .B(new_n408_), .C1(new_n424_), .C2(new_n425_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n406_), .A2(new_n407_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n413_), .B1(new_n456_), .B2(new_n420_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n305_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT98), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(KEYINPUT33), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n422_), .A2(new_n460_), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n426_), .B(new_n415_), .C1(new_n459_), .C2(KEYINPUT33), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n458_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n288_), .A2(KEYINPUT32), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT99), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n464_), .B1(new_n303_), .B2(new_n465_), .ZN(new_n466_));
  OAI211_X1 g265(.A(KEYINPUT32), .B(new_n288_), .C1(new_n303_), .C2(KEYINPUT99), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n466_), .B1(new_n467_), .B2(new_n283_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n413_), .B1(new_n426_), .B2(new_n409_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n421_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n417_), .B(new_n423_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n414_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n468_), .B1(new_n469_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n463_), .A2(new_n473_), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n451_), .A2(new_n307_), .B1(new_n454_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n444_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n446_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n478_));
  INV_X1    g277(.A(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT64), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT6), .ZN(new_n484_));
  INV_X1    g283(.A(G85gat), .ZN(new_n485_));
  INV_X1    g284(.A(G92gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G85gat), .A2(G92gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(KEYINPUT9), .A3(new_n488_), .ZN(new_n489_));
  OR3_X1    g288(.A1(new_n485_), .A2(new_n486_), .A3(KEYINPUT9), .ZN(new_n490_));
  AND3_X1   g289(.A1(new_n484_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n482_), .A2(KEYINPUT65), .A3(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(KEYINPUT65), .B1(new_n482_), .B2(new_n491_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n494_), .A2(KEYINPUT66), .ZN(new_n495_));
  OR3_X1    g294(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(KEYINPUT66), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n484_), .A2(new_n495_), .A3(new_n496_), .A4(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT8), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n487_), .A2(new_n488_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n499_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n503_));
  OAI22_X1  g302(.A1(new_n492_), .A2(new_n493_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT67), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n482_), .A2(new_n491_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT65), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n482_), .A2(new_n491_), .A3(KEYINPUT65), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n503_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n501_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT67), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n510_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G29gat), .B(G36gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G43gat), .B(G50gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n505_), .A2(new_n514_), .A3(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(KEYINPUT15), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n504_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G232gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT34), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n518_), .B(new_n520_), .C1(KEYINPUT35), .C2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n522_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n520_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n526_), .B1(new_n527_), .B2(KEYINPUT73), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n518_), .A2(KEYINPUT73), .A3(new_n520_), .A4(new_n526_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G190gat), .B(G218gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G134gat), .B(G162gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT74), .B(KEYINPUT36), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n531_), .A2(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(KEYINPUT75), .B(KEYINPUT36), .Z(new_n538_));
  XNOR2_X1  g337(.A(new_n534_), .B(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n529_), .A2(new_n539_), .A3(new_n530_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n477_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G127gat), .B(G155gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G183gat), .B(G211gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G57gat), .B(G64gat), .Z(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT69), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT11), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G57gat), .B(G64gat), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT69), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n552_), .A2(new_n553_), .A3(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(KEYINPUT68), .B(G71gat), .ZN(new_n558_));
  INV_X1    g357(.A(G78gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT70), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n552_), .A2(new_n556_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n562_), .B1(new_n563_), .B2(KEYINPUT11), .ZN(new_n564_));
  AOI211_X1 g363(.A(KEYINPUT70), .B(new_n553_), .C1(new_n552_), .C2(new_n556_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n561_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n554_), .B(KEYINPUT69), .ZN(new_n567_));
  OAI21_X1  g366(.A(KEYINPUT70), .B1(new_n567_), .B2(new_n553_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n563_), .A2(new_n562_), .A3(KEYINPUT11), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n568_), .A2(new_n557_), .A3(new_n569_), .A4(new_n560_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G15gat), .B(G22gat), .ZN(new_n572_));
  INV_X1    g371(.A(G8gat), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G1gat), .B(G8gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n575_), .B(new_n576_), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n571_), .B(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G231gat), .A2(G233gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n580_), .A2(new_n549_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n550_), .B1(new_n581_), .B2(new_n548_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT79), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n583_), .A3(new_n580_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n583_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n585_), .B(new_n550_), .C1(new_n581_), .C2(new_n548_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n566_), .A2(new_n570_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(new_n505_), .B2(new_n514_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n590_), .A2(KEYINPUT12), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G230gat), .A2(G233gat), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n505_), .A2(new_n514_), .A3(new_n589_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n571_), .A2(KEYINPUT12), .A3(new_n504_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n591_), .A2(new_n592_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n592_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n593_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n597_), .B1(new_n598_), .B2(new_n590_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G120gat), .B(G148gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(KEYINPUT5), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G176gat), .B(G204gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT71), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n600_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n596_), .A2(new_n599_), .A3(new_n604_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(KEYINPUT72), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT72), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n600_), .A2(new_n609_), .A3(new_n605_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT13), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT13), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n608_), .A2(new_n613_), .A3(new_n610_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n577_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n519_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n577_), .A2(new_n517_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n621_), .A2(KEYINPUT80), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(KEYINPUT80), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n577_), .B(new_n517_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(G229gat), .A3(G233gat), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n622_), .A2(new_n623_), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G113gat), .B(G141gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G169gat), .B(G197gat), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n627_), .B(new_n628_), .Z(new_n629_));
  XNOR2_X1  g428(.A(new_n626_), .B(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(KEYINPUT103), .B1(new_n615_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT103), .ZN(new_n632_));
  INV_X1    g431(.A(new_n630_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n612_), .A2(new_n632_), .A3(new_n633_), .A4(new_n614_), .ZN(new_n634_));
  AND4_X1   g433(.A1(new_n543_), .A2(new_n588_), .A3(new_n631_), .A4(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n202_), .B1(new_n635_), .B2(new_n428_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT104), .Z(new_n637_));
  AND3_X1   g436(.A1(new_n445_), .A2(new_n454_), .A3(new_n307_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n474_), .A2(new_n454_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n469_), .A2(new_n472_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n386_), .A2(new_n640_), .A3(new_n307_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n638_), .B1(new_n642_), .B2(new_n444_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(new_n630_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n531_), .A2(new_n536_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n539_), .B(KEYINPUT76), .Z(new_n646_));
  NOR2_X1   g445(.A1(new_n531_), .A2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT37), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT37), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n537_), .A2(new_n649_), .A3(new_n540_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n650_), .A3(KEYINPUT77), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT77), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n652_), .B(KEYINPUT37), .C1(new_n645_), .C2(new_n647_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n615_), .A2(new_n654_), .A3(new_n587_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n644_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n202_), .A3(new_n428_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT38), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n637_), .A2(new_n659_), .ZN(G1324gat));
  NAND3_X1  g459(.A1(new_n657_), .A2(new_n573_), .A3(new_n308_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT39), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n635_), .A2(new_n308_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n663_), .B2(G8gat), .ZN(new_n664_));
  AOI211_X1 g463(.A(KEYINPUT39), .B(new_n573_), .C1(new_n635_), .C2(new_n308_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n661_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT40), .Z(G1325gat));
  AOI21_X1  g466(.A(new_n430_), .B1(new_n635_), .B2(new_n476_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n668_), .B(KEYINPUT41), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n657_), .A2(new_n430_), .A3(new_n476_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1326gat));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n635_), .B2(new_n386_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT42), .Z(new_n674_));
  NAND3_X1  g473(.A1(new_n657_), .A2(new_n672_), .A3(new_n386_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1327gat));
  NOR3_X1   g475(.A1(new_n615_), .A2(new_n588_), .A3(new_n541_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n644_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G29gat), .B1(new_n679_), .B2(new_n428_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT105), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n477_), .A2(new_n681_), .A3(new_n682_), .A4(new_n654_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n476_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n682_), .B(new_n654_), .C1(new_n684_), .C2(new_n638_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT105), .ZN(new_n686_));
  INV_X1    g485(.A(new_n654_), .ZN(new_n687_));
  OAI21_X1  g486(.A(KEYINPUT43), .B1(new_n643_), .B2(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n683_), .A2(new_n686_), .A3(new_n688_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n631_), .A2(new_n587_), .A3(new_n634_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n689_), .A2(KEYINPUT44), .A3(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n428_), .A2(G29gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n680_), .B1(new_n696_), .B2(new_n697_), .ZN(G1328gat));
  NOR3_X1   g497(.A1(new_n678_), .A2(G36gat), .A3(new_n307_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT45), .Z(new_n700_));
  NAND3_X1  g499(.A1(new_n693_), .A2(new_n308_), .A3(new_n694_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT106), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n701_), .A2(new_n702_), .A3(G36gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n701_), .B2(G36gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT46), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n700_), .B(KEYINPUT46), .C1(new_n703_), .C2(new_n704_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1329gat));
  NAND2_X1  g508(.A1(new_n476_), .A2(G43gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n678_), .A2(new_n444_), .ZN(new_n711_));
  OAI22_X1  g510(.A1(new_n695_), .A2(new_n710_), .B1(G43gat), .B2(new_n711_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g512(.A(G50gat), .B1(new_n679_), .B2(new_n386_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n386_), .A2(G50gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n696_), .B2(new_n715_), .ZN(G1331gat));
  INV_X1    g515(.A(new_n615_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(new_n633_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n543_), .A2(new_n588_), .A3(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G57gat), .B1(new_n719_), .B2(new_n640_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n643_), .A2(new_n717_), .A3(new_n633_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(new_n588_), .A3(new_n687_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n640_), .A2(G57gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT107), .Z(G1332gat));
  OAI21_X1  g524(.A(G64gat), .B1(new_n719_), .B2(new_n307_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT48), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n307_), .A2(G64gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n722_), .B2(new_n728_), .ZN(G1333gat));
  OAI21_X1  g528(.A(G71gat), .B1(new_n719_), .B2(new_n444_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n730_), .B(new_n731_), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n444_), .A2(G71gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n722_), .B2(new_n733_), .ZN(G1334gat));
  OAI21_X1  g533(.A(G78gat), .B1(new_n719_), .B2(new_n454_), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n735_), .B(KEYINPUT50), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n386_), .A2(new_n559_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n722_), .B2(new_n737_), .ZN(G1335gat));
  NOR2_X1   g537(.A1(new_n588_), .A2(new_n541_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n721_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n485_), .B1(new_n740_), .B2(new_n640_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT109), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n718_), .A2(new_n587_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n689_), .A2(new_n744_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n745_), .A2(new_n485_), .A3(new_n640_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n742_), .A2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT110), .ZN(G1336gat));
  OAI21_X1  g547(.A(G92gat), .B1(new_n745_), .B2(new_n307_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n740_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n486_), .A3(new_n308_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1337gat));
  OAI21_X1  g551(.A(G99gat), .B1(new_n745_), .B2(new_n444_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n476_), .A2(new_n478_), .A3(new_n480_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n740_), .B2(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g555(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n689_), .A2(new_n744_), .A3(new_n386_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G106gat), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(KEYINPUT52), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(KEYINPUT52), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n750_), .A2(new_n479_), .A3(new_n386_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n757_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n763_), .B(new_n757_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  INV_X1    g566(.A(KEYINPUT57), .ZN(new_n768_));
  INV_X1    g567(.A(new_n629_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n626_), .A2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n619_), .A2(G229gat), .A3(G233gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n629_), .B1(new_n624_), .B2(new_n620_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n608_), .A2(new_n610_), .A3(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n593_), .B(new_n594_), .C1(new_n590_), .C2(KEYINPUT12), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n597_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(KEYINPUT112), .B(new_n775_), .C1(new_n776_), .C2(new_n597_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n591_), .A2(KEYINPUT55), .A3(new_n592_), .A4(new_n595_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n776_), .A2(new_n597_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .A4(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n605_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n605_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(KEYINPUT113), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT113), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n783_), .A2(new_n789_), .A3(KEYINPUT56), .A4(new_n605_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n607_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n630_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n774_), .B1(new_n788_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n541_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n768_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n787_), .A2(KEYINPUT113), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n793_), .B1(new_n798_), .B2(new_n786_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT57), .B(new_n541_), .C1(new_n799_), .C2(new_n774_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n773_), .A2(new_n607_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n605_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(new_n787_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n783_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n605_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n801_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(KEYINPUT115), .A2(KEYINPUT58), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n654_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n787_), .A2(new_n803_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(new_n786_), .A3(new_n805_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(new_n607_), .A3(new_n773_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(new_n807_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n797_), .B(new_n800_), .C1(new_n809_), .C2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n587_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n655_), .A2(new_n816_), .A3(new_n630_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n816_), .B1(new_n655_), .B2(new_n630_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n815_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n387_), .A2(new_n428_), .A3(new_n476_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT59), .ZN(new_n825_));
  INV_X1    g624(.A(G113gat), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n630_), .A2(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT118), .ZN(new_n828_));
  INV_X1    g627(.A(new_n800_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n797_), .B1(new_n809_), .B2(new_n813_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(KEYINPUT117), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n832_), .B(new_n797_), .C1(new_n809_), .C2(new_n813_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n588_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n834_), .A2(new_n819_), .ZN(new_n835_));
  XOR2_X1   g634(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n836_));
  NAND2_X1  g635(.A1(new_n823_), .A2(new_n836_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n825_), .B(new_n828_), .C1(new_n835_), .C2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n826_), .B1(new_n824_), .B2(new_n630_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(G1340gat));
  OAI211_X1 g639(.A(new_n825_), .B(new_n615_), .C1(new_n835_), .C2(new_n837_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(G120gat), .ZN(new_n842_));
  INV_X1    g641(.A(G120gat), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n717_), .B2(KEYINPUT60), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(KEYINPUT60), .B2(new_n843_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n824_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n846_), .ZN(G1341gat));
  NAND2_X1  g646(.A1(new_n588_), .A2(G127gat), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT119), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n825_), .B(new_n849_), .C1(new_n835_), .C2(new_n837_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n394_), .B1(new_n824_), .B2(new_n587_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1342gat));
  XOR2_X1   g651(.A(KEYINPUT120), .B(G134gat), .Z(new_n853_));
  NOR2_X1   g652(.A1(new_n687_), .A2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n825_), .B(new_n854_), .C1(new_n835_), .C2(new_n837_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n392_), .B1(new_n824_), .B2(new_n541_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(G1343gat));
  AOI21_X1  g656(.A(new_n819_), .B1(new_n587_), .B2(new_n814_), .ZN(new_n858_));
  NOR4_X1   g657(.A1(new_n308_), .A2(new_n454_), .A3(new_n640_), .A4(new_n476_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n633_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT121), .B(G141gat), .Z(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1344gat));
  NAND2_X1  g663(.A1(new_n861_), .A2(new_n615_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT122), .B(G148gat), .Z(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1345gat));
  NAND3_X1  g666(.A1(new_n861_), .A2(KEYINPUT123), .A3(new_n588_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n821_), .A2(new_n588_), .A3(new_n859_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT123), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n868_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1346gat));
  AOI21_X1  g674(.A(G162gat), .B1(new_n861_), .B2(new_n796_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n654_), .A2(G162gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT124), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n861_), .B2(new_n878_), .ZN(G1347gat));
  NAND3_X1  g678(.A1(new_n445_), .A2(new_n308_), .A3(new_n454_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n835_), .A2(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n633_), .A2(new_n224_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT125), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n880_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n633_), .B(new_n885_), .C1(new_n834_), .C2(new_n819_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT62), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n886_), .A2(new_n887_), .A3(G169gat), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n886_), .B2(G169gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n884_), .B1(new_n888_), .B2(new_n889_), .ZN(G1348gat));
  NOR4_X1   g689(.A1(new_n858_), .A2(new_n225_), .A3(new_n717_), .A4(new_n880_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n881_), .A2(new_n615_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n225_), .ZN(G1349gat));
  NOR2_X1   g692(.A1(new_n587_), .A2(new_n252_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n821_), .A2(new_n588_), .A3(new_n885_), .ZN(new_n895_));
  AOI22_X1  g694(.A1(new_n881_), .A2(new_n894_), .B1(new_n208_), .B2(new_n895_), .ZN(G1350gat));
  NAND3_X1  g695(.A1(new_n881_), .A2(new_n253_), .A3(new_n796_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n835_), .A2(new_n687_), .A3(new_n880_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n212_), .B2(new_n898_), .ZN(G1351gat));
  NAND3_X1  g698(.A1(new_n451_), .A2(new_n308_), .A3(new_n444_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n858_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n633_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g702(.A(new_n900_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n821_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n717_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1353gat));
  NAND2_X1  g707(.A1(new_n901_), .A2(new_n588_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n910_));
  AND2_X1   g709(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n909_), .A2(new_n910_), .A3(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n909_), .B2(new_n910_), .ZN(G1354gat));
  INV_X1    g712(.A(G218gat), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n901_), .A2(new_n914_), .A3(new_n796_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n905_), .A2(new_n687_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n914_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT127), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n915_), .B(KEYINPUT127), .C1(new_n916_), .C2(new_n914_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(G1355gat));
endmodule


