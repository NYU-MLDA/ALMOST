//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n777_, new_n778_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n878_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT9), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n206_), .A2(KEYINPUT65), .A3(G85gat), .ZN(new_n207_));
  OR2_X1    g006(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(G92gat), .ZN(new_n210_));
  INV_X1    g009(.A(G92gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(G85gat), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G92gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT9), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n210_), .A2(new_n216_), .A3(KEYINPUT66), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n211_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n206_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G106gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT10), .B(G99gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n224_), .A2(new_n225_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n223_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT6), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n222_), .A2(new_n228_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT7), .ZN(new_n236_));
  INV_X1    g035(.A(G99gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n223_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n238_), .A2(new_n231_), .A3(new_n232_), .A4(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(KEYINPUT67), .B1(new_n212_), .B2(new_n214_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT8), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT8), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n244_), .A3(new_n241_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G29gat), .B(G36gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G43gat), .B(G50gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n235_), .A2(new_n246_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT70), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n233_), .B1(new_n217_), .B2(new_n221_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n252_), .A2(new_n228_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT70), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(new_n249_), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT35), .ZN(new_n257_));
  INV_X1    g056(.A(new_n245_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n244_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260_));
  NOR3_X1   g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT69), .B1(new_n243_), .B2(new_n245_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n235_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n249_), .B(KEYINPUT15), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT72), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n256_), .A2(new_n257_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n265_), .A2(new_n267_), .A3(new_n251_), .A4(new_n255_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G232gat), .A2(G233gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n269_), .B(KEYINPUT34), .Z(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n256_), .A2(new_n267_), .A3(new_n265_), .A4(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n266_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n271_), .A2(new_n273_), .A3(KEYINPUT35), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n205_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n271_), .A2(new_n273_), .A3(KEYINPUT35), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n280_), .A2(new_n274_), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT73), .B1(new_n281_), .B2(new_n205_), .ZN(new_n282_));
  AND4_X1   g081(.A1(KEYINPUT73), .A2(new_n275_), .A3(new_n205_), .A4(new_n276_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n279_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT74), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n285_), .A2(KEYINPUT37), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n285_), .A2(KEYINPUT37), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n284_), .A2(new_n287_), .A3(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n275_), .A2(new_n205_), .A3(new_n276_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n281_), .A2(KEYINPUT73), .A3(new_n205_), .ZN(new_n294_));
  AOI22_X1  g093(.A1(new_n293_), .A2(new_n294_), .B1(new_n278_), .B2(new_n277_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(new_n285_), .A3(KEYINPUT37), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n290_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(G190gat), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT25), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT79), .B1(new_n300_), .B2(G183gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT25), .B(G183gat), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n299_), .B(new_n301_), .C1(new_n302_), .C2(KEYINPUT79), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT80), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305_));
  INV_X1    g104(.A(G169gat), .ZN(new_n306_));
  INV_X1    g105(.A(G176gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT24), .ZN(new_n310_));
  NOR2_X1   g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n308_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(KEYINPUT23), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n312_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT79), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n300_), .A2(G183gat), .ZN(new_n320_));
  INV_X1    g119(.A(G183gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n321_), .A2(KEYINPUT25), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n319_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT80), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n323_), .A2(new_n324_), .A3(new_n299_), .A4(new_n301_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n304_), .A2(new_n318_), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n306_), .A2(KEYINPUT22), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n327_), .A2(KEYINPUT82), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(KEYINPUT82), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT22), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(G169gat), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n328_), .A2(new_n329_), .A3(new_n307_), .A4(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n314_), .A2(KEYINPUT23), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(KEYINPUT81), .B(KEYINPUT23), .Z(new_n335_));
  INV_X1    g134(.A(new_n314_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n334_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(G183gat), .A2(G190gat), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n332_), .B(new_n309_), .C1(new_n337_), .C2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n326_), .A2(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT30), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n340_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G227gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT83), .ZN(new_n345_));
  XOR2_X1   g144(.A(G71gat), .B(G99gat), .Z(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n343_), .B(new_n347_), .Z(new_n348_));
  XNOR2_X1  g147(.A(G127gat), .B(G134gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G113gat), .B(G120gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G15gat), .B(G43gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n348_), .B(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(G155gat), .ZN(new_n355_));
  INV_X1    g154(.A(G162gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(new_n356_), .A3(KEYINPUT86), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT86), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(G155gat), .B2(G162gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT1), .B1(new_n355_), .B2(new_n356_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT87), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n355_), .A2(new_n356_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT1), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT87), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n360_), .A2(new_n367_), .A3(new_n361_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n363_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G141gat), .A2(G148gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(KEYINPUT85), .A2(G141gat), .A3(G148gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(G141gat), .A2(G148gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n364_), .B1(new_n359_), .B2(new_n357_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT88), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n378_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT2), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n372_), .A2(new_n382_), .A3(new_n373_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n380_), .A2(new_n379_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n381_), .A2(new_n383_), .A3(new_n384_), .A4(new_n385_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n369_), .A2(new_n376_), .B1(new_n377_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n388_));
  OAI21_X1  g187(.A(KEYINPUT89), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT89), .ZN(new_n390_));
  INV_X1    g189(.A(new_n376_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n360_), .A2(new_n367_), .A3(new_n361_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n367_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n391_), .B1(new_n394_), .B2(new_n366_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n386_), .A2(new_n377_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n390_), .B(KEYINPUT29), .C1(new_n395_), .C2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT92), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G211gat), .A2(G218gat), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(G211gat), .A2(G218gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n399_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G211gat), .ZN(new_n404_));
  INV_X1    g203(.A(G218gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(KEYINPUT92), .A3(new_n400_), .ZN(new_n407_));
  INV_X1    g206(.A(G197gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(G204gat), .ZN(new_n409_));
  INV_X1    g208(.A(G204gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(G197gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n403_), .A2(new_n407_), .A3(KEYINPUT21), .A4(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT21), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n408_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n415_), .A2(new_n411_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT90), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(new_n410_), .B2(G197gat), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n414_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n406_), .A2(new_n400_), .ZN(new_n420_));
  XOR2_X1   g219(.A(KEYINPUT91), .B(KEYINPUT21), .Z(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(new_n421_), .B2(new_n412_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n413_), .B1(new_n419_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(KEYINPUT93), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n418_), .A2(new_n415_), .A3(new_n411_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT21), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G197gat), .B(G204gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n420_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT93), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n413_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n424_), .A2(new_n432_), .B1(G228gat), .B2(G233gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n389_), .A2(new_n398_), .A3(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n423_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(G228gat), .A3(G233gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G78gat), .B(G106gat), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n434_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n438_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n369_), .A2(new_n376_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(new_n388_), .A3(new_n396_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT28), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT28), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n387_), .A2(new_n444_), .A3(new_n388_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G22gat), .B(G50gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n443_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n447_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n449_));
  OAI22_X1  g248(.A1(new_n439_), .A2(new_n440_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n434_), .A2(new_n436_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n437_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n448_), .A2(new_n449_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n434_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n450_), .A2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G8gat), .B(G36gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(G92gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT18), .B(G64gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G226gat), .A2(G233gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT19), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n327_), .A2(new_n331_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(new_n307_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n316_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n465_), .B(new_n309_), .C1(new_n466_), .C2(new_n338_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n333_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n310_), .A2(new_n311_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n302_), .A2(new_n299_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n308_), .A4(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n467_), .A2(new_n471_), .A3(new_n430_), .A4(new_n413_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT94), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT20), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n424_), .A2(new_n432_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n475_), .B1(new_n476_), .B2(new_n340_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n463_), .B1(new_n474_), .B2(new_n477_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n424_), .A2(new_n432_), .A3(new_n339_), .A4(new_n326_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n467_), .A2(new_n471_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n423_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n479_), .A2(KEYINPUT20), .A3(new_n463_), .A4(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n461_), .B1(new_n478_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT95), .ZN(new_n485_));
  INV_X1    g284(.A(new_n463_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n430_), .A2(new_n431_), .A3(new_n413_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n431_), .B1(new_n430_), .B2(new_n413_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n340_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT20), .ZN(new_n490_));
  INV_X1    g289(.A(new_n423_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n491_), .A2(new_n473_), .A3(new_n467_), .A4(new_n471_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n472_), .A2(KEYINPUT94), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n486_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(new_n482_), .A3(new_n460_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n484_), .A2(new_n485_), .A3(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n482_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(KEYINPUT95), .A3(new_n461_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n351_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n501_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n387_), .A2(new_n351_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G225gat), .A2(G233gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n502_), .A2(new_n503_), .A3(KEYINPUT4), .ZN(new_n508_));
  OR3_X1    g307(.A1(new_n387_), .A2(KEYINPUT4), .A3(new_n351_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n508_), .A2(new_n509_), .A3(new_n505_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G1gat), .B(G29gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(new_n213_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT0), .B(G57gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n512_), .B(new_n513_), .Z(new_n514_));
  NAND3_X1  g313(.A1(new_n507_), .A2(new_n510_), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n514_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n504_), .A2(new_n506_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n505_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n518_));
  OAI221_X1 g317(.A(new_n516_), .B1(KEYINPUT96), .B2(KEYINPUT33), .C1(new_n517_), .C2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n516_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n500_), .A2(new_n515_), .A3(new_n519_), .A4(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT32), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n498_), .B1(new_n524_), .B2(new_n460_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n477_), .A2(new_n463_), .A3(new_n472_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n479_), .A2(KEYINPUT20), .A3(new_n481_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n486_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n526_), .A2(new_n528_), .A3(KEYINPUT32), .A4(new_n461_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n520_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n517_), .A2(new_n518_), .A3(new_n516_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n525_), .B(new_n529_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n456_), .B1(new_n523_), .B2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n530_), .A2(new_n531_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT27), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n497_), .A2(new_n535_), .A3(new_n499_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n526_), .A2(new_n528_), .A3(new_n460_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n484_), .A2(KEYINPUT27), .A3(new_n537_), .ZN(new_n538_));
  AND4_X1   g337(.A1(new_n534_), .A2(new_n456_), .A3(new_n536_), .A4(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n354_), .B1(new_n533_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT97), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n536_), .A2(new_n538_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(new_n456_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n534_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n545_), .A2(new_n354_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(KEYINPUT97), .B(new_n354_), .C1(new_n533_), .C2(new_n539_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n542_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT12), .ZN(new_n550_));
  INV_X1    g349(.A(G57gat), .ZN(new_n551_));
  INV_X1    g350(.A(G64gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G57gat), .A2(G64gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G71gat), .B(G78gat), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT11), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n553_), .A2(new_n559_), .A3(new_n554_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(new_n558_), .A3(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n555_), .A2(new_n557_), .A3(KEYINPUT11), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n561_), .A2(KEYINPUT68), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(KEYINPUT68), .B1(new_n561_), .B2(new_n562_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n550_), .B1(new_n253_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n253_), .A2(new_n565_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G230gat), .A2(G233gat), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n561_), .A2(new_n562_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n263_), .A2(KEYINPUT12), .A3(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n569_), .A2(new_n570_), .A3(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n570_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n567_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n253_), .A2(new_n565_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n574_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G120gat), .B(G148gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(G204gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT5), .B(G176gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n580_), .B(new_n581_), .Z(new_n582_));
  NAND2_X1  g381(.A1(new_n578_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n573_), .A2(new_n577_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT13), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n583_), .A2(KEYINPUT13), .A3(new_n585_), .ZN(new_n589_));
  AND2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G15gat), .B(G22gat), .Z(new_n593_));
  NAND2_X1  g392(.A1(G1gat), .A2(G8gat), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n593_), .B1(KEYINPUT14), .B2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT75), .ZN(new_n596_));
  XOR2_X1   g395(.A(G1gat), .B(G8gat), .Z(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT75), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n595_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n249_), .B1(new_n598_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n598_), .A2(new_n602_), .A3(new_n249_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n604_), .A2(KEYINPUT77), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT77), .B1(new_n604_), .B2(new_n605_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n592_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n605_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n598_), .A2(new_n602_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n264_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n591_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(G113gat), .B(G141gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(new_n408_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT78), .B(G169gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n616_), .B(new_n617_), .Z(new_n618_));
  NAND2_X1  g417(.A1(new_n614_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n618_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n609_), .A2(new_n613_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n590_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n611_), .B(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(new_n571_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G183gat), .B(G211gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(G127gat), .B(G155gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT17), .ZN(new_n632_));
  OAI21_X1  g431(.A(KEYINPUT68), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n626_), .B(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n632_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n623_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n298_), .A2(new_n549_), .A3(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT98), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT99), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(G1gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n545_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n641_), .A2(KEYINPUT38), .A3(new_n642_), .A4(new_n545_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n637_), .B(KEYINPUT100), .Z(new_n647_));
  AND3_X1   g446(.A1(new_n542_), .A2(new_n547_), .A3(new_n548_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n647_), .A2(new_n295_), .A3(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n642_), .B1(new_n649_), .B2(new_n545_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT101), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n645_), .A2(new_n646_), .A3(new_n651_), .ZN(G1324gat));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n649_), .A2(new_n543_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(G8gat), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n655_), .A2(KEYINPUT39), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(KEYINPUT39), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n543_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n659_), .A2(G8gat), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n640_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n653_), .B1(new_n658_), .B2(new_n661_), .ZN(new_n662_));
  OAI221_X1 g461(.A(KEYINPUT40), .B1(new_n640_), .B2(new_n660_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1325gat));
  NOR3_X1   g463(.A1(new_n639_), .A2(G15gat), .A3(new_n354_), .ZN(new_n665_));
  XOR2_X1   g464(.A(new_n665_), .B(KEYINPUT102), .Z(new_n666_));
  INV_X1    g465(.A(new_n354_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n649_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(G15gat), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT41), .Z(new_n670_));
  NAND2_X1  g469(.A1(new_n666_), .A2(new_n670_), .ZN(G1326gat));
  XOR2_X1   g470(.A(new_n456_), .B(KEYINPUT103), .Z(new_n672_));
  NAND2_X1  g471(.A1(new_n649_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(G22gat), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT42), .ZN(new_n675_));
  INV_X1    g474(.A(new_n672_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n676_), .A2(G22gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n675_), .B1(new_n639_), .B2(new_n677_), .ZN(G1327gat));
  INV_X1    g477(.A(G29gat), .ZN(new_n679_));
  INV_X1    g478(.A(new_n636_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n680_), .A2(new_n623_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n549_), .A2(new_n295_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n679_), .B1(new_n683_), .B2(new_n534_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n681_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n549_), .A2(new_n297_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT104), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n297_), .B2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n549_), .B(new_n297_), .C1(new_n688_), .C2(new_n687_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n685_), .B1(new_n690_), .B2(new_n691_), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n692_), .A2(KEYINPUT44), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(G29gat), .A3(new_n545_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n690_), .A2(new_n691_), .ZN(new_n696_));
  AND4_X1   g495(.A1(new_n695_), .A2(new_n696_), .A3(KEYINPUT44), .A4(new_n681_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n695_), .B1(new_n692_), .B2(KEYINPUT44), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n684_), .B1(new_n694_), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT106), .ZN(G1328gat));
  OAI21_X1  g500(.A(KEYINPUT109), .B1(KEYINPUT108), .B2(KEYINPUT46), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706_));
  INV_X1    g505(.A(G36gat), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n682_), .A2(new_n706_), .A3(new_n707_), .A4(new_n543_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT45), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n549_), .A2(new_n707_), .A3(new_n295_), .A4(new_n681_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT107), .B1(new_n710_), .B2(new_n659_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n708_), .A2(new_n709_), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n709_), .B1(new_n708_), .B2(new_n711_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n705_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n543_), .B(new_n693_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n715_));
  AOI211_X1 g514(.A(new_n703_), .B(new_n714_), .C1(G36gat), .C2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(G36gat), .ZN(new_n717_));
  INV_X1    g516(.A(new_n714_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n702_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n716_), .A2(new_n719_), .ZN(G1329gat));
  INV_X1    g519(.A(G43gat), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n354_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n693_), .B(new_n722_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n721_), .B1(new_n683_), .B2(new_n354_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g525(.A1(new_n683_), .A2(G50gat), .A3(new_n676_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n456_), .B(new_n693_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n728_), .A2(new_n729_), .A3(G50gat), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n729_), .B1(new_n728_), .B2(G50gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1331gat));
  INV_X1    g531(.A(new_n590_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n636_), .A2(new_n622_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n549_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(new_n284_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n736_), .A2(KEYINPUT112), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(KEYINPUT112), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n545_), .A3(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(G57gat), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n735_), .A2(new_n298_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n742_), .A2(KEYINPUT111), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(KEYINPUT111), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n743_), .A2(new_n551_), .A3(new_n545_), .A4(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT113), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n740_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n740_), .B2(new_n745_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1332gat));
  NAND3_X1  g548(.A1(new_n737_), .A2(new_n543_), .A3(new_n738_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT48), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(G64gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n750_), .B2(G64gat), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n743_), .A2(new_n744_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n543_), .A2(new_n552_), .ZN(new_n755_));
  OAI22_X1  g554(.A1(new_n752_), .A2(new_n753_), .B1(new_n754_), .B2(new_n755_), .ZN(G1333gat));
  NAND3_X1  g555(.A1(new_n737_), .A2(new_n667_), .A3(new_n738_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT49), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n757_), .A2(new_n758_), .A3(G71gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n757_), .B2(G71gat), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n354_), .A2(G71gat), .ZN(new_n761_));
  OAI22_X1  g560(.A1(new_n759_), .A2(new_n760_), .B1(new_n754_), .B2(new_n761_), .ZN(G1334gat));
  NAND3_X1  g561(.A1(new_n737_), .A2(new_n672_), .A3(new_n738_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT50), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(G78gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G78gat), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n676_), .A2(G78gat), .ZN(new_n767_));
  OAI22_X1  g566(.A1(new_n765_), .A2(new_n766_), .B1(new_n754_), .B2(new_n767_), .ZN(G1335gat));
  NOR3_X1   g567(.A1(new_n680_), .A2(new_n590_), .A3(new_n622_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n549_), .A2(new_n295_), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(G85gat), .B1(new_n770_), .B2(new_n545_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n696_), .A2(new_n769_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n534_), .B1(new_n208_), .B2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n771_), .B1(new_n773_), .B2(new_n775_), .ZN(G1336gat));
  AOI21_X1  g575(.A(G92gat), .B1(new_n770_), .B2(new_n543_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n659_), .A2(new_n211_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n773_), .B2(new_n778_), .ZN(G1337gat));
  OAI21_X1  g578(.A(G99gat), .B1(new_n772_), .B2(new_n354_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n770_), .B(new_n667_), .C1(new_n227_), .C2(new_n226_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT114), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n781_), .A2(new_n782_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n780_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n785_), .B(new_n786_), .Z(G1338gat));
  AND3_X1   g586(.A1(new_n696_), .A2(new_n456_), .A3(new_n769_), .ZN(new_n788_));
  OAI21_X1  g587(.A(KEYINPUT116), .B1(new_n788_), .B2(new_n223_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT116), .ZN(new_n790_));
  INV_X1    g589(.A(new_n456_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n790_), .B(G106gat), .C1(new_n772_), .C2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(KEYINPUT52), .A3(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n770_), .A2(new_n223_), .A3(new_n456_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795_));
  OAI211_X1 g594(.A(KEYINPUT116), .B(new_n795_), .C1(new_n788_), .C2(new_n223_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(new_n794_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT53), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n793_), .A2(new_n799_), .A3(new_n794_), .A4(new_n796_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1339gat));
  NAND3_X1  g600(.A1(new_n544_), .A2(new_n545_), .A3(new_n667_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT117), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n290_), .A2(new_n296_), .A3(new_n734_), .A4(new_n590_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  INV_X1    g606(.A(new_n585_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n263_), .A2(KEYINPUT12), .A3(new_n571_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n574_), .B1(new_n568_), .B2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT55), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n573_), .ZN(new_n812_));
  AND4_X1   g611(.A1(new_n570_), .A2(new_n572_), .A3(new_n566_), .A4(new_n567_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n810_), .A2(new_n813_), .A3(KEYINPUT55), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n812_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(KEYINPUT56), .A3(new_n582_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n813_), .B1(new_n810_), .B2(KEYINPUT55), .ZN(new_n817_));
  AND4_X1   g616(.A1(KEYINPUT55), .A2(new_n569_), .A3(new_n570_), .A4(new_n572_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n582_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n808_), .B1(new_n816_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n591_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n612_), .A2(new_n592_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n618_), .A3(new_n824_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n621_), .A2(new_n825_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n822_), .A2(new_n622_), .B1(new_n586_), .B2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n807_), .B1(new_n827_), .B2(new_n295_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n586_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT56), .B1(new_n815_), .B2(new_n582_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n819_), .A2(new_n820_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n585_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n622_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n829_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(KEYINPUT57), .A3(new_n284_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n828_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n621_), .A2(new_n825_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n832_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n822_), .A2(KEYINPUT58), .A3(new_n826_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n297_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n680_), .B1(new_n836_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n803_), .B1(new_n806_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G113gat), .B1(new_n844_), .B2(new_n622_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n804_), .B(KEYINPUT54), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n839_), .A2(new_n840_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n848_), .B1(new_n290_), .B2(new_n296_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n828_), .A2(new_n835_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n636_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n847_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT59), .B1(new_n852_), .B2(new_n803_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT59), .ZN(new_n854_));
  INV_X1    g653(.A(new_n803_), .ZN(new_n855_));
  AOI211_X1 g654(.A(new_n854_), .B(new_n855_), .C1(new_n847_), .C2(new_n851_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n846_), .B1(new_n853_), .B2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n843_), .A2(new_n854_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n852_), .A2(KEYINPUT59), .A3(new_n803_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(KEYINPUT118), .A3(new_n859_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n857_), .A2(new_n860_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n622_), .A2(G113gat), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n845_), .B1(new_n861_), .B2(new_n862_), .ZN(G1340gat));
  NOR2_X1   g662(.A1(new_n590_), .A2(G120gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n844_), .B1(KEYINPUT60), .B2(new_n864_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n865_), .B(new_n733_), .C1(new_n853_), .C2(new_n856_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(G120gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(KEYINPUT60), .B2(new_n865_), .ZN(G1341gat));
  INV_X1    g667(.A(G127gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n636_), .A2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n857_), .A2(new_n860_), .A3(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n869_), .B1(new_n843_), .B2(new_n636_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT119), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT119), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n871_), .A2(new_n875_), .A3(new_n872_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(G1342gat));
  AOI21_X1  g676(.A(G134gat), .B1(new_n844_), .B2(new_n295_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n297_), .A2(G134gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT120), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n861_), .B2(new_n880_), .ZN(G1343gat));
  NAND4_X1  g680(.A1(new_n659_), .A2(new_n545_), .A3(new_n456_), .A4(new_n354_), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n882_), .B(KEYINPUT121), .Z(new_n883_));
  AOI21_X1  g682(.A(new_n883_), .B1(new_n847_), .B2(new_n851_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n622_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n733_), .ZN(new_n887_));
  XOR2_X1   g686(.A(KEYINPUT122), .B(G148gat), .Z(new_n888_));
  XNOR2_X1  g687(.A(new_n887_), .B(new_n888_), .ZN(G1345gat));
  NAND2_X1  g688(.A1(new_n884_), .A2(new_n680_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  AOI21_X1  g691(.A(G162gat), .B1(new_n884_), .B2(new_n295_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT123), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n298_), .A2(new_n356_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n884_), .B2(new_n895_), .ZN(G1347gat));
  NAND3_X1  g695(.A1(new_n852_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n897_), .A2(new_n833_), .A3(new_n672_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT62), .ZN(new_n899_));
  OR3_X1    g698(.A1(new_n898_), .A2(new_n899_), .A3(new_n306_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n464_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n899_), .B1(new_n898_), .B2(new_n306_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(G1348gat));
  NOR2_X1   g702(.A1(new_n897_), .A2(new_n672_), .ZN(new_n904_));
  AOI21_X1  g703(.A(G176gat), .B1(new_n904_), .B2(new_n733_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n897_), .A2(new_n456_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n590_), .A2(new_n307_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(G1349gat));
  OAI211_X1 g707(.A(new_n904_), .B(new_n680_), .C1(new_n320_), .C2(new_n322_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT124), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n909_), .A2(new_n910_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G183gat), .B1(new_n906_), .B2(new_n680_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n911_), .A2(new_n912_), .A3(new_n913_), .ZN(G1350gat));
  AND2_X1   g713(.A1(new_n295_), .A2(new_n299_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n904_), .A2(new_n915_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n897_), .A2(new_n298_), .A3(new_n672_), .ZN(new_n917_));
  INV_X1    g716(.A(G190gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n916_), .B1(new_n917_), .B2(new_n918_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(KEYINPUT125), .ZN(G1351gat));
  NOR3_X1   g719(.A1(new_n667_), .A2(new_n791_), .A3(new_n545_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n852_), .A2(new_n543_), .A3(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n852_), .A2(KEYINPUT126), .A3(new_n543_), .A4(new_n921_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n622_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n733_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  NAND2_X1  g730(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n932_));
  AND4_X1   g731(.A1(new_n680_), .A2(new_n926_), .A3(new_n931_), .A4(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n931_), .B1(new_n926_), .B2(new_n680_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1354gat));
  AOI21_X1  g734(.A(new_n405_), .B1(new_n926_), .B2(new_n297_), .ZN(new_n936_));
  AOI211_X1 g735(.A(G218gat), .B(new_n284_), .C1(new_n924_), .C2(new_n925_), .ZN(new_n937_));
  OAI21_X1  g736(.A(KEYINPUT127), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n926_), .A2(new_n405_), .A3(new_n295_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n298_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n939_), .B(new_n940_), .C1(new_n405_), .C2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n938_), .A2(new_n942_), .ZN(G1355gat));
endmodule


