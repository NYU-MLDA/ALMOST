//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n940_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n954_, new_n955_, new_n957_, new_n958_, new_n959_,
    new_n961_, new_n962_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n970_, new_n971_, new_n972_, new_n974_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_;
  NAND2_X1  g000(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n202_));
  OR2_X1    g001(.A1(KEYINPUT74), .A2(KEYINPUT13), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT64), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT64), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n210_));
  AND3_X1   g009(.A1(new_n206_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n206_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n204_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n208_), .A2(new_n210_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(new_n205_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n206_), .A2(new_n208_), .A3(new_n210_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(KEYINPUT65), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT10), .B(G99gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G106gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT9), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(G85gat), .A3(G92gat), .ZN(new_n224_));
  XOR2_X1   g023(.A(G85gat), .B(G92gat), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT9), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n218_), .A2(new_n222_), .A3(new_n224_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n230_));
  NAND2_X1  g029(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n231_));
  INV_X1    g030(.A(G99gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(new_n232_), .A3(new_n221_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n230_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n236_));
  OR2_X1    g035(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n237_));
  NOR2_X1   g036(.A1(G99gat), .A2(G106gat), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n237_), .A2(KEYINPUT67), .A3(new_n238_), .A4(new_n231_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n235_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n215_), .A2(new_n216_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n225_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n229_), .B1(new_n242_), .B2(KEYINPUT8), .ZN(new_n243_));
  INV_X1    g042(.A(new_n225_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n244_), .A2(KEYINPUT8), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n240_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n246_), .B1(new_n218_), .B2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n243_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n242_), .A2(new_n229_), .A3(KEYINPUT8), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n228_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G57gat), .B(G64gat), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n252_), .A2(KEYINPUT11), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(KEYINPUT11), .ZN(new_n254_));
  XOR2_X1   g053(.A(G71gat), .B(G78gat), .Z(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n254_), .A2(new_n255_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT12), .B1(new_n251_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n242_), .A2(KEYINPUT8), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT68), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n218_), .A2(new_n247_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(new_n245_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n250_), .A3(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n227_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT12), .ZN(new_n266_));
  INV_X1    g065(.A(new_n258_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n259_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n264_), .A2(new_n258_), .A3(new_n227_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G230gat), .A2(G233gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT70), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n270_), .A2(KEYINPUT70), .A3(new_n271_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n269_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n265_), .A2(new_n267_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(KEYINPUT69), .A3(new_n270_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n271_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n265_), .A2(new_n280_), .A3(new_n267_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n278_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G176gat), .B(G204gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT72), .ZN(new_n284_));
  XOR2_X1   g083(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G120gat), .B(G148gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n286_), .B(new_n287_), .Z(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n276_), .A2(new_n282_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n289_), .B1(new_n276_), .B2(new_n282_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n293_));
  NOR3_X1   g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n276_), .A2(new_n282_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n288_), .ZN(new_n296_));
  AOI21_X1  g095(.A(KEYINPUT73), .B1(new_n296_), .B2(new_n290_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n202_), .B(new_n203_), .C1(new_n294_), .C2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n293_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n296_), .A2(KEYINPUT73), .A3(new_n290_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(KEYINPUT74), .A4(KEYINPUT13), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n298_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G8gat), .B(G36gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT18), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G64gat), .B(G92gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT20), .ZN(new_n307_));
  NOR2_X1   g106(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n308_));
  INV_X1    g107(.A(G169gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT23), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n311_), .A2(G183gat), .A3(G190gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT88), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT88), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n314_), .A2(new_n311_), .A3(G183gat), .A4(G190gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G183gat), .A2(G190gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT87), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n316_), .A2(new_n317_), .A3(KEYINPUT23), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n316_), .B2(KEYINPUT23), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n313_), .B(new_n315_), .C1(new_n318_), .C2(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n310_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT25), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n324_), .A2(G183gat), .ZN(new_n325_));
  INV_X1    g124(.A(G183gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n326_), .A2(KEYINPUT25), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT98), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT26), .B(G190gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n326_), .A2(KEYINPUT25), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(G183gat), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT98), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n328_), .A2(new_n329_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G176gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n309_), .A2(new_n335_), .A3(KEYINPUT86), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT86), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(G169gat), .B2(G176gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT24), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n316_), .A2(KEYINPUT23), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n312_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n340_), .B1(G169gat), .B2(G176gat), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n343_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n323_), .B1(new_n334_), .B2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G197gat), .A2(G204gat), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G197gat), .A2(G204gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(KEYINPUT21), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT21), .ZN(new_n353_));
  INV_X1    g152(.A(new_n351_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n353_), .B1(new_n354_), .B2(new_n349_), .ZN(new_n355_));
  INV_X1    g154(.A(G211gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(G218gat), .ZN(new_n357_));
  INV_X1    g156(.A(G218gat), .ZN(new_n358_));
  AOI21_X1  g157(.A(KEYINPUT96), .B1(new_n358_), .B2(G211gat), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n352_), .A2(new_n355_), .A3(new_n357_), .A4(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n357_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n361_), .A2(KEYINPUT21), .A3(new_n350_), .A4(new_n351_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n307_), .B1(new_n348_), .B2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n329_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n320_), .A2(new_n341_), .A3(new_n345_), .A4(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n310_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n343_), .A2(new_n322_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT99), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n360_), .A2(new_n362_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n371_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n364_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT19), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n376_), .A2(KEYINPUT101), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n334_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n380_), .A2(new_n346_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n372_), .B1(new_n381_), .B2(new_n323_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n378_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n363_), .A2(new_n369_), .A3(new_n366_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n382_), .A2(KEYINPUT20), .A3(new_n383_), .A4(new_n384_), .ZN(new_n385_));
  AOI22_X1  g184(.A1(new_n376_), .A2(new_n378_), .B1(KEYINPUT101), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n306_), .B1(new_n379_), .B2(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n364_), .B(new_n383_), .C1(new_n374_), .C2(new_n375_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n306_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n382_), .A2(KEYINPUT20), .A3(new_n384_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n378_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n387_), .A2(KEYINPUT103), .A3(KEYINPUT27), .A4(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT103), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n385_), .A2(KEYINPUT101), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n320_), .A2(new_n322_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n367_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n334_), .A2(new_n343_), .A3(new_n341_), .A4(new_n345_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n363_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT20), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n370_), .A2(new_n372_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT99), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n400_), .B1(new_n402_), .B2(new_n373_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n395_), .B1(new_n403_), .B2(new_n383_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n376_), .A2(KEYINPUT101), .A3(new_n378_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n389_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n392_), .A2(KEYINPUT27), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n394_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n388_), .A2(new_n391_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n306_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n392_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT27), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n393_), .A2(new_n408_), .A3(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G78gat), .B(G106gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT94), .B(G228gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT95), .B(G233gat), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT3), .ZN(new_n421_));
  INV_X1    g220(.A(G141gat), .ZN(new_n422_));
  INV_X1    g221(.A(G148gat), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(new_n422_), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G141gat), .A2(G148gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT2), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n424_), .A2(new_n427_), .A3(new_n428_), .A4(new_n429_), .ZN(new_n430_));
  OR2_X1    g229(.A1(G155gat), .A2(G162gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G155gat), .A2(G162gat), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(KEYINPUT1), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT1), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(G155gat), .A3(G162gat), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n437_), .A3(new_n431_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G141gat), .B(G148gat), .Z(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n434_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT29), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n420_), .B1(new_n442_), .B2(new_n372_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n372_), .A3(new_n420_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n416_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT97), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G22gat), .B(G50gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT29), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n434_), .A2(new_n440_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT91), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n430_), .A2(new_n433_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(KEYINPUT91), .A3(new_n451_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT93), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n454_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n457_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n450_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n454_), .A2(new_n456_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT93), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n454_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n449_), .A3(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n460_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n465_), .B1(new_n460_), .B2(new_n464_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n448_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n444_), .A2(new_n445_), .A3(new_n416_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n469_), .A2(new_n446_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n470_), .B(new_n448_), .C1(new_n466_), .C2(new_n467_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n414_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT89), .ZN(new_n477_));
  INV_X1    g276(.A(G134gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(G127gat), .ZN(new_n479_));
  INV_X1    g278(.A(G127gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(G134gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(G120gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(G113gat), .ZN(new_n484_));
  INV_X1    g283(.A(G113gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(G120gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n477_), .B1(new_n482_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n482_), .A2(new_n487_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n479_), .A2(new_n481_), .A3(new_n484_), .A4(new_n486_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n488_), .B1(new_n491_), .B2(new_n477_), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n492_), .B(KEYINPUT31), .Z(new_n493_));
  INV_X1    g292(.A(KEYINPUT90), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G227gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(G15gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT30), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G71gat), .B(G99gat), .ZN(new_n500_));
  INV_X1    g299(.A(G43gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n499_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(new_n370_), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n495_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n494_), .A3(new_n493_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G1gat), .B(G29gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(G85gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT0), .B(G57gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n482_), .A2(new_n487_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n479_), .A2(new_n481_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n477_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n488_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n441_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n455_), .A2(new_n491_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(KEYINPUT4), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT4), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n514_), .A2(new_n441_), .A3(new_n519_), .A4(new_n515_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT100), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT100), .ZN(new_n522_));
  NAND4_X1  g321(.A1(new_n492_), .A2(new_n522_), .A3(new_n519_), .A4(new_n441_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n518_), .A2(new_n521_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G225gat), .A2(G233gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n526_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n511_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n511_), .ZN(new_n531_));
  AOI211_X1 g330(.A(new_n531_), .B(new_n528_), .C1(new_n524_), .C2(new_n526_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n507_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n476_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n472_), .A2(new_n473_), .A3(new_n533_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n414_), .A2(new_n537_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n518_), .A2(new_n521_), .A3(new_n523_), .A4(new_n525_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n516_), .A2(new_n526_), .A3(new_n517_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n540_), .A2(new_n511_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT33), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n528_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n544_));
  OAI22_X1  g343(.A1(new_n542_), .A2(new_n543_), .B1(new_n544_), .B2(new_n511_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n527_), .A2(new_n529_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(KEYINPUT33), .A3(new_n531_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n389_), .A2(KEYINPUT32), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n388_), .A2(new_n391_), .A3(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n550_), .B1(new_n530_), .B2(new_n532_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n549_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n552_));
  OAI22_X1  g351(.A1(new_n548_), .A2(new_n411_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT102), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n474_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n553_), .B2(new_n474_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n538_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n507_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n536_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G15gat), .B(G22gat), .Z(new_n561_));
  NAND2_X1  g360(.A1(G1gat), .A2(G8gat), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(KEYINPUT14), .B2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT81), .ZN(new_n564_));
  XOR2_X1   g363(.A(G1gat), .B(G8gat), .Z(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT81), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n563_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n565_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G29gat), .B(G36gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G43gat), .B(G50gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n566_), .A2(new_n570_), .A3(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n574_), .A2(KEYINPUT84), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(KEYINPUT84), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G229gat), .A2(G233gat), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n566_), .A2(new_n570_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n573_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n577_), .A2(new_n579_), .A3(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n573_), .B(KEYINPUT15), .ZN(new_n584_));
  AOI22_X1  g383(.A1(new_n575_), .A2(new_n576_), .B1(new_n580_), .B2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n583_), .B1(new_n579_), .B2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G113gat), .B(G141gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT85), .ZN(new_n588_));
  XOR2_X1   g387(.A(G169gat), .B(G197gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  OR2_X1    g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n590_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(KEYINPUT104), .B1(new_n560_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT104), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n559_), .A2(new_n596_), .A3(new_n593_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n302_), .B1(new_n595_), .B2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n258_), .B(new_n599_), .Z(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(new_n580_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G127gat), .B(G155gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT16), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT17), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n601_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(KEYINPUT17), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT82), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n601_), .A2(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT83), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(KEYINPUT83), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n607_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT34), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT35), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n251_), .A2(new_n573_), .B1(new_n618_), .B2(new_n617_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT75), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n622_), .B1(new_n265_), .B2(new_n584_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n584_), .ZN(new_n624_));
  AOI211_X1 g423(.A(KEYINPUT75), .B(new_n624_), .C1(new_n264_), .C2(new_n227_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n620_), .B(new_n621_), .C1(new_n623_), .C2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n264_), .A2(new_n573_), .A3(new_n227_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n617_), .A2(new_n618_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT75), .B1(new_n251_), .B2(new_n624_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n265_), .A2(new_n622_), .A3(new_n584_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n629_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n632_), .A2(KEYINPUT76), .A3(new_n620_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT76), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n621_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n635_), .B2(new_n619_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n626_), .B1(new_n633_), .B2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G190gat), .B(G218gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G134gat), .B(G162gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT36), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n637_), .A2(KEYINPUT79), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT79), .ZN(new_n644_));
  INV_X1    g443(.A(new_n626_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT76), .B1(new_n632_), .B2(new_n620_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n635_), .A2(new_n634_), .A3(new_n619_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n645_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n644_), .B1(new_n648_), .B2(new_n641_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n647_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT78), .ZN(new_n651_));
  XOR2_X1   g450(.A(KEYINPUT77), .B(KEYINPUT36), .Z(new_n652_));
  NOR2_X1   g451(.A1(new_n640_), .A2(new_n652_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n626_), .A2(new_n653_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n650_), .A2(new_n651_), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n651_), .B1(new_n650_), .B2(new_n654_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n643_), .B(new_n649_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(KEYINPUT37), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n641_), .B1(new_n650_), .B2(new_n626_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n654_), .B1(new_n633_), .B2(new_n636_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT78), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n650_), .A2(new_n651_), .A3(new_n654_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(KEYINPUT80), .B(KEYINPUT37), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n614_), .B1(new_n658_), .B2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n598_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(G1gat), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(new_n534_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT38), .ZN(new_n670_));
  OR2_X1    g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n302_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n593_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n663_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n559_), .A2(new_n613_), .A3(new_n674_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G1gat), .B1(new_n677_), .B2(new_n533_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n669_), .A2(new_n670_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n671_), .A2(new_n678_), .A3(new_n679_), .ZN(G1324gat));
  INV_X1    g479(.A(new_n414_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n681_), .A2(G8gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n667_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT105), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT105), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n667_), .A2(new_n685_), .A3(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G8gat), .B1(new_n677_), .B2(new_n681_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT39), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT40), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n687_), .A2(KEYINPUT40), .A3(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1325gat));
  NAND3_X1  g493(.A1(new_n667_), .A2(new_n497_), .A3(new_n558_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n497_), .B1(new_n676_), .B2(new_n558_), .ZN(new_n696_));
  XOR2_X1   g495(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n697_));
  OR2_X1    g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n697_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n695_), .A2(new_n698_), .A3(new_n699_), .ZN(G1326gat));
  INV_X1    g499(.A(G22gat), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n676_), .B2(new_n475_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT42), .Z(new_n703_));
  NAND3_X1  g502(.A1(new_n667_), .A2(new_n701_), .A3(new_n475_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(G1327gat));
  NAND2_X1  g504(.A1(new_n663_), .A2(new_n614_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n598_), .A2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G29gat), .B1(new_n708_), .B2(new_n534_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n559_), .A2(new_n658_), .A3(new_n665_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT43), .ZN(new_n711_));
  AOI22_X1  g510(.A1(new_n657_), .A2(KEYINPUT37), .B1(new_n663_), .B2(new_n664_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n712_), .A2(new_n713_), .A3(new_n559_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n302_), .A2(new_n613_), .A3(new_n594_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT44), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  AND4_X1   g516(.A1(new_n713_), .A2(new_n559_), .A3(new_n658_), .A4(new_n665_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n713_), .B1(new_n712_), .B2(new_n559_), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT44), .B(new_n716_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n715_), .A2(KEYINPUT107), .A3(KEYINPUT44), .A4(new_n716_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n717_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n534_), .A2(G29gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n709_), .B1(new_n724_), .B2(new_n725_), .ZN(G1328gat));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n414_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G36gat), .ZN(new_n728_));
  INV_X1    g527(.A(G36gat), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n414_), .A2(KEYINPUT108), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n414_), .A2(KEYINPUT108), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n598_), .A2(new_n729_), .A3(new_n707_), .A4(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n733_), .B(new_n734_), .Z(new_n735_));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n728_), .A2(new_n735_), .A3(KEYINPUT110), .A4(new_n736_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n736_), .A2(KEYINPUT110), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(KEYINPUT110), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n729_), .B1(new_n724_), .B2(new_n414_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n733_), .B(new_n734_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n738_), .B(new_n739_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n737_), .A2(new_n742_), .ZN(G1329gat));
  NAND3_X1  g542(.A1(new_n598_), .A2(new_n558_), .A3(new_n707_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n501_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT112), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n744_), .A2(KEYINPUT112), .A3(new_n501_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n722_), .A2(new_n723_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n717_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n507_), .A2(new_n501_), .ZN(new_n752_));
  AND4_X1   g551(.A1(KEYINPUT111), .A2(new_n750_), .A3(new_n751_), .A4(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT111), .B1(new_n724_), .B2(new_n752_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n749_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT47), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT47), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(new_n749_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1330gat));
  INV_X1    g558(.A(G50gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n708_), .A2(new_n760_), .A3(new_n475_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n724_), .A2(KEYINPUT113), .A3(new_n475_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G50gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT113), .B1(new_n724_), .B2(new_n475_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n763_), .B2(new_n764_), .ZN(G1331gat));
  NOR2_X1   g564(.A1(new_n672_), .A2(new_n593_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n767_), .A2(new_n560_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n768_), .A2(new_n666_), .ZN(new_n769_));
  INV_X1    g568(.A(G57gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n534_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n767_), .A2(new_n675_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G57gat), .B1(new_n773_), .B2(new_n533_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n771_), .A2(new_n774_), .ZN(G1332gat));
  INV_X1    g574(.A(G64gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n769_), .A2(new_n776_), .A3(new_n732_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n772_), .B2(new_n732_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n778_), .A2(new_n779_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n777_), .B1(new_n780_), .B2(new_n781_), .ZN(G1333gat));
  INV_X1    g581(.A(G71gat), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n769_), .A2(new_n783_), .A3(new_n558_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n772_), .A2(new_n558_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(G71gat), .ZN(new_n787_));
  AOI211_X1 g586(.A(KEYINPUT49), .B(new_n783_), .C1(new_n772_), .C2(new_n558_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  XOR2_X1   g588(.A(new_n789_), .B(KEYINPUT115), .Z(G1334gat));
  INV_X1    g589(.A(G78gat), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n769_), .A2(new_n791_), .A3(new_n475_), .ZN(new_n792_));
  OAI21_X1  g591(.A(G78gat), .B1(new_n773_), .B2(new_n474_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(KEYINPUT50), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(KEYINPUT50), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n792_), .B1(new_n794_), .B2(new_n795_), .ZN(G1335gat));
  NAND3_X1  g595(.A1(new_n715_), .A2(new_n614_), .A3(new_n766_), .ZN(new_n797_));
  OAI21_X1  g596(.A(G85gat), .B1(new_n797_), .B2(new_n533_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n768_), .A2(new_n707_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n533_), .A2(G85gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n798_), .B1(new_n799_), .B2(new_n800_), .ZN(G1336gat));
  INV_X1    g600(.A(new_n732_), .ZN(new_n802_));
  OAI21_X1  g601(.A(G92gat), .B1(new_n797_), .B2(new_n802_), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n681_), .A2(G92gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n799_), .B2(new_n804_), .ZN(G1337gat));
  OAI21_X1  g604(.A(G99gat), .B1(new_n797_), .B2(new_n507_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n558_), .A2(new_n220_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n799_), .B2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT51), .ZN(G1338gat));
  OR2_X1    g608(.A1(new_n797_), .A2(new_n474_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n810_), .A2(new_n811_), .A3(G106gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n810_), .B2(G106gat), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n475_), .A2(new_n221_), .ZN(new_n814_));
  OAI22_X1  g613(.A1(new_n812_), .A2(new_n813_), .B1(new_n799_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT53), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817_));
  OAI221_X1 g616(.A(new_n817_), .B1(new_n799_), .B2(new_n814_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1339gat));
  NAND2_X1  g618(.A1(new_n593_), .A2(G113gat), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(KEYINPUT120), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n266_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n823_));
  AOI211_X1 g622(.A(KEYINPUT12), .B(new_n258_), .C1(new_n264_), .C2(new_n227_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n270_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n279_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n269_), .A2(new_n274_), .A3(KEYINPUT55), .A4(new_n275_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n275_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT70), .B1(new_n270_), .B2(new_n271_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n829_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT117), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n276_), .A2(new_n834_), .A3(new_n829_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n828_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n822_), .B1(new_n836_), .B2(new_n289_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n289_), .A2(new_n822_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n838_), .B1(new_n836_), .B2(new_n840_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n276_), .A2(new_n834_), .A3(new_n829_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n834_), .B1(new_n276_), .B2(new_n829_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n827_), .B(new_n826_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(KEYINPUT118), .A3(new_n839_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n837_), .A2(new_n841_), .A3(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n594_), .A2(new_n291_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n577_), .A2(new_n582_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n590_), .B1(new_n849_), .B2(new_n578_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n585_), .A2(new_n579_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n592_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n848_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n663_), .A2(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(KEYINPUT119), .A3(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n854_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n857_), .B1(new_n860_), .B2(new_n663_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT119), .ZN(new_n862_));
  INV_X1    g661(.A(new_n858_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n860_), .B2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n853_), .A2(new_n291_), .ZN(new_n865_));
  AOI21_X1  g664(.A(KEYINPUT56), .B1(new_n844_), .B2(new_n288_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n836_), .A2(new_n840_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OAI211_X1 g669(.A(KEYINPUT58), .B(new_n865_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n870_), .A2(new_n712_), .A3(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n859_), .A2(new_n861_), .A3(new_n864_), .A4(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n614_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n593_), .B1(KEYINPUT116), .B2(KEYINPUT54), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n298_), .A2(new_n876_), .A3(new_n301_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n875_), .B1(new_n666_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n875_), .ZN(new_n880_));
  NOR4_X1   g679(.A1(new_n712_), .A2(new_n877_), .A3(new_n614_), .A4(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n879_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n874_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n476_), .A2(new_n534_), .A3(new_n558_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(KEYINPUT59), .B1(new_n884_), .B2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n882_), .B1(new_n873_), .B2(new_n614_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n888_), .A2(new_n889_), .A3(new_n885_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n821_), .B1(new_n887_), .B2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n884_), .A2(new_n886_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n485_), .B1(new_n892_), .B2(new_n594_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n891_), .A2(KEYINPUT121), .A3(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT121), .ZN(new_n895_));
  INV_X1    g694(.A(new_n821_), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT119), .B1(new_n856_), .B2(new_n858_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n860_), .A2(new_n863_), .A3(new_n862_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n861_), .A2(new_n872_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n613_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  OAI211_X1 g700(.A(KEYINPUT59), .B(new_n886_), .C1(new_n901_), .C2(new_n882_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n889_), .B1(new_n888_), .B2(new_n885_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n896_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n888_), .A2(new_n885_), .ZN(new_n905_));
  AOI21_X1  g704(.A(G113gat), .B1(new_n905_), .B2(new_n593_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n895_), .B1(new_n904_), .B2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n894_), .A2(new_n907_), .ZN(G1340gat));
  AOI21_X1  g707(.A(new_n672_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n483_), .B1(new_n672_), .B2(KEYINPUT60), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n910_), .B1(KEYINPUT60), .B2(new_n483_), .ZN(new_n911_));
  OAI22_X1  g710(.A1(new_n909_), .A2(new_n483_), .B1(new_n892_), .B2(new_n911_), .ZN(G1341gat));
  NAND3_X1  g711(.A1(new_n905_), .A2(new_n480_), .A3(new_n613_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n614_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n480_), .ZN(G1342gat));
  NAND3_X1  g714(.A1(new_n905_), .A2(new_n478_), .A3(new_n663_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n712_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n916_), .B1(new_n918_), .B2(new_n478_), .ZN(G1343gat));
  NOR3_X1   g718(.A1(new_n474_), .A2(new_n558_), .A3(new_n533_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n802_), .A2(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n874_), .B2(new_n883_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n593_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n302_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g725(.A(KEYINPUT61), .B(G155gat), .ZN(new_n927_));
  INV_X1    g726(.A(new_n921_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n884_), .A2(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(KEYINPUT122), .B1(new_n929_), .B2(new_n614_), .ZN(new_n930_));
  NOR4_X1   g729(.A1(new_n888_), .A2(KEYINPUT122), .A3(new_n614_), .A4(new_n921_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n931_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n927_), .B1(new_n930_), .B2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n934_), .B1(new_n922_), .B2(new_n613_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n927_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n935_), .A2(new_n931_), .A3(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n933_), .A2(new_n937_), .ZN(G1346gat));
  OR3_X1    g737(.A1(new_n929_), .A2(G162gat), .A3(new_n674_), .ZN(new_n939_));
  OAI21_X1  g738(.A(G162gat), .B1(new_n929_), .B2(new_n917_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1347gat));
  INV_X1    g740(.A(KEYINPUT22), .ZN(new_n942_));
  NAND3_X1  g741(.A1(new_n732_), .A2(new_n474_), .A3(new_n535_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n943_), .ZN(new_n944_));
  NAND4_X1  g743(.A1(new_n884_), .A2(new_n942_), .A3(new_n593_), .A4(new_n944_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  NAND3_X1  g746(.A1(new_n945_), .A2(new_n309_), .A3(new_n947_), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n945_), .A2(new_n947_), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n884_), .A2(new_n593_), .A3(new_n946_), .A4(new_n944_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(G169gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n948_), .B1(new_n949_), .B2(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(G1348gat));
  NAND2_X1  g752(.A1(new_n884_), .A2(new_n944_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n954_), .A2(new_n672_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(new_n335_), .ZN(G1349gat));
  NOR2_X1   g755(.A1(new_n954_), .A2(new_n614_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n957_), .A2(G183gat), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n328_), .A2(new_n333_), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n958_), .B1(new_n959_), .B2(new_n957_), .ZN(G1350gat));
  OAI21_X1  g759(.A(G190gat), .B1(new_n954_), .B2(new_n917_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n663_), .A2(new_n329_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n961_), .B1(new_n954_), .B2(new_n962_), .ZN(G1351gat));
  NOR2_X1   g762(.A1(new_n537_), .A2(new_n558_), .ZN(new_n964_));
  XOR2_X1   g763(.A(new_n964_), .B(KEYINPUT124), .Z(new_n965_));
  NOR3_X1   g764(.A1(new_n888_), .A2(new_n802_), .A3(new_n965_), .ZN(new_n966_));
  INV_X1    g765(.A(G197gat), .ZN(new_n967_));
  OR2_X1    g766(.A1(new_n967_), .A2(KEYINPUT125), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n967_), .A2(KEYINPUT125), .ZN(new_n969_));
  AOI22_X1  g768(.A1(new_n966_), .A2(new_n593_), .B1(new_n968_), .B2(new_n969_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n966_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n971_), .A2(new_n594_), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n970_), .B1(new_n972_), .B2(new_n969_), .ZN(G1352gat));
  NAND2_X1  g772(.A1(new_n966_), .A2(new_n302_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g774(.A(new_n614_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n966_), .A2(new_n976_), .ZN(new_n977_));
  NOR2_X1   g776(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n978_));
  XOR2_X1   g777(.A(new_n978_), .B(KEYINPUT126), .Z(new_n979_));
  XOR2_X1   g778(.A(new_n979_), .B(KEYINPUT127), .Z(new_n980_));
  INV_X1    g779(.A(new_n980_), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n977_), .B(new_n981_), .ZN(G1354gat));
  OAI21_X1  g781(.A(G218gat), .B1(new_n971_), .B2(new_n917_), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n966_), .A2(new_n358_), .A3(new_n663_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n983_), .A2(new_n984_), .ZN(G1355gat));
endmodule


