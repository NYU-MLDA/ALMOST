//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT20), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT24), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT89), .B1(G169gat), .B2(G176gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR3_X1   g007(.A1(KEYINPUT89), .A2(G169gat), .A3(G176gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n206_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT90), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n210_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT89), .ZN(new_n219_));
  INV_X1    g018(.A(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT24), .B1(new_n222_), .B2(new_n207_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT90), .B1(new_n223_), .B2(new_n215_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT25), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G183gat), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n226_), .A2(KEYINPUT88), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT26), .B(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n226_), .A2(KEYINPUT88), .ZN(new_n229_));
  INV_X1    g028(.A(G183gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT25), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .A4(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n222_), .A2(KEYINPUT24), .A3(new_n207_), .A4(new_n233_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n218_), .A2(new_n224_), .A3(new_n232_), .A4(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT91), .ZN(new_n236_));
  NOR2_X1   g035(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(G169gat), .ZN(new_n238_));
  OR2_X1    g037(.A1(G183gat), .A2(G190gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n213_), .A2(new_n239_), .A3(new_n214_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n235_), .A2(new_n236_), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n236_), .B1(new_n235_), .B2(new_n241_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XOR2_X1   g043(.A(G211gat), .B(G218gat), .Z(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT100), .ZN(new_n246_));
  INV_X1    g045(.A(G204gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT97), .B1(new_n247_), .B2(G197gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT97), .ZN(new_n249_));
  INV_X1    g048(.A(G197gat), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(new_n250_), .A3(G204gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n247_), .A2(G197gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n248_), .A2(new_n251_), .A3(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G211gat), .B(G218gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT100), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n246_), .A2(KEYINPUT21), .A3(new_n253_), .A4(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G197gat), .B(G204gat), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT21), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n254_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n248_), .A2(new_n251_), .A3(new_n260_), .A4(new_n252_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT98), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n263_), .A2(new_n264_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n262_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT99), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n251_), .A2(new_n252_), .ZN(new_n269_));
  NAND4_X1  g068(.A1(new_n269_), .A2(KEYINPUT98), .A3(new_n260_), .A4(new_n248_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n263_), .A2(new_n264_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT99), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n262_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n258_), .B1(new_n268_), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n205_), .B1(new_n244_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n206_), .A2(KEYINPUT101), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT101), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT24), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n280_), .A2(new_n222_), .A3(new_n207_), .A4(new_n233_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n277_), .B(new_n279_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n228_), .A2(new_n231_), .A3(new_n226_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n216_), .A4(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT102), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n240_), .A2(new_n285_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n213_), .A2(new_n239_), .A3(KEYINPUT102), .A4(new_n214_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n238_), .A3(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n284_), .A2(new_n257_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n273_), .B1(new_n272_), .B2(new_n262_), .ZN(new_n291_));
  AOI211_X1 g090(.A(KEYINPUT99), .B(new_n261_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n290_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT103), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n268_), .A2(new_n274_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(KEYINPUT103), .A3(new_n290_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT104), .B1(new_n276_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n205_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n235_), .A2(new_n241_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT91), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n235_), .A2(new_n236_), .A3(new_n241_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n257_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n300_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT104), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(new_n295_), .A4(new_n297_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n299_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n203_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n284_), .A2(new_n288_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n204_), .B1(new_n305_), .B2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n275_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n310_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G8gat), .B(G36gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(KEYINPUT18), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G64gat), .B(G92gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n317_), .B(new_n318_), .Z(new_n319_));
  NAND3_X1  g118(.A1(new_n309_), .A2(new_n315_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT27), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n244_), .A2(new_n275_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n293_), .A2(KEYINPUT20), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n203_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n312_), .A2(new_n313_), .A3(new_n310_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n319_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n321_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n320_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G22gat), .B(G50gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333_));
  INV_X1    g132(.A(G141gat), .ZN(new_n334_));
  INV_X1    g133(.A(G148gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT95), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n336_), .B(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340_));
  XOR2_X1   g139(.A(new_n340_), .B(KEYINPUT2), .Z(new_n341_));
  OAI211_X1 g140(.A(new_n332_), .B(new_n333_), .C1(new_n339_), .C2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n333_), .A2(KEYINPUT1), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n332_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n333_), .A2(KEYINPUT1), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n336_), .B(new_n340_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n347_), .A2(KEYINPUT29), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(KEYINPUT29), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G228gat), .A2(G233gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n352_), .B(new_n353_), .Z(new_n354_));
  NAND3_X1  g153(.A1(new_n305_), .A2(new_n351_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT96), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n305_), .A2(new_n351_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n354_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n350_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n361_));
  AND4_X1   g160(.A1(new_n356_), .A2(new_n360_), .A3(new_n350_), .A4(new_n355_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n331_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(new_n356_), .A3(new_n355_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n350_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n357_), .A2(new_n350_), .A3(new_n360_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n330_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n363_), .A2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G127gat), .B(G134gat), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n370_), .A2(KEYINPUT93), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(KEYINPUT93), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G113gat), .B(G120gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(new_n347_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n376_), .A2(new_n342_), .A3(new_n377_), .A4(new_n346_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G225gat), .A2(G233gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n379_), .A2(KEYINPUT4), .A3(new_n380_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT4), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n378_), .A2(new_n347_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n382_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G85gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT0), .B(G57gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  OR3_X1    g191(.A1(new_n384_), .A2(new_n388_), .A3(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n392_), .B1(new_n384_), .B2(new_n388_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n329_), .A2(new_n369_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT107), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n276_), .A2(new_n298_), .A3(KEYINPUT104), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT103), .B1(new_n296_), .B2(new_n290_), .ZN(new_n401_));
  AOI211_X1 g200(.A(new_n294_), .B(new_n289_), .C1(new_n268_), .C2(new_n274_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n307_), .B1(new_n403_), .B2(new_n306_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n315_), .B1(new_n400_), .B2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n327_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n320_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n399_), .B1(new_n407_), .B2(new_n321_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n319_), .B1(new_n309_), .B2(new_n315_), .ZN(new_n409_));
  AOI211_X1 g208(.A(new_n314_), .B(new_n327_), .C1(new_n299_), .C2(new_n308_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n399_), .B(new_n321_), .C1(new_n409_), .C2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n398_), .B1(new_n408_), .B2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n392_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n385_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n416_), .B1(new_n394_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n394_), .A2(new_n417_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT105), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT105), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n394_), .A2(new_n421_), .A3(new_n417_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n418_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(new_n320_), .A3(new_n406_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n319_), .A2(KEYINPUT32), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n309_), .A2(new_n315_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT106), .ZN(new_n427_));
  INV_X1    g226(.A(new_n425_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n427_), .B1(new_n326_), .B2(new_n428_), .ZN(new_n429_));
  AOI211_X1 g228(.A(KEYINPUT106), .B(new_n425_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n395_), .B(new_n426_), .C1(new_n429_), .C2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n424_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n369_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n413_), .A2(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G71gat), .B(G99gat), .Z(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT92), .B(G43gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n438_), .B(KEYINPUT30), .Z(new_n439_));
  XNOR2_X1  g238(.A(new_n304_), .B(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(G15gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT94), .B1(new_n440_), .B2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n244_), .B(new_n439_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n443_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT31), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT31), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n444_), .A2(new_n450_), .A3(new_n447_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n378_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n449_), .A2(new_n377_), .A3(new_n451_), .A4(new_n376_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n329_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n321_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT107), .ZN(new_n459_));
  AOI211_X1 g258(.A(new_n369_), .B(new_n457_), .C1(new_n459_), .C2(new_n411_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n395_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n435_), .A2(new_n456_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT78), .B(G1gat), .ZN(new_n463_));
  INV_X1    g262(.A(G8gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT14), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G15gat), .B(G22gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT79), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G8gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n467_), .B(KEYINPUT79), .ZN(new_n472_));
  INV_X1    g271(.A(new_n470_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G29gat), .B(G36gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G43gat), .B(G50gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT15), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT84), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n471_), .A2(new_n474_), .A3(new_n478_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G229gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT85), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n481_), .A2(new_n482_), .A3(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n475_), .B(new_n478_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n487_), .A2(new_n483_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G113gat), .B(G141gat), .Z(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT87), .ZN(new_n491_));
  XOR2_X1   g290(.A(G169gat), .B(G197gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT86), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n489_), .B(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n462_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(G85gat), .ZN(new_n499_));
  INV_X1    g298(.A(G92gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G85gat), .A2(G92gat), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT9), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n501_), .A2(new_n502_), .B1(new_n503_), .B2(G92gat), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT66), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n501_), .A2(new_n503_), .A3(new_n502_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n507_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT66), .B1(new_n509_), .B2(new_n504_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT6), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(KEYINPUT10), .B(G99gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT64), .B(G106gat), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT65), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n515_), .A2(KEYINPUT65), .A3(new_n516_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n514_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n511_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT8), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT6), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT68), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT68), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT6), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n512_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT69), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n526_), .A3(new_n512_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n524_), .A2(new_n526_), .A3(new_n512_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT69), .B1(new_n532_), .B2(new_n527_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(G99gat), .A2(G106gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT7), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n531_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n501_), .A2(new_n502_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n522_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n522_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n535_), .A2(new_n513_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT67), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n535_), .A2(KEYINPUT67), .A3(new_n513_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n540_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n521_), .B1(new_n539_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G57gat), .B(G64gat), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n547_), .A2(KEYINPUT11), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(KEYINPUT11), .ZN(new_n549_));
  XOR2_X1   g348(.A(G71gat), .B(G78gat), .Z(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n549_), .A2(new_n550_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n546_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT12), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT72), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n555_), .A2(KEYINPUT72), .A3(new_n556_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT73), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n511_), .A2(new_n520_), .A3(KEYINPUT71), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT71), .ZN(new_n564_));
  INV_X1    g363(.A(new_n519_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n513_), .B1(new_n565_), .B2(new_n517_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n508_), .A2(new_n510_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n564_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n563_), .B(new_n568_), .C1(new_n539_), .C2(new_n545_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n569_), .A2(KEYINPUT12), .A3(new_n554_), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n553_), .B(new_n521_), .C1(new_n539_), .C2(new_n545_), .ZN(new_n571_));
  INV_X1    g370(.A(G230gat), .ZN(new_n572_));
  INV_X1    g371(.A(G233gat), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n571_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n561_), .A2(new_n562_), .A3(new_n570_), .A4(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT72), .B1(new_n555_), .B2(new_n556_), .ZN(new_n577_));
  AOI211_X1 g376(.A(new_n558_), .B(KEYINPUT12), .C1(new_n546_), .C2(new_n554_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n575_), .B(new_n570_), .C1(new_n577_), .C2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT73), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n571_), .B(KEYINPUT70), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(new_n555_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n572_), .A2(new_n573_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n576_), .A2(new_n580_), .A3(new_n584_), .ZN(new_n585_));
  XOR2_X1   g384(.A(G120gat), .B(G148gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G176gat), .B(G204gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n585_), .A2(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n576_), .A2(new_n580_), .A3(new_n584_), .A4(new_n590_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n594_), .A2(KEYINPUT13), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(KEYINPUT13), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT81), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n475_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(G231gat), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n600_), .A2(new_n573_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n471_), .A2(new_n474_), .A3(KEYINPUT81), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n599_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n602_), .B1(new_n599_), .B2(new_n603_), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n553_), .B(KEYINPUT80), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OR3_X1    g406(.A1(new_n604_), .A2(new_n605_), .A3(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n607_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n609_));
  XOR2_X1   g408(.A(G127gat), .B(G155gat), .Z(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT82), .B(KEYINPUT16), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n608_), .A2(new_n609_), .A3(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n608_), .A2(new_n609_), .A3(KEYINPUT83), .ZN(new_n617_));
  AOI22_X1  g416(.A1(KEYINPUT17), .A2(new_n616_), .B1(new_n617_), .B2(new_n614_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n617_), .A2(KEYINPUT17), .A3(new_n614_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n478_), .B(new_n521_), .C1(new_n539_), .C2(new_n545_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G232gat), .A2(G233gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT34), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT35), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n621_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n569_), .A2(KEYINPUT75), .A3(new_n479_), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT75), .B1(new_n569_), .B2(new_n479_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n628_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n624_), .A2(new_n625_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT76), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n632_), .B1(new_n627_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n631_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n569_), .A2(new_n479_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT75), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n569_), .A2(KEYINPUT75), .A3(new_n479_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(new_n628_), .A3(new_n634_), .ZN(new_n642_));
  XOR2_X1   g441(.A(G190gat), .B(G218gat), .Z(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT77), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G134gat), .B(G162gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(KEYINPUT36), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n636_), .A2(new_n642_), .A3(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n646_), .B(KEYINPUT36), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n649_), .B1(new_n636_), .B2(new_n642_), .ZN(new_n650_));
  OAI21_X1  g449(.A(KEYINPUT37), .B1(new_n648_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n649_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n631_), .A2(new_n635_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n634_), .B1(new_n641_), .B2(new_n628_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n652_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT37), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n636_), .A2(new_n642_), .A3(new_n647_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n651_), .A2(new_n658_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n597_), .A2(new_n620_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n498_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n395_), .A3(new_n463_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT38), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n397_), .B1(new_n459_), .B2(new_n411_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n369_), .B1(new_n424_), .B2(new_n431_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n456_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n457_), .B1(new_n459_), .B2(new_n411_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n433_), .A3(new_n461_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n655_), .A2(new_n657_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n620_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n597_), .A2(new_n497_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n673_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G1gat), .B1(new_n676_), .B2(new_n396_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n663_), .A2(new_n664_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n665_), .A2(new_n677_), .A3(new_n678_), .ZN(G1324gat));
  INV_X1    g478(.A(new_n669_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n662_), .A2(new_n464_), .A3(new_n680_), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n676_), .A2(new_n669_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT39), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(new_n683_), .A3(G8gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n682_), .B2(G8gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1325gat));
  OAI21_X1  g487(.A(G15gat), .B1(new_n676_), .B2(new_n456_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT108), .B(KEYINPUT41), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n690_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n662_), .A2(new_n442_), .A3(new_n455_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n691_), .A2(new_n692_), .A3(new_n693_), .ZN(G1326gat));
  OAI21_X1  g493(.A(G22gat), .B1(new_n676_), .B2(new_n433_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT42), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n433_), .A2(G22gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n661_), .B2(new_n697_), .ZN(G1327gat));
  INV_X1    g497(.A(new_n597_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n674_), .A2(new_n672_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n498_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n701_), .A2(G29gat), .A3(new_n396_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n659_), .ZN(new_n703_));
  AOI211_X1 g502(.A(KEYINPUT43), .B(new_n703_), .C1(new_n668_), .C2(new_n670_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n651_), .A2(new_n658_), .A3(KEYINPUT109), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT109), .B1(new_n651_), .B2(new_n658_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n671_), .A2(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n706_), .B1(new_n711_), .B2(KEYINPUT43), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n709_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT43), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n713_), .A2(KEYINPUT110), .A3(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n705_), .B1(new_n712_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n675_), .A2(new_n620_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n716_), .A2(KEYINPUT44), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT44), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n706_), .B(KEYINPUT43), .C1(new_n462_), .C2(new_n709_), .ZN(new_n721_));
  OAI21_X1  g520(.A(KEYINPUT110), .B1(new_n713_), .B2(new_n714_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n704_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n720_), .B1(new_n723_), .B2(new_n717_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(new_n724_), .A3(new_n395_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n725_), .A2(KEYINPUT111), .A3(G29gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(KEYINPUT111), .B1(new_n725_), .B2(G29gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n702_), .B1(new_n726_), .B2(new_n727_), .ZN(G1328gat));
  NAND3_X1  g527(.A1(new_n719_), .A2(new_n724_), .A3(new_n680_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(G36gat), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n701_), .A2(G36gat), .A3(new_n669_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT45), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT46), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n730_), .A2(new_n733_), .A3(KEYINPUT46), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(G1329gat));
  NAND4_X1  g537(.A1(new_n719_), .A2(new_n724_), .A3(G43gat), .A4(new_n455_), .ZN(new_n739_));
  INV_X1    g538(.A(G43gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n740_), .B1(new_n701_), .B2(new_n456_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(G1330gat));
  NAND4_X1  g543(.A1(new_n719_), .A2(new_n724_), .A3(G50gat), .A4(new_n369_), .ZN(new_n745_));
  INV_X1    g544(.A(G50gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n701_), .B2(new_n433_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1331gat));
  NAND2_X1  g547(.A1(new_n597_), .A2(new_n497_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(new_n620_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n673_), .A2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G57gat), .B1(new_n751_), .B2(new_n396_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n462_), .A2(new_n749_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n620_), .A2(new_n659_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n396_), .A2(G57gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(G1332gat));
  OAI21_X1  g556(.A(G64gat), .B1(new_n751_), .B2(new_n669_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT48), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n669_), .A2(G64gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n759_), .B1(new_n755_), .B2(new_n760_), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n751_), .B2(new_n456_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT49), .ZN(new_n763_));
  OR2_X1    g562(.A1(new_n456_), .A2(G71gat), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n755_), .B2(new_n764_), .ZN(G1334gat));
  OAI21_X1  g564(.A(G78gat), .B1(new_n751_), .B2(new_n433_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT50), .ZN(new_n767_));
  OR3_X1    g566(.A1(new_n755_), .A2(G78gat), .A3(new_n433_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n769_), .B(new_n770_), .ZN(G1335gat));
  NAND3_X1  g570(.A1(new_n597_), .A2(new_n497_), .A3(new_n620_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n716_), .A2(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G85gat), .B1(new_n774_), .B2(new_n396_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n753_), .A2(KEYINPUT114), .A3(new_n700_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT114), .B1(new_n753_), .B2(new_n700_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n395_), .A2(new_n499_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1336gat));
  INV_X1    g579(.A(new_n778_), .ZN(new_n781_));
  AOI21_X1  g580(.A(G92gat), .B1(new_n781_), .B2(new_n680_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n680_), .A2(G92gat), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT115), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n774_), .A2(new_n785_), .ZN(new_n786_));
  OR3_X1    g585(.A1(new_n782_), .A2(new_n783_), .A3(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n782_), .B2(new_n786_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1337gat));
  NAND3_X1  g588(.A1(new_n781_), .A2(new_n455_), .A3(new_n515_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G99gat), .B1(new_n774_), .B2(new_n456_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g592(.A1(new_n781_), .A2(new_n369_), .A3(new_n516_), .ZN(new_n794_));
  INV_X1    g593(.A(G106gat), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n721_), .A2(new_n722_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n772_), .B1(new_n796_), .B2(new_n705_), .ZN(new_n797_));
  AOI211_X1 g596(.A(KEYINPUT52), .B(new_n795_), .C1(new_n797_), .C2(new_n369_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n716_), .A2(new_n369_), .A3(new_n773_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(G106gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n794_), .B1(new_n798_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT53), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n804_), .B(new_n794_), .C1(new_n798_), .C2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1339gat));
  NAND3_X1  g605(.A1(new_n699_), .A2(new_n754_), .A3(new_n497_), .ZN(new_n807_));
  XOR2_X1   g606(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n660_), .A2(new_n497_), .A3(new_n808_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n576_), .A2(new_n580_), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n579_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n581_), .B(new_n570_), .C1(new_n577_), .C2(new_n578_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n815_), .A2(KEYINPUT55), .B1(new_n583_), .B2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n590_), .B1(new_n814_), .B2(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n818_), .A2(KEYINPUT56), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n591_), .A2(KEYINPUT56), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n814_), .B2(new_n817_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n496_), .B(new_n593_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n481_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n487_), .A2(new_n485_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n494_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n594_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT118), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT118), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n594_), .A2(new_n829_), .A3(new_n826_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n822_), .A2(new_n828_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n672_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n826_), .A2(new_n593_), .ZN(new_n835_));
  OAI22_X1  g634(.A1(KEYINPUT120), .A2(new_n821_), .B1(new_n818_), .B2(KEYINPUT56), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n821_), .A2(KEYINPUT120), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n835_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT58), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT58), .B(new_n835_), .C1(new_n836_), .C2(new_n837_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n659_), .A3(new_n841_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n831_), .B(new_n672_), .C1(KEYINPUT119), .C2(KEYINPUT57), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n834_), .A2(new_n842_), .A3(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n812_), .B1(new_n844_), .B2(new_n620_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n460_), .A2(new_n395_), .A3(new_n455_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n847_), .A2(KEYINPUT121), .ZN(new_n848_));
  OR3_X1    g647(.A1(new_n845_), .A2(new_n846_), .A3(new_n848_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n847_), .A2(KEYINPUT121), .ZN(new_n850_));
  OAI22_X1  g649(.A1(new_n845_), .A2(new_n846_), .B1(new_n850_), .B2(new_n848_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n849_), .A2(new_n496_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G113gat), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n845_), .A2(new_n846_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  OR3_X1    g654(.A1(new_n855_), .A2(G113gat), .A3(new_n497_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n853_), .A2(new_n856_), .ZN(G1340gat));
  INV_X1    g656(.A(G120gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n699_), .B2(KEYINPUT60), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n854_), .B(new_n859_), .C1(KEYINPUT60), .C2(new_n858_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n849_), .A2(new_n597_), .A3(new_n851_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n858_), .ZN(G1341gat));
  AOI21_X1  g661(.A(G127gat), .B1(new_n854_), .B2(new_n674_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n849_), .A2(new_n851_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n620_), .A2(KEYINPUT122), .ZN(new_n865_));
  MUX2_X1   g664(.A(KEYINPUT122), .B(new_n865_), .S(G127gat), .Z(new_n866_));
  AOI21_X1  g665(.A(new_n863_), .B1(new_n864_), .B2(new_n866_), .ZN(G1342gat));
  NAND3_X1  g666(.A1(new_n849_), .A2(new_n659_), .A3(new_n851_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(G134gat), .ZN(new_n869_));
  OR3_X1    g668(.A1(new_n855_), .A2(G134gat), .A3(new_n672_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1343gat));
  NOR2_X1   g670(.A1(new_n845_), .A2(new_n455_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n680_), .A2(new_n396_), .A3(new_n433_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(new_n334_), .A3(new_n496_), .ZN(new_n876_));
  OAI21_X1  g675(.A(G141gat), .B1(new_n874_), .B2(new_n497_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1344gat));
  NAND3_X1  g677(.A1(new_n875_), .A2(new_n335_), .A3(new_n597_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G148gat), .B1(new_n874_), .B2(new_n699_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(G1345gat));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  OR3_X1    g681(.A1(new_n874_), .A2(new_n620_), .A3(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n874_), .B2(new_n620_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1346gat));
  INV_X1    g684(.A(G162gat), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n874_), .A2(new_n886_), .A3(new_n709_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n874_), .A2(new_n672_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n886_), .B2(new_n888_), .ZN(G1347gat));
  INV_X1    g688(.A(KEYINPUT62), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n680_), .A2(new_n433_), .A3(new_n461_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n845_), .A2(new_n497_), .A3(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT22), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n890_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(G169gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n220_), .B1(new_n892_), .B2(new_n890_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n894_), .B2(new_n896_), .ZN(G1348gat));
  NOR2_X1   g696(.A1(new_n845_), .A2(new_n891_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n597_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G176gat), .ZN(G1349gat));
  INV_X1    g699(.A(new_n898_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n620_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n231_), .A2(new_n226_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(KEYINPUT123), .B2(new_n230_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(KEYINPUT123), .A2(G183gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n902_), .B2(new_n906_), .ZN(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n901_), .B2(new_n703_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n655_), .A2(new_n228_), .A3(new_n657_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n901_), .B2(new_n909_), .ZN(G1351gat));
  NOR3_X1   g709(.A1(new_n669_), .A2(new_n395_), .A3(new_n433_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n872_), .A2(new_n911_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n250_), .B1(new_n912_), .B2(new_n497_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n872_), .A2(G197gat), .A3(new_n496_), .A4(new_n911_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(KEYINPUT124), .ZN(new_n915_));
  INV_X1    g714(.A(new_n911_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n845_), .A2(new_n455_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n917_), .A2(new_n918_), .A3(G197gat), .A4(new_n496_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n913_), .A2(new_n915_), .A3(new_n919_), .ZN(G1352gat));
  NOR2_X1   g719(.A1(new_n247_), .A2(KEYINPUT125), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n247_), .A2(KEYINPUT125), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n917_), .B(new_n597_), .C1(new_n921_), .C2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n912_), .A2(new_n699_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n924_), .B2(new_n922_), .ZN(G1353gat));
  NAND2_X1  g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n917_), .A2(new_n674_), .A3(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(KEYINPUT126), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n927_), .B(new_n929_), .ZN(G1354gat));
  INV_X1    g729(.A(new_n845_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n672_), .A2(G218gat), .ZN(new_n932_));
  NAND4_X1  g731(.A1(new_n931_), .A2(new_n456_), .A3(new_n911_), .A4(new_n932_), .ZN(new_n933_));
  NOR4_X1   g732(.A1(new_n845_), .A2(new_n455_), .A3(new_n703_), .A4(new_n916_), .ZN(new_n934_));
  INV_X1    g733(.A(G218gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n933_), .B1(new_n934_), .B2(new_n935_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT127), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n936_), .A2(new_n937_), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n933_), .B(KEYINPUT127), .C1(new_n934_), .C2(new_n935_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1355gat));
endmodule


