//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n897_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n203_), .B(KEYINPUT90), .Z(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n204_), .B1(G176gat), .B2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT85), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(KEYINPUT85), .A3(KEYINPUT23), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G183gat), .A3(G190gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n211_), .A2(new_n212_), .A3(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(G183gat), .B2(G190gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT91), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n216_), .A2(new_n217_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n207_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G211gat), .B(G218gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT87), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G197gat), .B(G204gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n222_), .A2(KEYINPUT21), .A3(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(new_n223_), .B(KEYINPUT21), .Z(new_n226_));
  OAI21_X1  g025(.A(new_n225_), .B1(new_n222_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n203_), .A2(KEYINPUT24), .ZN(new_n228_));
  INV_X1    g027(.A(G169gat), .ZN(new_n229_));
  INV_X1    g028(.A(G176gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  MUX2_X1   g030(.A(KEYINPUT24), .B(new_n228_), .S(new_n231_), .Z(new_n232_));
  NAND2_X1  g031(.A1(new_n209_), .A2(new_n214_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT25), .B(G183gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT26), .B(G190gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  AND3_X1   g035(.A1(new_n232_), .A2(new_n233_), .A3(new_n236_), .ZN(new_n237_));
  NOR3_X1   g036(.A1(new_n220_), .A2(new_n227_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT20), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G226gat), .A2(G233gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT84), .ZN(new_n245_));
  INV_X1    g044(.A(G190gat), .ZN(new_n246_));
  OR3_X1    g045(.A1(new_n245_), .A2(new_n246_), .A3(KEYINPUT26), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT26), .B1(new_n245_), .B2(new_n246_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n247_), .A2(new_n234_), .A3(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n232_), .A2(new_n215_), .A3(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n233_), .B1(G183gat), .B2(G190gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n205_), .A2(KEYINPUT86), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n229_), .A2(KEYINPUT22), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT86), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n230_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n251_), .B(new_n203_), .C1(new_n252_), .C2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n250_), .A2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n227_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n240_), .A2(new_n244_), .A3(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n227_), .B1(new_n220_), .B2(new_n237_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n260_), .B(KEYINPUT20), .C1(new_n227_), .C2(new_n257_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT92), .ZN(new_n262_));
  AND3_X1   g061(.A1(new_n261_), .A2(new_n262_), .A3(new_n243_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n262_), .B1(new_n261_), .B2(new_n243_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n259_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G8gat), .B(G36gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT18), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G64gat), .B(G92gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(new_n268_), .Z(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n265_), .A2(new_n270_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n259_), .B(new_n269_), .C1(new_n263_), .C2(new_n264_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G155gat), .A2(G162gat), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G141gat), .A2(G148gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n278_), .B(KEYINPUT3), .Z(new_n279_));
  NAND2_X1  g078(.A1(G141gat), .A2(G148gat), .ZN(new_n280_));
  XOR2_X1   g079(.A(new_n280_), .B(KEYINPUT2), .Z(new_n281_));
  OAI211_X1 g080(.A(new_n275_), .B(new_n277_), .C1(new_n279_), .C2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n276_), .B1(KEYINPUT1), .B2(new_n275_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(KEYINPUT1), .B2(new_n275_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n278_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(new_n280_), .A3(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n282_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G127gat), .B(G134gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G113gat), .B(G120gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n282_), .A2(new_n286_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n290_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n291_), .A2(KEYINPUT4), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G225gat), .A2(G233gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT93), .B(KEYINPUT4), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n296_), .A2(KEYINPUT94), .A3(new_n298_), .A4(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT94), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n298_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n302_), .B1(new_n303_), .B2(new_n295_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n301_), .A2(new_n304_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n291_), .A2(new_n294_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n297_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G1gat), .B(G29gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT0), .ZN(new_n309_));
  INV_X1    g108(.A(G57gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(G85gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n305_), .A2(new_n307_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT95), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT33), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n301_), .A2(new_n304_), .B1(new_n306_), .B2(new_n297_), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT95), .B1(new_n317_), .B2(new_n312_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT33), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n296_), .A2(new_n297_), .A3(new_n300_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n312_), .B1(new_n306_), .B2(new_n298_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n318_), .A2(new_n319_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n274_), .A2(new_n316_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT97), .ZN(new_n324_));
  OR3_X1    g123(.A1(new_n317_), .A2(new_n324_), .A3(new_n312_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n324_), .B1(new_n317_), .B2(new_n312_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(new_n326_), .A3(new_n313_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n261_), .A2(new_n243_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n240_), .A2(KEYINPUT96), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT96), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n329_), .A2(new_n258_), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n328_), .B1(new_n332_), .B2(new_n243_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n269_), .A2(KEYINPUT32), .ZN(new_n334_));
  MUX2_X1   g133(.A(new_n333_), .B(new_n265_), .S(new_n334_), .Z(new_n335_));
  NAND2_X1  g134(.A1(new_n327_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n323_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n257_), .B(KEYINPUT30), .ZN(new_n338_));
  XOR2_X1   g137(.A(G71gat), .B(G99gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(G43gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G227gat), .A2(G233gat), .ZN(new_n341_));
  INV_X1    g140(.A(G15gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n340_), .B(new_n343_), .Z(new_n344_));
  XNOR2_X1  g143(.A(new_n338_), .B(new_n344_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n345_), .A2(KEYINPUT31), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(KEYINPUT31), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n346_), .A2(new_n290_), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n290_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT29), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n287_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G22gat), .B(G50gat), .Z(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n352_), .B(KEYINPUT28), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n355_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n292_), .A2(KEYINPUT29), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(new_n227_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G78gat), .B(G106gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n362_), .B1(G228gat), .B2(G233gat), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n363_), .B1(new_n361_), .B2(new_n227_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n365_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n367_), .A2(KEYINPUT88), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n360_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n357_), .A2(new_n359_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n367_), .B(new_n370_), .C1(new_n374_), .C2(KEYINPUT88), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n350_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT27), .ZN(new_n379_));
  OR2_X1    g178(.A1(new_n333_), .A2(new_n269_), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n272_), .A2(KEYINPUT27), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n379_), .A2(new_n273_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n375_), .B(new_n373_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n346_), .A2(new_n347_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n293_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n346_), .A2(new_n347_), .A3(new_n290_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n376_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n327_), .B1(new_n383_), .B2(new_n387_), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n337_), .A2(new_n378_), .B1(new_n382_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G229gat), .A2(G233gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G36gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G29gat), .ZN(new_n393_));
  INV_X1    g192(.A(G29gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(G36gat), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n393_), .A2(new_n395_), .A3(KEYINPUT73), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT73), .B1(new_n393_), .B2(new_n395_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G43gat), .B(G50gat), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G43gat), .B(G50gat), .Z(new_n400_));
  INV_X1    g199(.A(KEYINPUT73), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n394_), .A2(G36gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n392_), .A2(G29gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n401_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n393_), .A2(new_n395_), .A3(KEYINPUT73), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n400_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT15), .B1(new_n399_), .B2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n398_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n404_), .A2(new_n405_), .A3(new_n400_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT15), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n408_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n407_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT80), .B(G8gat), .ZN(new_n413_));
  INV_X1    g212(.A(G1gat), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT14), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G15gat), .B(G22gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(G1gat), .B(G8gat), .Z(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n418_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n412_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n408_), .A2(new_n409_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n391_), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n421_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n427_), .A2(new_n409_), .A3(new_n408_), .A4(new_n419_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n425_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n429_), .A2(new_n390_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G113gat), .B(G141gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G169gat), .B(G197gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n434_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n436_), .B1(new_n426_), .B2(new_n430_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT83), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n202_), .B1(new_n389_), .B2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n313_), .A2(new_n314_), .A3(new_n319_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n320_), .A2(new_n321_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n318_), .A2(new_n319_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n445_), .A2(new_n274_), .B1(new_n335_), .B2(new_n327_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n378_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n383_), .A2(new_n387_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n327_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n380_), .A2(new_n381_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(new_n274_), .B2(KEYINPUT27), .ZN(new_n452_));
  OAI22_X1  g251(.A1(new_n446_), .A2(new_n447_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n439_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(KEYINPUT98), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n440_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT67), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G99gat), .A2(G106gat), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT6), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  AND2_X1   g262(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(G106gat), .ZN(new_n467_));
  AOI21_X1  g266(.A(KEYINPUT65), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT65), .ZN(new_n469_));
  NOR4_X1   g268(.A1(new_n464_), .A2(new_n465_), .A3(new_n469_), .A4(G106gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n463_), .B1(new_n468_), .B2(new_n470_), .ZN(new_n471_));
  OR2_X1    g270(.A1(G85gat), .A2(G92gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  OR2_X1    g273(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(G85gat), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT9), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n474_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n457_), .B1(new_n471_), .B2(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(new_n467_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n469_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n482_), .A2(KEYINPUT65), .A3(new_n467_), .A4(new_n483_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n472_), .A2(new_n473_), .ZN(new_n488_));
  INV_X1    g287(.A(G85gat), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n489_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n490_), .B2(KEYINPUT9), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n487_), .A2(new_n491_), .A3(KEYINPUT67), .A4(new_n463_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT7), .ZN(new_n493_));
  INV_X1    g292(.A(G99gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(new_n467_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n495_), .A2(new_n460_), .A3(new_n461_), .A4(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G85gat), .B(G92gat), .Z(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(KEYINPUT8), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT8), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n497_), .A2(new_n501_), .A3(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n481_), .A2(new_n492_), .A3(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT35), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G232gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT34), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n504_), .A2(new_n412_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n481_), .A2(new_n492_), .A3(new_n503_), .A4(new_n424_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT74), .B1(new_n504_), .B2(new_n412_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n507_), .A2(KEYINPUT35), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n509_), .B(new_n510_), .C1(new_n511_), .C2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n503_), .A2(new_n492_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n462_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n515_));
  AOI21_X1  g314(.A(KEYINPUT67), .B1(new_n515_), .B2(new_n491_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n412_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT74), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n512_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n508_), .A2(new_n505_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(new_n510_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT79), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n513_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n513_), .B2(new_n522_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G190gat), .B(G218gat), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n526_), .A2(KEYINPUT75), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(KEYINPUT75), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G134gat), .B(G162gat), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n529_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT36), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n532_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT36), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n530_), .ZN(new_n536_));
  AND3_X1   g335(.A1(new_n533_), .A2(new_n536_), .A3(KEYINPUT77), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT77), .B1(new_n533_), .B2(new_n536_), .ZN(new_n538_));
  OAI22_X1  g337(.A1(new_n524_), .A2(new_n525_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n536_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n513_), .A2(new_n522_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT76), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n513_), .A2(new_n522_), .A3(KEYINPUT76), .A4(new_n540_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n539_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT37), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n537_), .A2(new_n538_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT78), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n513_), .A2(new_n522_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n547_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n546_), .A2(new_n547_), .B1(new_n545_), .B2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(G64gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(G57gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n310_), .A2(G64gat), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT68), .ZN(new_n556_));
  AND3_X1   g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT11), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n310_), .A2(G64gat), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n553_), .A2(G57gat), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT68), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT11), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  AND2_X1   g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566_));
  NOR2_X1   g365(.A1(G71gat), .A2(G78gat), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n559_), .A2(new_n565_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n562_), .A2(new_n564_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n568_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(KEYINPUT11), .A3(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(new_n422_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT81), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G127gat), .B(G155gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT16), .ZN(new_n579_));
  XOR2_X1   g378(.A(G183gat), .B(G211gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT17), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  OR3_X1    g382(.A1(new_n576_), .A2(new_n577_), .A3(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n583_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n576_), .A2(new_n582_), .A3(new_n581_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n552_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(G230gat), .A2(G233gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT64), .Z(new_n590_));
  NOR2_X1   g389(.A1(new_n514_), .A2(new_n516_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n590_), .B1(new_n591_), .B2(new_n573_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n593_));
  AOI211_X1 g392(.A(new_n563_), .B(new_n568_), .C1(new_n562_), .C2(new_n564_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n571_), .B1(new_n570_), .B2(KEYINPUT11), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n594_), .B1(new_n595_), .B2(new_n565_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n593_), .B(new_n596_), .C1(new_n514_), .C2(new_n516_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n504_), .B2(new_n596_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n592_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT70), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n596_), .B1(new_n514_), .B2(new_n516_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n573_), .A2(new_n481_), .A3(new_n492_), .A4(new_n503_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n590_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n592_), .B(KEYINPUT70), .C1(new_n598_), .C2(new_n600_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n603_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(G176gat), .B(G204gat), .Z(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(G120gat), .B(G148gat), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT72), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n612_), .B(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n609_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n615_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n603_), .A2(new_n607_), .A3(new_n608_), .A4(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT13), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n588_), .A2(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT82), .Z(new_n622_));
  NAND2_X1  g421(.A1(new_n456_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(new_n414_), .A3(new_n327_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT38), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n546_), .B(KEYINPUT99), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n620_), .A2(new_n438_), .A3(new_n587_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n453_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G1gat), .B1(new_n630_), .B2(new_n449_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n626_), .A2(new_n631_), .ZN(G1324gat));
  NAND2_X1  g431(.A1(new_n452_), .A2(new_n413_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n453_), .A2(new_n627_), .A3(new_n452_), .A4(new_n629_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n634_), .A2(new_n635_), .A3(G8gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n634_), .B2(G8gat), .ZN(new_n637_));
  OAI22_X1  g436(.A1(new_n623_), .A2(new_n633_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT101), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT101), .ZN(new_n640_));
  OAI221_X1 g439(.A(new_n640_), .B1(new_n636_), .B2(new_n637_), .C1(new_n623_), .C2(new_n633_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n639_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n639_), .B2(new_n641_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(G1325gat));
  INV_X1    g444(.A(new_n350_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G15gat), .B1(new_n630_), .B2(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT41), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n624_), .A2(new_n342_), .A3(new_n350_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1326gat));
  OAI21_X1  g449(.A(G22gat), .B1(new_n630_), .B2(new_n376_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n651_), .A2(KEYINPUT42), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(KEYINPUT42), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n376_), .A2(G22gat), .ZN(new_n654_));
  OAI22_X1  g453(.A1(new_n652_), .A2(new_n653_), .B1(new_n623_), .B2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT102), .ZN(G1327gat));
  OAI21_X1  g455(.A(KEYINPUT43), .B1(new_n389_), .B2(new_n552_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  INV_X1    g457(.A(new_n552_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n453_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n657_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n587_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n620_), .A2(new_n438_), .A3(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT103), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n661_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n661_), .A2(KEYINPUT44), .A3(new_n665_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n668_), .A2(G29gat), .A3(new_n327_), .A4(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n546_), .A2(new_n587_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n620_), .A2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n672_), .B1(new_n440_), .B2(new_n455_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n394_), .B1(new_n674_), .B2(new_n449_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n670_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT104), .ZN(G1328gat));
  NOR2_X1   g476(.A1(new_n382_), .A2(G36gat), .ZN(new_n678_));
  XOR2_X1   g477(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n673_), .A2(new_n678_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n673_), .B2(new_n678_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT44), .B1(new_n661_), .B2(new_n665_), .ZN(new_n684_));
  AOI211_X1 g483(.A(new_n667_), .B(new_n664_), .C1(new_n657_), .C2(new_n660_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n684_), .A2(new_n685_), .A3(new_n382_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n686_), .B2(new_n392_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT46), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n683_), .B(KEYINPUT46), .C1(new_n686_), .C2(new_n392_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1329gat));
  NAND4_X1  g490(.A1(new_n668_), .A2(G43gat), .A3(new_n350_), .A4(new_n669_), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT106), .B(G43gat), .Z(new_n693_));
  OAI21_X1  g492(.A(new_n693_), .B1(new_n674_), .B2(new_n646_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n696_));
  XNOR2_X1  g495(.A(new_n695_), .B(new_n696_), .ZN(G1330gat));
  AOI21_X1  g496(.A(G50gat), .B1(new_n673_), .B2(new_n377_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n668_), .A2(G50gat), .A3(new_n377_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n699_), .B2(new_n669_), .ZN(G1331gat));
  NAND2_X1  g499(.A1(new_n453_), .A2(new_n627_), .ZN(new_n701_));
  NOR4_X1   g500(.A1(new_n701_), .A2(new_n620_), .A3(new_n662_), .A4(new_n454_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G57gat), .B1(new_n703_), .B2(new_n449_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n389_), .A2(new_n438_), .A3(new_n620_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n705_), .A2(new_n588_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(new_n310_), .A3(new_n327_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n707_), .ZN(G1332gat));
  AOI21_X1  g507(.A(new_n553_), .B1(new_n702_), .B2(new_n452_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT48), .Z(new_n710_));
  NOR2_X1   g509(.A1(new_n382_), .A2(G64gat), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT108), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n706_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n710_), .A2(new_n713_), .ZN(G1333gat));
  INV_X1    g513(.A(G71gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n702_), .B2(new_n350_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT49), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n706_), .A2(new_n715_), .A3(new_n350_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1334gat));
  INV_X1    g518(.A(G78gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n702_), .B2(new_n377_), .ZN(new_n721_));
  XOR2_X1   g520(.A(new_n721_), .B(KEYINPUT50), .Z(new_n722_));
  NAND3_X1  g521(.A1(new_n706_), .A2(new_n720_), .A3(new_n377_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1335gat));
  NAND2_X1  g523(.A1(new_n705_), .A2(new_n671_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(new_n489_), .A3(new_n327_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n661_), .A2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n657_), .A2(new_n660_), .A3(KEYINPUT109), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n620_), .A2(new_n438_), .A3(new_n587_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n729_), .A2(new_n730_), .A3(new_n731_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n732_), .A2(new_n327_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n727_), .B1(new_n733_), .B2(new_n489_), .ZN(G1336gat));
  AOI21_X1  g533(.A(G92gat), .B1(new_n726_), .B2(new_n452_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n382_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n732_), .B2(new_n736_), .ZN(G1337gat));
  NAND4_X1  g536(.A1(new_n729_), .A2(new_n350_), .A3(new_n730_), .A4(new_n731_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(G99gat), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n350_), .A2(new_n466_), .ZN(new_n740_));
  AOI21_X1  g539(.A(KEYINPUT110), .B1(new_n726_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g542(.A1(new_n705_), .A2(new_n467_), .A3(new_n377_), .A4(new_n671_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT111), .Z(new_n745_));
  NAND2_X1  g544(.A1(new_n731_), .A2(new_n377_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n389_), .A2(KEYINPUT43), .A3(new_n552_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n658_), .B1(new_n453_), .B2(new_n659_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT52), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n751_), .A3(G106gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n750_), .B2(G106gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(KEYINPUT112), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n746_), .B1(new_n657_), .B2(new_n660_), .ZN(new_n755_));
  OAI211_X1 g554(.A(KEYINPUT112), .B(KEYINPUT52), .C1(new_n755_), .C2(new_n467_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n745_), .B1(new_n754_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT53), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n745_), .B(new_n760_), .C1(new_n754_), .C2(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1339gat));
  NAND2_X1  g561(.A1(new_n618_), .A2(new_n438_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n603_), .A2(new_n764_), .A3(new_n608_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n605_), .B1(new_n598_), .B2(new_n600_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n590_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n605_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(new_n599_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n604_), .A2(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n768_), .B1(new_n770_), .B2(new_n597_), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n590_), .A2(new_n766_), .B1(new_n771_), .B2(KEYINPUT55), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n765_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(new_n615_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT56), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n773_), .A2(KEYINPUT56), .A3(new_n615_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n763_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n423_), .A2(new_n391_), .A3(new_n425_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n429_), .A2(new_n390_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(new_n434_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n437_), .A2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT113), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT113), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n437_), .A2(new_n784_), .A3(new_n781_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n619_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n546_), .B1(new_n778_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n786_), .A2(new_n618_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT56), .B1(new_n773_), .B2(new_n615_), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n775_), .B(new_n617_), .C1(new_n765_), .C2(new_n772_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n792_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n552_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n776_), .A2(new_n777_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n798_), .A2(KEYINPUT114), .A3(KEYINPUT58), .A4(new_n792_), .ZN(new_n799_));
  OAI211_X1 g598(.A(KEYINPUT58), .B(new_n792_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n797_), .A2(new_n799_), .A3(new_n802_), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n438_), .B(new_n618_), .C1(new_n793_), .C2(new_n794_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n787_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(KEYINPUT57), .A3(new_n546_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n791_), .A2(new_n803_), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n662_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n620_), .A2(new_n587_), .A3(new_n439_), .A4(new_n552_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n588_), .A2(KEYINPUT54), .A3(new_n620_), .A4(new_n439_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n808_), .A2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n452_), .A2(new_n449_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(new_n387_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n815_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n815_), .A2(KEYINPUT59), .A3(new_n818_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n439_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(G113gat), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n438_), .A2(new_n824_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n819_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT115), .B1(new_n825_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n829_));
  OAI221_X1 g628(.A(new_n829_), .B1(new_n819_), .B2(new_n826_), .C1(new_n823_), .C2(new_n824_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(G1340gat));
  INV_X1    g630(.A(new_n819_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n620_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT60), .ZN(new_n834_));
  XOR2_X1   g633(.A(KEYINPUT116), .B(G120gat), .Z(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n832_), .A2(new_n837_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n821_), .A2(new_n822_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n620_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n838_), .B1(new_n840_), .B2(new_n835_), .ZN(G1341gat));
  OR2_X1    g640(.A1(KEYINPUT117), .A2(G127gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n587_), .A2(KEYINPUT117), .A3(G127gat), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n839_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G127gat), .B1(new_n832_), .B2(new_n587_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(G1342gat));
  OAI21_X1  g645(.A(G134gat), .B1(new_n839_), .B2(new_n552_), .ZN(new_n847_));
  OR2_X1    g646(.A1(new_n627_), .A2(G134gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n819_), .B2(new_n848_), .ZN(G1343gat));
  AOI21_X1  g648(.A(new_n383_), .B1(new_n808_), .B2(new_n814_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n816_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n438_), .ZN(new_n852_));
  OR3_X1    g651(.A1(new_n851_), .A2(KEYINPUT119), .A3(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT119), .B1(new_n851_), .B2(new_n852_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  XOR2_X1   g654(.A(KEYINPUT118), .B(G141gat), .Z(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(G1344gat));
  NOR2_X1   g656(.A1(new_n851_), .A2(new_n620_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT120), .B(G148gat), .Z(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1345gat));
  OR3_X1    g659(.A1(new_n851_), .A2(KEYINPUT121), .A3(new_n662_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT121), .B1(new_n851_), .B2(new_n662_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1346gat));
  OAI21_X1  g664(.A(G162gat), .B1(new_n851_), .B2(new_n552_), .ZN(new_n866_));
  OR2_X1    g665(.A1(new_n627_), .A2(G162gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n866_), .B1(new_n851_), .B2(new_n867_), .ZN(G1347gat));
  NAND2_X1  g667(.A1(new_n452_), .A2(new_n449_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n869_), .A2(new_n646_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n438_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT122), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n813_), .B1(new_n807_), .B2(new_n662_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n377_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n229_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  XOR2_X1   g674(.A(new_n875_), .B(KEYINPUT62), .Z(new_n876_));
  NAND3_X1  g675(.A1(new_n815_), .A2(new_n376_), .A3(new_n870_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT123), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT123), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n874_), .A2(new_n879_), .A3(new_n870_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(new_n205_), .A3(new_n438_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n876_), .A2(new_n882_), .ZN(G1348gat));
  NAND4_X1  g682(.A1(new_n874_), .A2(G176gat), .A3(new_n833_), .A4(new_n870_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n620_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(G176gat), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI211_X1 g687(.A(KEYINPUT124), .B(new_n884_), .C1(new_n885_), .C2(G176gat), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1349gat));
  NOR3_X1   g689(.A1(new_n877_), .A2(KEYINPUT125), .A3(new_n662_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(G183gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(KEYINPUT125), .B1(new_n877_), .B2(new_n662_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n662_), .A2(new_n234_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n892_), .A2(new_n893_), .B1(new_n881_), .B2(new_n894_), .ZN(G1350gat));
  INV_X1    g694(.A(new_n235_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n627_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n881_), .A2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n552_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n246_), .ZN(G1351gat));
  INV_X1    g699(.A(new_n383_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n869_), .ZN(new_n902_));
  AOI21_X1  g701(.A(KEYINPUT57), .B1(new_n805_), .B2(new_n546_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n546_), .ZN(new_n904_));
  AOI211_X1 g703(.A(new_n790_), .B(new_n904_), .C1(new_n804_), .C2(new_n787_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n587_), .B1(new_n906_), .B2(new_n803_), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n901_), .B(new_n902_), .C1(new_n907_), .C2(new_n813_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(KEYINPUT126), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT126), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n850_), .A2(new_n910_), .A3(new_n902_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n438_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n833_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g715(.A(KEYINPUT63), .B(G211gat), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n910_), .B1(new_n850_), .B2(new_n902_), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n873_), .A2(KEYINPUT126), .A3(new_n383_), .A4(new_n869_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n587_), .B(new_n917_), .C1(new_n918_), .C2(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT127), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n662_), .B1(new_n909_), .B2(new_n911_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  OAI211_X1 g722(.A(new_n920_), .B(new_n921_), .C1(new_n922_), .C2(new_n923_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n587_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n923_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n921_), .B1(new_n928_), .B2(new_n920_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n925_), .A2(new_n929_), .ZN(G1354gat));
  INV_X1    g729(.A(new_n912_), .ZN(new_n931_));
  OAI21_X1  g730(.A(G218gat), .B1(new_n931_), .B2(new_n552_), .ZN(new_n932_));
  OR2_X1    g731(.A1(new_n627_), .A2(G218gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n931_), .B2(new_n933_), .ZN(G1355gat));
endmodule


