//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n786_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n936_,
    new_n937_, new_n939_, new_n940_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_;
  XOR2_X1   g000(.A(G85gat), .B(G92gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT8), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NOR3_X1   g005(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT7), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n206_), .B1(new_n209_), .B2(KEYINPUT67), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n207_), .B(KEYINPUT7), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n203_), .B1(new_n210_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n202_), .B1(new_n209_), .B2(new_n206_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT8), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n202_), .A2(KEYINPUT65), .ZN(new_n219_));
  INV_X1    g018(.A(G85gat), .ZN(new_n220_));
  INV_X1    g019(.A(G92gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT9), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n206_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT10), .B(G99gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n225_));
  OR3_X1    g024(.A1(new_n224_), .A2(new_n225_), .A3(G106gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n202_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n225_), .B1(new_n224_), .B2(G106gat), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n223_), .A2(new_n226_), .A3(new_n227_), .A4(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n215_), .A2(new_n218_), .A3(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(G29gat), .B(G36gat), .Z(new_n231_));
  XOR2_X1   g030(.A(G43gat), .B(G50gat), .Z(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT74), .B(KEYINPUT15), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n230_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n229_), .A2(new_n218_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(new_n214_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n233_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G232gat), .A2(G233gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(KEYINPUT35), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(KEYINPUT35), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT73), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT75), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n243_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n236_), .A2(new_n239_), .A3(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n246_), .A2(new_n247_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n250_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G190gat), .B(G218gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G134gat), .B(G162gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n256_), .A2(KEYINPUT36), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n256_), .B(KEYINPUT36), .Z(new_n259_));
  NAND3_X1  g058(.A1(new_n251_), .A2(new_n252_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n258_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT37), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT76), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n262_), .B1(new_n260_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n258_), .B(new_n260_), .C1(new_n263_), .C2(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G57gat), .B(G64gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT11), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT68), .B(G71gat), .ZN(new_n271_));
  INV_X1    g070(.A(G78gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n271_), .B(G78gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n269_), .A2(KEYINPUT11), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n238_), .A2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n278_), .B1(new_n237_), .B2(new_n214_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(KEYINPUT69), .ZN(new_n282_));
  AND2_X1   g081(.A1(G230gat), .A2(G233gat), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n282_), .B(new_n283_), .C1(KEYINPUT69), .C2(new_n281_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT12), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(new_n279_), .B2(KEYINPUT70), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT70), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n278_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n230_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n283_), .B1(new_n238_), .B2(new_n279_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n281_), .A2(new_n285_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n284_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G120gat), .B(G148gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT5), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G176gat), .B(G204gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n295_), .B(new_n296_), .Z(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT71), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n293_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n297_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n284_), .A2(new_n292_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(KEYINPUT13), .B1(new_n299_), .B2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n293_), .A2(new_n298_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT13), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n305_), .A3(new_n301_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n303_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G1gat), .B(G8gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT14), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT77), .B(G1gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(G8gat), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT78), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G15gat), .B(G22gat), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n309_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n315_), .A3(new_n309_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G231gat), .A2(G233gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n278_), .B(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n319_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G127gat), .B(G155gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT16), .ZN(new_n325_));
  XOR2_X1   g124(.A(G183gat), .B(G211gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(KEYINPUT70), .A3(KEYINPUT17), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n323_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n329_), .B1(KEYINPUT17), .B2(new_n328_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n322_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n268_), .A2(new_n308_), .A3(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G113gat), .B(G141gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G169gat), .B(G197gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n318_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n233_), .B1(new_n340_), .B2(new_n316_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n317_), .A2(new_n235_), .A3(new_n318_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G229gat), .A2(G233gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n233_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n317_), .A2(new_n346_), .A3(new_n318_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n343_), .B1(new_n341_), .B2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n339_), .B1(new_n345_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n341_), .A2(new_n347_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n343_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(new_n344_), .A3(new_n338_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(KEYINPUT79), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT79), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n355_), .B(new_n339_), .C1(new_n345_), .C2(new_n348_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G15gat), .B(G43gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT86), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT30), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT31), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT84), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT22), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(G169gat), .ZN(new_n366_));
  INV_X1    g165(.A(G169gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT22), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n364_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n364_), .B1(new_n367_), .B2(KEYINPUT22), .ZN(new_n370_));
  INV_X1    g169(.A(G176gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n363_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(G176gat), .B1(new_n366_), .B2(new_n364_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT22), .B(G169gat), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n374_), .B(KEYINPUT85), .C1(new_n364_), .C2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT23), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(KEYINPUT83), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT83), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT23), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  AND2_X1   g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n380_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(G183gat), .A2(G190gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n379_), .B1(new_n387_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n377_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT26), .ZN(new_n392_));
  INV_X1    g191(.A(G190gat), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n392_), .B1(new_n393_), .B2(KEYINPUT81), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT81), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n395_), .A2(KEYINPUT26), .A3(G190gat), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT80), .ZN(new_n398_));
  INV_X1    g197(.A(G183gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n398_), .B1(new_n399_), .B2(KEYINPUT25), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT25), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n401_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n399_), .A2(KEYINPUT25), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT82), .B1(new_n397_), .B2(new_n404_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n402_), .A2(new_n403_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT82), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n394_), .A2(new_n396_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .A4(new_n400_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(G169gat), .A2(G176gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(KEYINPUT24), .A3(new_n378_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT24), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G183gat), .A2(G190gat), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n416_), .A2(KEYINPUT23), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n382_), .A2(new_n384_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n418_), .B1(new_n419_), .B2(new_n386_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n405_), .A2(new_n409_), .A3(new_n415_), .A4(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n391_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G227gat), .A2(G233gat), .ZN(new_n423_));
  INV_X1    g222(.A(G71gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(G99gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n422_), .B(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(G127gat), .B(G134gat), .Z(new_n428_));
  XOR2_X1   g227(.A(G113gat), .B(G120gat), .Z(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n427_), .A2(new_n430_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n362_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n433_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(new_n361_), .A3(new_n431_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT87), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT29), .ZN(new_n440_));
  OR2_X1    g239(.A1(G141gat), .A2(G148gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G141gat), .A2(G148gat), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G155gat), .A2(G162gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT1), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT1), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(G155gat), .A3(G162gat), .ZN(new_n447_));
  OR2_X1    g246(.A1(G155gat), .A2(G162gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n445_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT88), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT88), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n443_), .A2(new_n449_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT89), .B1(G141gat), .B2(G148gat), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT3), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NOR3_X1   g256(.A1(KEYINPUT89), .A2(G141gat), .A3(G148gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT90), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G141gat), .A2(G148gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT89), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT90), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(new_n456_), .A4(new_n455_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n442_), .A2(KEYINPUT2), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT2), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(G141gat), .A3(G148gat), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n465_), .A2(new_n467_), .B1(new_n441_), .B2(KEYINPUT3), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n459_), .A2(new_n464_), .A3(new_n468_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n448_), .A2(new_n444_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT91), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n454_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n472_), .B1(new_n454_), .B2(new_n471_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n440_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G22gat), .B(G50gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n476_), .B(new_n477_), .Z(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT97), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n440_), .B(new_n478_), .C1(new_n473_), .C2(new_n474_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n480_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT94), .ZN(new_n484_));
  INV_X1    g283(.A(G197gat), .ZN(new_n485_));
  INV_X1    g284(.A(G204gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT93), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT93), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(G204gat), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n485_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(G197gat), .A2(G204gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n484_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n491_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT93), .B(G204gat), .ZN(new_n494_));
  OAI211_X1 g293(.A(KEYINPUT94), .B(new_n493_), .C1(new_n494_), .C2(new_n485_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(G211gat), .B(G218gat), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT21), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n492_), .A2(new_n495_), .A3(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n497_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n487_), .A2(new_n489_), .A3(new_n485_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n497_), .B1(G197gat), .B2(G204gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n500_), .A2(new_n503_), .A3(new_n496_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n499_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT96), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n504_), .A2(new_n499_), .A3(KEYINPUT96), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n454_), .A2(new_n471_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n509_), .B1(new_n440_), .B2(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(G228gat), .A2(G233gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n483_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n510_), .A2(KEYINPUT91), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n454_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(KEYINPUT29), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n505_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(new_n513_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n519_), .A2(KEYINPUT95), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT95), .B1(new_n519_), .B2(new_n521_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n517_), .A2(new_n518_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n478_), .B1(new_n526_), .B2(new_n440_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n482_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT97), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(G78gat), .B(G106gat), .Z(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n480_), .A2(new_n482_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n530_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n532_), .A2(KEYINPUT97), .A3(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n516_), .A2(new_n525_), .A3(new_n531_), .A4(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n532_), .B2(KEYINPUT97), .ZN(new_n536_));
  AOI211_X1 g335(.A(new_n481_), .B(new_n530_), .C1(new_n480_), .C2(new_n482_), .ZN(new_n537_));
  OAI22_X1  g336(.A1(new_n536_), .A2(new_n537_), .B1(new_n515_), .B2(new_n524_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n430_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n517_), .A2(new_n518_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(G225gat), .ZN(new_n542_));
  INV_X1    g341(.A(G233gat), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n430_), .A2(KEYINPUT101), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n430_), .A2(KEYINPUT101), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n511_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n541_), .A2(new_n545_), .A3(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G1gat), .B(G29gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(G85gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT0), .B(G57gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n541_), .A2(KEYINPUT4), .A3(new_n548_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT4), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n517_), .A2(new_n556_), .A3(new_n518_), .A4(new_n540_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n544_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n549_), .B(new_n554_), .C1(new_n555_), .C2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT33), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G226gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n366_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT99), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n565_), .A2(new_n566_), .A3(new_n378_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n417_), .B1(new_n385_), .B2(new_n416_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n567_), .B1(new_n568_), .B2(new_n388_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n566_), .B1(new_n565_), .B2(new_n378_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n401_), .A2(G183gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n403_), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT26), .B(G190gat), .Z(new_n573_));
  OAI21_X1  g372(.A(new_n387_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n412_), .A2(new_n414_), .ZN(new_n575_));
  OAI22_X1  g374(.A1(new_n569_), .A2(new_n570_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  OAI211_X1 g375(.A(KEYINPUT20), .B(new_n564_), .C1(new_n576_), .C2(new_n505_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT100), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n397_), .A2(new_n404_), .A3(KEYINPUT82), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n386_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n412_), .B(new_n414_), .C1(new_n580_), .C2(new_n417_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n582_), .A2(new_n405_), .B1(new_n377_), .B2(new_n390_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n578_), .B1(new_n583_), .B2(new_n520_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n422_), .A2(KEYINPUT100), .A3(new_n505_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n577_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT20), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n587_), .B1(new_n576_), .B2(new_n505_), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n391_), .A2(new_n421_), .A3(new_n504_), .A4(new_n499_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n564_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G8gat), .B(G36gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT18), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G64gat), .B(G92gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n586_), .A2(new_n590_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n594_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n564_), .A2(KEYINPUT20), .ZN(new_n597_));
  INV_X1    g396(.A(new_n576_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n598_), .B2(new_n520_), .ZN(new_n599_));
  AOI221_X4 g398(.A(new_n578_), .B1(new_n499_), .B2(new_n504_), .C1(new_n391_), .C2(new_n421_), .ZN(new_n600_));
  AOI21_X1  g399(.A(KEYINPUT100), .B1(new_n422_), .B2(new_n505_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n599_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n588_), .A2(new_n589_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n564_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n596_), .B1(new_n602_), .B2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n595_), .A2(new_n606_), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n541_), .A2(new_n548_), .A3(KEYINPUT4), .A4(new_n545_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n541_), .A2(new_n548_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n557_), .B(new_n608_), .C1(new_n609_), .C2(new_n545_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n553_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n541_), .A2(KEYINPUT4), .A3(new_n548_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(new_n544_), .A3(new_n557_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n613_), .A2(KEYINPUT33), .A3(new_n549_), .A4(new_n554_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n561_), .A2(new_n607_), .A3(new_n611_), .A4(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n596_), .A2(KEYINPUT32), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n598_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n618_), .A2(KEYINPUT20), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n584_), .A2(new_n585_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n564_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n588_), .A2(new_n564_), .A3(new_n589_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n617_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n602_), .A2(new_n605_), .A3(new_n616_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n559_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n554_), .B1(new_n613_), .B2(new_n549_), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n623_), .B(new_n624_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n539_), .B1(new_n615_), .B2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n602_), .A2(new_n605_), .A3(new_n596_), .ZN(new_n629_));
  OAI211_X1 g428(.A(KEYINPUT20), .B(new_n618_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n622_), .B1(new_n630_), .B2(new_n604_), .ZN(new_n631_));
  OAI211_X1 g430(.A(KEYINPUT27), .B(new_n629_), .C1(new_n631_), .C2(new_n596_), .ZN(new_n632_));
  XOR2_X1   g431(.A(KEYINPUT102), .B(KEYINPUT27), .Z(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n595_), .B2(new_n606_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n613_), .A2(new_n549_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n553_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n632_), .A2(new_n634_), .A3(new_n636_), .A4(new_n559_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n535_), .B2(new_n538_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n439_), .B1(new_n628_), .B2(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n535_), .A2(new_n538_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n625_), .A2(new_n626_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n632_), .A2(new_n634_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n640_), .A2(new_n641_), .A3(new_n437_), .A4(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n357_), .B1(new_n639_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n335_), .A2(new_n645_), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n646_), .A2(new_n641_), .A3(new_n311_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT38), .Z(new_n648_));
  NAND2_X1  g447(.A1(new_n639_), .A2(new_n644_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n261_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT103), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(KEYINPUT103), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n649_), .A2(KEYINPUT104), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT104), .B1(new_n649_), .B2(new_n653_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n357_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n307_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n334_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n657_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G1gat), .B1(new_n661_), .B2(new_n641_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n648_), .A2(new_n662_), .ZN(G1324gat));
  INV_X1    g462(.A(G8gat), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n645_), .A2(new_n335_), .A3(new_n664_), .A4(new_n642_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT105), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n642_), .B(new_n660_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT39), .ZN(new_n668_));
  AND4_X1   g467(.A1(new_n666_), .A2(new_n667_), .A3(new_n668_), .A4(G8gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n664_), .B1(KEYINPUT105), .B2(KEYINPUT39), .ZN(new_n670_));
  AOI22_X1  g469(.A1(new_n667_), .A2(new_n670_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n665_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(KEYINPUT40), .B(new_n665_), .C1(new_n669_), .C2(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1325gat));
  OR3_X1    g475(.A1(new_n646_), .A2(G15gat), .A3(new_n439_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n657_), .A2(new_n438_), .A3(new_n660_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n678_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT41), .B1(new_n678_), .B2(G15gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n677_), .B1(new_n679_), .B2(new_n680_), .ZN(G1326gat));
  OR3_X1    g480(.A1(new_n646_), .A2(G22gat), .A3(new_n640_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n657_), .A2(new_n539_), .A3(new_n660_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(G22gat), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n683_), .B2(G22gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(G1327gat));
  NOR2_X1   g486(.A1(new_n261_), .A2(new_n333_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n307_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n645_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n641_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G29gat), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n615_), .A2(new_n627_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n640_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n643_), .A2(new_n539_), .A3(new_n641_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n438_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n644_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n694_), .B(new_n268_), .C1(new_n698_), .C2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n267_), .B1(new_n639_), .B2(new_n644_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n700_), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n659_), .A2(new_n333_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(KEYINPUT44), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT44), .B1(new_n703_), .B2(new_n704_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n692_), .A2(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n693_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  AOI21_X1  g508(.A(KEYINPUT109), .B1(KEYINPUT110), .B2(KEYINPUT46), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n703_), .A2(new_n704_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n703_), .A2(KEYINPUT44), .A3(new_n704_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n642_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(G36gat), .ZN(new_n716_));
  INV_X1    g515(.A(G36gat), .ZN(new_n717_));
  OR2_X1    g516(.A1(new_n642_), .A2(KEYINPUT108), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n642_), .A2(KEYINPUT108), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  AND4_X1   g519(.A1(new_n717_), .A2(new_n645_), .A3(new_n689_), .A4(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT45), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n721_), .B(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n710_), .B1(new_n716_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n705_), .A2(new_n706_), .A3(new_n643_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n725_), .B(new_n723_), .C1(new_n726_), .C2(new_n717_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT110), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n724_), .B1(new_n728_), .B2(new_n729_), .ZN(G1329gat));
  INV_X1    g529(.A(new_n437_), .ZN(new_n731_));
  INV_X1    g530(.A(G43gat), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n707_), .A2(KEYINPUT111), .A3(new_n733_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n713_), .A2(new_n714_), .A3(new_n733_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT111), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n732_), .B1(new_n690_), .B2(new_n439_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n734_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n734_), .A2(new_n737_), .A3(new_n738_), .A4(new_n740_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1330gat));
  NOR3_X1   g543(.A1(new_n705_), .A2(new_n706_), .A3(new_n640_), .ZN(new_n745_));
  INV_X1    g544(.A(G50gat), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n539_), .A2(new_n746_), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT113), .Z(new_n748_));
  OAI22_X1  g547(.A1(new_n745_), .A2(new_n746_), .B1(new_n690_), .B2(new_n748_), .ZN(G1331gat));
  NOR3_X1   g548(.A1(new_n307_), .A2(new_n334_), .A3(new_n658_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n657_), .A2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G57gat), .B1(new_n751_), .B2(new_n641_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n307_), .A2(new_n658_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n649_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n333_), .A3(new_n267_), .ZN(new_n755_));
  OR3_X1    g554(.A1(new_n755_), .A2(G57gat), .A3(new_n641_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n752_), .A2(new_n756_), .ZN(G1332gat));
  INV_X1    g556(.A(new_n720_), .ZN(new_n758_));
  OR3_X1    g557(.A1(new_n755_), .A2(G64gat), .A3(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G64gat), .B1(new_n751_), .B2(new_n758_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n760_), .A2(KEYINPUT48), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n760_), .A2(KEYINPUT48), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n759_), .B1(new_n761_), .B2(new_n762_), .ZN(G1333gat));
  OR3_X1    g562(.A1(new_n755_), .A2(G71gat), .A3(new_n439_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n438_), .B(new_n750_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n765_));
  XOR2_X1   g564(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(G71gat), .A3(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(G71gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT115), .ZN(G1334gat));
  OAI21_X1  g569(.A(G78gat), .B1(new_n751_), .B2(new_n640_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n771_), .A2(KEYINPUT50), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(KEYINPUT50), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n539_), .A2(new_n272_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT116), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n772_), .A2(new_n773_), .B1(new_n755_), .B2(new_n775_), .ZN(G1335gat));
  NAND2_X1  g575(.A1(new_n754_), .A2(new_n688_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n220_), .B1(new_n777_), .B2(new_n641_), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT117), .Z(new_n779_));
  AND3_X1   g578(.A1(new_n703_), .A2(new_n334_), .A3(new_n753_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n781_), .A2(new_n220_), .A3(new_n641_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n779_), .A2(new_n782_), .ZN(G1336gat));
  OAI21_X1  g582(.A(G92gat), .B1(new_n781_), .B2(new_n758_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n777_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(new_n221_), .A3(new_n642_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1337gat));
  INV_X1    g586(.A(G99gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n788_), .B1(new_n780_), .B2(new_n438_), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n777_), .A2(new_n224_), .A3(new_n731_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791_));
  OAI22_X1  g590(.A1(new_n789_), .A2(new_n790_), .B1(new_n791_), .B2(KEYINPUT51), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(KEYINPUT51), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(G1338gat));
  OR3_X1    g593(.A1(new_n777_), .A2(G106gat), .A3(new_n640_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n703_), .A2(new_n539_), .A3(new_n334_), .A4(new_n753_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n796_), .A2(new_n797_), .A3(G106gat), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n796_), .B2(G106gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g600(.A1(new_n267_), .A2(new_n307_), .A3(new_n333_), .A4(new_n357_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n802_), .B(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n292_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n289_), .A2(new_n291_), .A3(new_n280_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(new_n283_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n289_), .A2(new_n290_), .A3(KEYINPUT55), .A4(new_n291_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n298_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n810_), .A2(KEYINPUT56), .A3(new_n298_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n813_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT56), .B1(new_n810_), .B2(new_n298_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT120), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n350_), .A2(new_n343_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n341_), .A2(new_n342_), .A3(new_n351_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n339_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n353_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n302_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n816_), .A2(new_n818_), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n816_), .A2(KEYINPUT58), .A3(new_n818_), .A4(new_n823_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n268_), .A3(new_n827_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n354_), .A2(new_n356_), .A3(new_n301_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n815_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n817_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n822_), .B1(new_n304_), .B2(new_n301_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n650_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT119), .B1(new_n834_), .B2(KEYINPUT57), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n354_), .A2(new_n356_), .A3(new_n301_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n261_), .B1(new_n837_), .B2(new_n832_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n834_), .A2(KEYINPUT57), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n828_), .A2(new_n835_), .A3(new_n841_), .A4(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n804_), .B1(new_n843_), .B2(new_n334_), .ZN(new_n844_));
  NOR4_X1   g643(.A1(new_n539_), .A2(new_n642_), .A3(new_n731_), .A4(new_n641_), .ZN(new_n845_));
  XOR2_X1   g644(.A(new_n845_), .B(KEYINPUT121), .Z(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n844_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(G113gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n658_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n838_), .A2(new_n840_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n828_), .A2(new_n842_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n334_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n804_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n856_), .A3(new_n846_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT59), .B1(new_n844_), .B2(new_n847_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n857_), .A2(new_n858_), .A3(new_n658_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n850_), .B1(new_n859_), .B2(new_n849_), .ZN(G1340gat));
  NAND2_X1  g659(.A1(new_n843_), .A2(new_n334_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n854_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n856_), .B1(new_n862_), .B2(new_n846_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n804_), .B1(new_n334_), .B2(new_n852_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n846_), .A2(new_n856_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n308_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT122), .B1(new_n863_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT122), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n857_), .A2(new_n858_), .A3(new_n868_), .A4(new_n308_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n867_), .A2(G120gat), .A3(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n307_), .B2(KEYINPUT60), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n848_), .B(new_n872_), .C1(KEYINPUT60), .C2(new_n871_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(G1341gat));
  INV_X1    g673(.A(G127gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n848_), .A2(new_n875_), .A3(new_n333_), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n857_), .A2(new_n858_), .A3(new_n333_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n875_), .ZN(G1342gat));
  INV_X1    g677(.A(G134gat), .ZN(new_n879_));
  INV_X1    g678(.A(new_n653_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n848_), .A2(new_n879_), .A3(new_n880_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n857_), .A2(new_n858_), .A3(new_n268_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(new_n879_), .ZN(G1343gat));
  NOR2_X1   g682(.A1(new_n438_), .A2(new_n640_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n885_), .A2(new_n720_), .A3(new_n641_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n844_), .A2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(new_n658_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n308_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g691(.A1(new_n862_), .A2(new_n333_), .A3(new_n886_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT123), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n888_), .A2(KEYINPUT123), .A3(new_n333_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(KEYINPUT61), .B(G155gat), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n895_), .A2(new_n896_), .A3(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n895_), .B2(new_n896_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1346gat));
  NAND2_X1  g699(.A1(new_n862_), .A2(new_n886_), .ZN(new_n901_));
  OAI21_X1  g700(.A(G162gat), .B1(new_n901_), .B2(new_n267_), .ZN(new_n902_));
  INV_X1    g701(.A(G162gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n880_), .A2(new_n903_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n902_), .B(KEYINPUT124), .C1(new_n901_), .C2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT124), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n901_), .A2(new_n904_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n903_), .B1(new_n888_), .B2(new_n268_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n905_), .A2(new_n909_), .ZN(G1347gat));
  XNOR2_X1  g709(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n720_), .A2(new_n641_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n439_), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n855_), .A2(new_n640_), .A3(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n357_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n911_), .B1(new_n915_), .B2(new_n367_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n911_), .ZN(new_n917_));
  OAI211_X1 g716(.A(G169gat), .B(new_n917_), .C1(new_n914_), .C2(new_n357_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n915_), .A2(new_n375_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n916_), .A2(new_n918_), .A3(new_n919_), .ZN(G1348gat));
  INV_X1    g719(.A(new_n914_), .ZN(new_n921_));
  AOI21_X1  g720(.A(G176gat), .B1(new_n921_), .B2(new_n308_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n844_), .A2(new_n539_), .ZN(new_n923_));
  NOR4_X1   g722(.A1(new_n912_), .A2(new_n371_), .A3(new_n307_), .A4(new_n439_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1349gat));
  INV_X1    g724(.A(KEYINPUT126), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n913_), .A2(new_n333_), .ZN(new_n927_));
  NOR3_X1   g726(.A1(new_n844_), .A2(new_n539_), .A3(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(G183gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n855_), .A2(new_n640_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n913_), .A2(new_n572_), .A3(new_n333_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n926_), .B1(new_n929_), .B2(new_n932_), .ZN(new_n933_));
  OAI221_X1 g732(.A(KEYINPUT126), .B1(new_n930_), .B2(new_n931_), .C1(new_n928_), .C2(G183gat), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1350gat));
  OAI21_X1  g734(.A(G190gat), .B1(new_n914_), .B2(new_n267_), .ZN(new_n936_));
  OR2_X1    g735(.A1(new_n653_), .A2(new_n573_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n914_), .B2(new_n937_), .ZN(G1351gat));
  NOR3_X1   g737(.A1(new_n844_), .A2(new_n885_), .A3(new_n912_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n658_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n308_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n494_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n943_), .B1(new_n486_), .B2(new_n942_), .ZN(G1353gat));
  INV_X1    g743(.A(KEYINPUT63), .ZN(new_n945_));
  INV_X1    g744(.A(G211gat), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n945_), .A2(new_n946_), .A3(KEYINPUT127), .ZN(new_n947_));
  NAND2_X1  g746(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n939_), .A2(new_n333_), .A3(new_n947_), .A4(new_n948_), .ZN(new_n949_));
  AOI21_X1  g748(.A(KEYINPUT127), .B1(new_n945_), .B2(new_n946_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n949_), .B(new_n950_), .ZN(G1354gat));
  NAND4_X1  g750(.A1(new_n862_), .A2(new_n641_), .A3(new_n720_), .A4(new_n884_), .ZN(new_n952_));
  OR3_X1    g751(.A1(new_n952_), .A2(G218gat), .A3(new_n653_), .ZN(new_n953_));
  OAI21_X1  g752(.A(G218gat), .B1(new_n952_), .B2(new_n267_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(G1355gat));
endmodule


