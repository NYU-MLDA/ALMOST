//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_;
  XNOR2_X1  g000(.A(KEYINPUT25), .B(G183gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT83), .ZN(new_n203_));
  INV_X1    g002(.A(G190gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT26), .B1(new_n203_), .B2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT26), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G190gat), .ZN(new_n207_));
  OAI211_X1 g006(.A(new_n202_), .B(new_n205_), .C1(new_n203_), .C2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(G183gat), .A3(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  AND3_X1   g010(.A1(new_n211_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT84), .B1(new_n211_), .B2(KEYINPUT23), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n210_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NOR3_X1   g013(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n215_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n208_), .A2(new_n214_), .A3(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n211_), .A2(KEYINPUT23), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT86), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT86), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n211_), .A2(new_n224_), .A3(KEYINPUT23), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n221_), .B1(new_n226_), .B2(new_n210_), .ZN(new_n227_));
  INV_X1    g026(.A(G169gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT22), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT22), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G169gat), .ZN(new_n231_));
  INV_X1    g030(.A(G176gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n229_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT85), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G169gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(KEYINPUT85), .A3(new_n232_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n237_), .A3(new_n218_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n220_), .B1(new_n227_), .B2(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(G71gat), .B(G99gat), .Z(new_n240_));
  XNOR2_X1  g039(.A(G15gat), .B(G43gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n239_), .B(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G227gat), .A2(G233gat), .ZN(new_n244_));
  XOR2_X1   g043(.A(new_n244_), .B(KEYINPUT87), .Z(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT30), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n243_), .B(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT88), .ZN(new_n248_));
  INV_X1    g047(.A(G134gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G127gat), .ZN(new_n250_));
  INV_X1    g049(.A(G127gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G134gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(G120gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G113gat), .ZN(new_n255_));
  INV_X1    g054(.A(G113gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G120gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n250_), .A2(new_n252_), .A3(new_n255_), .A4(new_n257_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n261_), .B(KEYINPUT31), .Z(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n247_), .A2(new_n248_), .A3(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n247_), .A2(new_n248_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n262_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(G197gat), .A2(G204gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G197gat), .A2(G204gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(KEYINPUT21), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT21), .ZN(new_n271_));
  AND2_X1   g070(.A1(G197gat), .A2(G204gat), .ZN(new_n272_));
  NOR2_X1   g071(.A1(G197gat), .A2(G204gat), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n271_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G211gat), .B(G218gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n270_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NOR3_X1   g075(.A1(new_n272_), .A2(new_n273_), .A3(new_n271_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G211gat), .B(G218gat), .Z(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G141gat), .ZN(new_n281_));
  INV_X1    g080(.A(G148gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(new_n282_), .A3(KEYINPUT89), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT3), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT3), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(KEYINPUT89), .A3(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G141gat), .A2(G148gat), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT2), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n291_));
  NAND4_X1  g090(.A1(new_n284_), .A2(new_n287_), .A3(new_n290_), .A4(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(G155gat), .B(G162gat), .Z(new_n293_));
  INV_X1    g092(.A(KEYINPUT1), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n285_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n288_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n292_), .A2(new_n293_), .B1(new_n295_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT29), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n280_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(KEYINPUT91), .A2(G233gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(KEYINPUT91), .A2(G233gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(G228gat), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n302_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT90), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n309_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n293_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n290_), .A2(new_n291_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n286_), .B1(new_n285_), .B2(KEYINPUT89), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n311_), .B1(new_n314_), .B2(new_n287_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n298_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n316_));
  OAI211_X1 g115(.A(KEYINPUT90), .B(KEYINPUT29), .C1(new_n315_), .C2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n310_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n280_), .A2(new_n306_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT92), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT92), .ZN(new_n322_));
  AOI211_X1 g121(.A(new_n322_), .B(new_n319_), .C1(new_n310_), .C2(new_n317_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n308_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  XOR2_X1   g123(.A(G78gat), .B(G106gat), .Z(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n325_), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n327_), .B(new_n308_), .C1(new_n321_), .C2(new_n323_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n300_), .A2(new_n301_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT28), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G22gat), .B(G50gat), .Z(new_n333_));
  AND2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n332_), .A2(new_n333_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n329_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n326_), .A2(new_n336_), .A3(new_n328_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G183gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT25), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT25), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(G183gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n204_), .A2(KEYINPUT26), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n342_), .A2(new_n344_), .A3(new_n207_), .A4(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n219_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n210_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n348_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n233_), .A2(new_n218_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n221_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n351_), .B1(new_n214_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n280_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n218_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n355_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n237_), .B(new_n356_), .C1(new_n349_), .C2(new_n221_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n276_), .A2(new_n279_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(new_n358_), .A3(new_n220_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n354_), .A2(new_n359_), .A3(KEYINPUT20), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT19), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n239_), .A2(new_n280_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n353_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n226_), .A2(new_n210_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n366_), .A2(new_n219_), .A3(new_n346_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n365_), .A2(new_n358_), .A3(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n362_), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n364_), .A2(new_n368_), .A3(KEYINPUT20), .A4(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n370_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G8gat), .B(G36gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT18), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n371_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n363_), .A2(new_n375_), .A3(new_n370_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT93), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n259_), .A2(new_n260_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n380_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n292_), .A2(new_n293_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n295_), .A2(new_n299_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(KEYINPUT94), .B1(new_n383_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT94), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n300_), .B(new_n389_), .C1(new_n382_), .C2(new_n381_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n261_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  OR3_X1    g192(.A1(new_n388_), .A2(new_n393_), .A3(KEYINPUT96), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT96), .B1(new_n388_), .B2(new_n393_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n394_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G1gat), .B(G29gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(G85gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT0), .B(G57gat), .ZN(new_n401_));
  XOR2_X1   g200(.A(new_n400_), .B(new_n401_), .Z(new_n402_));
  NAND4_X1  g201(.A1(new_n387_), .A2(KEYINPUT4), .A3(new_n392_), .A4(new_n390_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n392_), .A2(KEYINPUT4), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n402_), .B1(new_n405_), .B2(new_n395_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n379_), .B1(new_n398_), .B2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n403_), .A2(new_n396_), .A3(new_n404_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n387_), .A2(new_n395_), .A3(new_n392_), .A4(new_n390_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n409_), .A3(new_n402_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT95), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(KEYINPUT33), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT95), .B1(new_n410_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n410_), .A2(new_n414_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n407_), .A2(new_n413_), .A3(new_n415_), .A4(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n375_), .A2(KEYINPUT32), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n363_), .A2(new_n418_), .A3(new_n370_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT20), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n420_), .B1(new_n239_), .B2(new_n280_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n369_), .B1(new_n421_), .B2(new_n368_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n354_), .A2(new_n359_), .A3(KEYINPUT20), .A4(new_n369_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n402_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n426_));
  OAI221_X1 g225(.A(new_n419_), .B1(new_n418_), .B2(new_n425_), .C1(new_n411_), .C2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n340_), .B1(new_n417_), .B2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n411_), .A2(new_n426_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n326_), .A2(new_n336_), .A3(new_n328_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n336_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n429_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n378_), .A2(KEYINPUT27), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n364_), .A2(KEYINPUT20), .A3(new_n368_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n362_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n375_), .B1(new_n435_), .B2(new_n423_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT97), .B1(new_n433_), .B2(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n376_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT97), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n438_), .A2(new_n439_), .A3(KEYINPUT27), .A4(new_n378_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT27), .ZN(new_n442_));
  AOI21_X1  g241(.A(KEYINPUT98), .B1(new_n379_), .B2(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n363_), .A2(new_n375_), .A3(new_n370_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n375_), .B1(new_n363_), .B2(new_n370_), .ZN(new_n445_));
  OAI211_X1 g244(.A(KEYINPUT98), .B(new_n442_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n441_), .B1(new_n443_), .B2(new_n447_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n432_), .A2(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n267_), .B1(new_n428_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n340_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n429_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n267_), .A2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n442_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT98), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(new_n446_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT99), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n457_), .A2(new_n458_), .A3(new_n441_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n457_), .B2(new_n441_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n451_), .B(new_n453_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n450_), .A2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G29gat), .B(G36gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G43gat), .B(G50gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(KEYINPUT82), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G15gat), .B(G22gat), .ZN(new_n467_));
  INV_X1    g266(.A(G1gat), .ZN(new_n468_));
  INV_X1    g267(.A(G8gat), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT14), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G1gat), .B(G8gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n466_), .B(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G229gat), .A2(G233gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n466_), .A2(new_n473_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT81), .B(KEYINPUT15), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n465_), .B(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n473_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n481_), .A3(new_n475_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n477_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G113gat), .B(G141gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G169gat), .B(G197gat), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n484_), .B(new_n485_), .Z(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n477_), .A2(new_n482_), .A3(new_n486_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n462_), .A2(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n491_), .A2(KEYINPUT100), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(KEYINPUT100), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT68), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT7), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n495_), .B(new_n496_), .C1(G99gat), .C2(G106gat), .ZN(new_n497_));
  INV_X1    g296(.A(G99gat), .ZN(new_n498_));
  INV_X1    g297(.A(G106gat), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n498_), .B(new_n499_), .C1(KEYINPUT68), .C2(KEYINPUT7), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT71), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n497_), .A2(new_n500_), .A3(KEYINPUT71), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G99gat), .A2(G106gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT6), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(G99gat), .A3(G106gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT70), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n506_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(new_n508_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT70), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n503_), .A2(new_n504_), .A3(new_n510_), .A4(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT8), .ZN(new_n514_));
  INV_X1    g313(.A(G85gat), .ZN(new_n515_));
  INV_X1    g314(.A(G92gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT69), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n517_), .A2(KEYINPUT69), .A3(new_n518_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n514_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n513_), .A2(new_n523_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n521_), .A2(new_n522_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n501_), .A2(new_n511_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n514_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  OR2_X1    g326(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n528_), .A2(KEYINPUT65), .A3(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT65), .B1(new_n528_), .B2(new_n529_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n499_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  OAI211_X1 g331(.A(KEYINPUT66), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n533_), .A2(KEYINPUT67), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(KEYINPUT67), .ZN(new_n535_));
  NOR2_X1   g334(.A1(KEYINPUT66), .A2(KEYINPUT9), .ZN(new_n536_));
  OAI22_X1  g335(.A1(new_n534_), .A2(new_n535_), .B1(new_n518_), .B2(new_n536_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n533_), .A2(KEYINPUT67), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n536_), .A2(new_n518_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n533_), .A2(KEYINPUT67), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n532_), .A2(new_n537_), .A3(new_n511_), .A4(new_n541_), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n524_), .A2(new_n527_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n465_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n524_), .A2(new_n527_), .A3(new_n542_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n480_), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT79), .B(KEYINPUT34), .Z(new_n547_));
  NAND2_X1  g346(.A1(G232gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n549_), .A2(KEYINPUT35), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n544_), .A2(new_n546_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n549_), .A2(KEYINPUT35), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(KEYINPUT80), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n551_), .B(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G190gat), .B(G218gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT36), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n554_), .A2(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n557_), .A2(KEYINPUT36), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n554_), .A2(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n559_), .A2(KEYINPUT37), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT37), .B1(new_n559_), .B2(new_n561_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(G64gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(G57gat), .ZN(new_n567_));
  INV_X1    g366(.A(G57gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(G64gat), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n567_), .A2(new_n569_), .A3(KEYINPUT72), .ZN(new_n570_));
  AOI21_X1  g369(.A(KEYINPUT72), .B1(new_n567_), .B2(new_n569_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT11), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT72), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n568_), .A2(G64gat), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n566_), .A2(G57gat), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT11), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n567_), .A2(new_n569_), .A3(KEYINPUT72), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G71gat), .B(G78gat), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n572_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  OAI211_X1 g381(.A(KEYINPUT11), .B(new_n580_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n582_), .A2(new_n585_), .A3(new_n583_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G231gat), .A2(G233gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n473_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n589_), .B(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(G127gat), .B(G155gat), .Z(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT16), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G183gat), .B(G211gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT17), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n596_), .A2(new_n597_), .ZN(new_n599_));
  OR3_X1    g398(.A1(new_n592_), .A2(new_n598_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n592_), .A2(new_n598_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n565_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT77), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT75), .B1(new_n589_), .B2(new_n545_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n582_), .A2(new_n585_), .A3(new_n583_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n585_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT75), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n609_), .A2(new_n610_), .A3(new_n543_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n545_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n606_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(G230gat), .A2(G233gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT64), .Z(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(KEYINPUT12), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT12), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n545_), .B(new_n617_), .C1(new_n607_), .C2(new_n608_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n615_), .B1(new_n609_), .B2(new_n543_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n613_), .A2(new_n615_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  XOR2_X1   g420(.A(G120gat), .B(G148gat), .Z(new_n622_));
  XNOR2_X1  g421(.A(G176gat), .B(G204gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(KEYINPUT76), .B(KEYINPUT5), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n624_), .B(new_n625_), .Z(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n605_), .B1(new_n621_), .B2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n613_), .A2(new_n615_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n617_), .B1(new_n589_), .B2(new_n545_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n618_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n620_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n629_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n626_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n628_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n633_), .A2(new_n605_), .A3(new_n626_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT13), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n635_), .A2(KEYINPUT13), .A3(new_n636_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(KEYINPUT78), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT78), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n635_), .A2(KEYINPUT13), .A3(new_n636_), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n642_), .B2(new_n637_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n604_), .A2(new_n644_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n494_), .A2(new_n468_), .A3(new_n452_), .A4(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n647_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n490_), .B1(new_n642_), .B2(new_n637_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n602_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n559_), .A2(new_n561_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n450_), .B2(new_n461_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n650_), .A2(new_n651_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n652_), .A2(new_n653_), .A3(new_n656_), .A4(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G1gat), .B1(new_n658_), .B2(new_n429_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n648_), .A2(new_n649_), .A3(new_n659_), .ZN(G1324gat));
  NOR2_X1   g459(.A1(new_n459_), .A2(new_n460_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G8gat), .B1(new_n658_), .B2(new_n662_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n663_), .A2(KEYINPUT103), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(KEYINPUT103), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(KEYINPUT39), .A3(new_n665_), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n665_), .A2(KEYINPUT39), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n494_), .A2(new_n469_), .A3(new_n661_), .A4(new_n645_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n666_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n666_), .A2(new_n667_), .A3(KEYINPUT40), .A4(new_n668_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(G1325gat));
  INV_X1    g472(.A(new_n658_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n267_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT41), .B1(new_n676_), .B2(G15gat), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n494_), .A2(new_n645_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n267_), .A2(G15gat), .ZN(new_n681_));
  OAI22_X1  g480(.A1(new_n678_), .A2(new_n679_), .B1(new_n680_), .B2(new_n681_), .ZN(G1326gat));
  NAND2_X1  g481(.A1(new_n674_), .A2(new_n340_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n683_), .A2(new_n684_), .A3(G22gat), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(new_n683_), .B2(G22gat), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n451_), .A2(G22gat), .ZN(new_n688_));
  OAI22_X1  g487(.A1(new_n686_), .A2(new_n687_), .B1(new_n680_), .B2(new_n688_), .ZN(G1327gat));
  NOR2_X1   g488(.A1(new_n654_), .A2(new_n653_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT106), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n642_), .A2(new_n637_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n494_), .A2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n429_), .A2(G29gat), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT107), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n462_), .A2(new_n565_), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n462_), .A2(new_n702_), .A3(new_n565_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n652_), .A2(new_n602_), .A3(new_n657_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n704_), .A2(new_n705_), .A3(KEYINPUT44), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT44), .B1(new_n704_), .B2(new_n705_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(KEYINPUT105), .A3(new_n452_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G29gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(KEYINPUT105), .B1(new_n708_), .B2(new_n452_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n698_), .B1(new_n710_), .B2(new_n711_), .ZN(G1328gat));
  NOR2_X1   g511(.A1(new_n662_), .A2(G36gat), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n694_), .B(new_n713_), .C1(new_n492_), .C2(new_n493_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT45), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n706_), .A2(new_n707_), .A3(new_n662_), .ZN(new_n716_));
  INV_X1    g515(.A(G36gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n715_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(G1329gat));
  INV_X1    g519(.A(G43gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n695_), .A2(new_n721_), .A3(new_n675_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n706_), .A2(new_n707_), .A3(new_n267_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n723_), .B2(new_n721_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n722_), .B(KEYINPUT47), .C1(new_n723_), .C2(new_n721_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1330gat));
  INV_X1    g527(.A(G50gat), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n340_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT108), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n695_), .A2(new_n731_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n706_), .A2(new_n707_), .A3(new_n451_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n729_), .ZN(G1331gat));
  NOR2_X1   g533(.A1(new_n602_), .A2(new_n490_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n644_), .A2(new_n656_), .A3(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  OAI21_X1  g536(.A(G57gat), .B1(new_n737_), .B2(new_n429_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n490_), .B1(new_n450_), .B2(new_n461_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NOR3_X1   g539(.A1(new_n740_), .A2(new_n604_), .A3(new_n693_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(new_n568_), .A3(new_n452_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n742_), .ZN(G1332gat));
  AOI21_X1  g542(.A(new_n566_), .B1(new_n736_), .B2(new_n661_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n741_), .A2(new_n566_), .A3(new_n661_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1333gat));
  INV_X1    g547(.A(G71gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n741_), .A2(new_n749_), .A3(new_n675_), .ZN(new_n750_));
  OAI21_X1  g549(.A(G71gat), .B1(new_n737_), .B2(new_n267_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n751_), .A2(KEYINPUT49), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n751_), .A2(KEYINPUT49), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n750_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT110), .ZN(G1334gat));
  INV_X1    g554(.A(G78gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n736_), .B2(new_n340_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT50), .Z(new_n758_));
  NAND3_X1  g557(.A1(new_n741_), .A2(new_n756_), .A3(new_n340_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1335gat));
  NAND2_X1  g559(.A1(new_n644_), .A2(new_n691_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n761_), .A2(new_n740_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n515_), .A3(new_n452_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n693_), .A2(new_n490_), .A3(new_n653_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(new_n452_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n767_), .B2(new_n515_), .ZN(G1336gat));
  AOI21_X1  g567(.A(new_n516_), .B1(new_n766_), .B2(new_n661_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n662_), .A2(G92gat), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n762_), .B2(new_n770_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT111), .Z(G1337gat));
  OAI21_X1  g571(.A(new_n675_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  AND4_X1   g573(.A1(new_n644_), .A2(new_n739_), .A3(new_n691_), .A4(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n700_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n462_), .B2(new_n565_), .ZN(new_n777_));
  AOI211_X1 g576(.A(KEYINPUT43), .B(new_n564_), .C1(new_n450_), .C2(new_n461_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n675_), .B(new_n764_), .C1(new_n777_), .C2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n775_), .B1(new_n779_), .B2(G99gat), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT51), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT113), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(G99gat), .ZN(new_n783_));
  INV_X1    g582(.A(new_n775_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT112), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n781_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  AOI211_X1 g586(.A(new_n786_), .B(new_n775_), .C1(new_n779_), .C2(G99gat), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n782_), .B1(new_n787_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT51), .B1(new_n780_), .B2(KEYINPUT112), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n791_), .A2(KEYINPUT113), .A3(new_n788_), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT114), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n782_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(new_n788_), .B2(new_n791_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n787_), .A2(new_n796_), .A3(new_n789_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT114), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n795_), .A2(new_n797_), .A3(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n793_), .A2(new_n799_), .ZN(G1338gat));
  NAND3_X1  g599(.A1(new_n762_), .A2(new_n499_), .A3(new_n340_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n766_), .A2(new_n340_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(G106gat), .ZN(new_n804_));
  AOI211_X1 g603(.A(KEYINPUT52), .B(new_n499_), .C1(new_n766_), .C2(new_n340_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n801_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT53), .ZN(G1339gat));
  OAI211_X1 g606(.A(new_n564_), .B(new_n735_), .C1(new_n642_), .C2(new_n637_), .ZN(new_n808_));
  XOR2_X1   g607(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n810_), .A2(KEYINPUT116), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n808_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n808_), .A2(new_n811_), .ZN(new_n813_));
  AOI22_X1  g612(.A1(new_n812_), .A2(new_n813_), .B1(KEYINPUT116), .B2(new_n810_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n490_), .B1(new_n633_), .B2(new_n626_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n630_), .A2(new_n631_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n606_), .A2(new_n611_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n615_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n819_), .B(new_n620_), .C1(new_n630_), .C2(new_n631_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n819_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n818_), .B(KEYINPUT117), .C1(new_n821_), .C2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n632_), .A2(KEYINPUT55), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n820_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT117), .B1(new_n826_), .B2(new_n818_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n626_), .B1(new_n824_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n818_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n823_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(KEYINPUT56), .A3(new_n626_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n815_), .B1(new_n830_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n474_), .A2(new_n475_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n478_), .A2(new_n481_), .A3(new_n476_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n487_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n489_), .A2(new_n839_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT118), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n841_), .A2(new_n636_), .A3(new_n635_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n654_), .B1(new_n836_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT57), .B(new_n654_), .C1(new_n836_), .C2(new_n842_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n841_), .B1(new_n633_), .B2(new_n626_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT56), .B1(new_n834_), .B2(new_n626_), .ZN(new_n849_));
  AOI211_X1 g648(.A(new_n829_), .B(new_n627_), .C1(new_n833_), .C2(new_n823_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n848_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT58), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n848_), .B(KEYINPUT58), .C1(new_n849_), .C2(new_n850_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n565_), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n845_), .A2(new_n846_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n814_), .B1(new_n856_), .B2(new_n602_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NOR4_X1   g657(.A1(new_n661_), .A2(new_n429_), .A3(new_n340_), .A4(new_n267_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(G113gat), .B1(new_n860_), .B2(new_n490_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n847_), .B1(new_n830_), .B2(new_n835_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n564_), .B1(new_n862_), .B2(KEYINPUT58), .ZN(new_n863_));
  AOI22_X1  g662(.A1(new_n844_), .A2(new_n843_), .B1(new_n863_), .B2(new_n853_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n653_), .B1(new_n864_), .B2(new_n846_), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT119), .B(new_n859_), .C1(new_n865_), .C2(new_n814_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT59), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n858_), .A2(KEYINPUT119), .A3(KEYINPUT59), .A4(new_n859_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n256_), .B1(new_n490_), .B2(KEYINPUT120), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(KEYINPUT120), .B2(new_n256_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n861_), .B1(new_n870_), .B2(new_n872_), .ZN(G1340gat));
  OAI21_X1  g672(.A(new_n254_), .B1(new_n693_), .B2(KEYINPUT60), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n860_), .B(new_n874_), .C1(KEYINPUT60), .C2(new_n254_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n644_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n875_), .B1(new_n877_), .B2(new_n254_), .ZN(G1341gat));
  AOI21_X1  g677(.A(G127gat), .B1(new_n860_), .B2(new_n653_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n602_), .A2(KEYINPUT121), .ZN(new_n880_));
  MUX2_X1   g679(.A(KEYINPUT121), .B(new_n880_), .S(G127gat), .Z(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n870_), .B2(new_n881_), .ZN(G1342gat));
  NAND3_X1  g681(.A1(new_n860_), .A2(new_n249_), .A3(new_n655_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n564_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n249_), .ZN(G1343gat));
  NOR2_X1   g684(.A1(new_n857_), .A2(new_n675_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n661_), .A2(new_n429_), .A3(new_n451_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n886_), .A2(new_n490_), .A3(new_n887_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT122), .B(G141gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1344gat));
  NAND3_X1  g689(.A1(new_n886_), .A2(new_n644_), .A3(new_n887_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT123), .B(G148gat), .ZN(new_n892_));
  XOR2_X1   g691(.A(new_n891_), .B(new_n892_), .Z(G1345gat));
  NAND3_X1  g692(.A1(new_n886_), .A2(new_n653_), .A3(new_n887_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT61), .B(G155gat), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n894_), .B(new_n895_), .ZN(G1346gat));
  AND4_X1   g695(.A1(G162gat), .A2(new_n886_), .A3(new_n565_), .A4(new_n887_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n887_), .ZN(new_n898_));
  NOR4_X1   g697(.A1(new_n857_), .A2(new_n675_), .A3(new_n654_), .A4(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(G162gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n900_), .A2(KEYINPUT124), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT124), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n899_), .B2(G162gat), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n897_), .B1(new_n902_), .B2(new_n904_), .ZN(G1347gat));
  AND3_X1   g704(.A1(new_n661_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n858_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n490_), .ZN(new_n908_));
  OAI21_X1  g707(.A(G169gat), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n910_), .ZN(new_n912_));
  OAI211_X1 g711(.A(G169gat), .B(new_n912_), .C1(new_n907_), .C2(new_n908_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n907_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n914_), .A2(new_n490_), .A3(new_n236_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n911_), .A2(new_n913_), .A3(new_n915_), .ZN(G1348gat));
  OAI21_X1  g715(.A(G176gat), .B1(new_n907_), .B2(new_n876_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n692_), .A2(new_n232_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n907_), .B2(new_n918_), .ZN(G1349gat));
  NOR3_X1   g718(.A1(new_n907_), .A2(new_n202_), .A3(new_n602_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n914_), .A2(new_n653_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n341_), .B2(new_n921_), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n907_), .B2(new_n564_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n655_), .A2(new_n207_), .A3(new_n345_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n907_), .B2(new_n924_), .ZN(G1351gat));
  NOR2_X1   g724(.A1(new_n662_), .A2(new_n432_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n886_), .A2(new_n490_), .A3(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(KEYINPUT126), .B(G197gat), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n927_), .B2(new_n930_), .ZN(G1352gat));
  NAND3_X1  g730(.A1(new_n886_), .A2(new_n644_), .A3(new_n926_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g732(.A1(new_n886_), .A2(new_n653_), .A3(new_n926_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(KEYINPUT63), .B(G211gat), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n934_), .B2(new_n937_), .ZN(G1354gat));
  NOR2_X1   g737(.A1(new_n654_), .A2(G218gat), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n858_), .A2(new_n267_), .A3(new_n926_), .A4(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(new_n926_), .ZN(new_n941_));
  NOR4_X1   g740(.A1(new_n857_), .A2(new_n675_), .A3(new_n564_), .A4(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(G218gat), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n940_), .B1(new_n942_), .B2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  OAI211_X1 g745(.A(new_n940_), .B(KEYINPUT127), .C1(new_n942_), .C2(new_n943_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(new_n947_), .ZN(G1355gat));
endmodule


