//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n595_, new_n596_, new_n597_, new_n598_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_;
  NAND2_X1  g000(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n202_));
  OR2_X1    g001(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G120gat), .B(G148gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT5), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G176gat), .B(G204gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G99gat), .A3(G106gat), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G85gat), .ZN(new_n213_));
  INV_X1    g012(.A(G92gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(KEYINPUT65), .A3(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(KEYINPUT9), .B1(new_n213_), .B2(new_n214_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n212_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221_));
  INV_X1    g020(.A(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .A4(new_n223_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n215_), .A2(KEYINPUT65), .A3(KEYINPUT9), .A4(new_n216_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n220_), .A2(new_n223_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT64), .B1(new_n226_), .B2(G106gat), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n219_), .A2(new_n224_), .A3(new_n225_), .A4(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G57gat), .B(G64gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n230_));
  XOR2_X1   g029(.A(G71gat), .B(G78gat), .Z(new_n231_));
  OR2_X1    g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n229_), .A2(KEYINPUT11), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n231_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n210_), .B1(G99gat), .B2(G106gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n208_), .A2(KEYINPUT6), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT67), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT7), .ZN(new_n242_));
  INV_X1    g041(.A(G99gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n243_), .A3(new_n222_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n240_), .A2(new_n241_), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n215_), .A2(new_n216_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n236_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n244_), .A2(new_n245_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n212_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n236_), .A2(KEYINPUT66), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n236_), .A2(KEYINPUT66), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n249_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n252_), .A2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n228_), .B(new_n235_), .C1(new_n250_), .C2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G230gat), .ZN(new_n258_));
  INV_X1    g057(.A(G233gat), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n227_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n217_), .A2(new_n218_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n209_), .A2(new_n211_), .A3(KEYINPUT67), .ZN(new_n267_));
  AOI21_X1  g066(.A(KEYINPUT67), .B1(new_n209_), .B2(new_n211_), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n267_), .A2(new_n268_), .A3(new_n251_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT8), .B1(new_n269_), .B2(new_n248_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n256_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n266_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(KEYINPUT12), .B1(new_n272_), .B2(new_n235_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n228_), .B1(new_n250_), .B2(new_n256_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT12), .ZN(new_n275_));
  INV_X1    g074(.A(new_n235_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n262_), .B1(new_n273_), .B2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n276_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n261_), .B1(new_n279_), .B2(new_n257_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n207_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n257_), .A2(new_n261_), .ZN(new_n282_));
  AND3_X1   g081(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n275_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n280_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n207_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n281_), .A2(KEYINPUT68), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT68), .B1(new_n281_), .B2(new_n288_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n202_), .B(new_n203_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT68), .ZN(new_n292_));
  NOR3_X1   g091(.A1(new_n278_), .A2(new_n280_), .A3(new_n207_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n287_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n292_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n281_), .A2(KEYINPUT68), .A3(new_n288_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n295_), .A2(KEYINPUT69), .A3(KEYINPUT13), .A4(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n298_), .A2(new_n299_), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G190gat), .B(G218gat), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT72), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G134gat), .B(G162gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT36), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G29gat), .B(G36gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G43gat), .B(G50gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(new_n228_), .B(new_n314_), .C1(new_n250_), .C2(new_n256_), .ZN(new_n315_));
  XOR2_X1   g114(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n313_), .B(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n315_), .B1(new_n272_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G232gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT34), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT35), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n320_), .B(KEYINPUT35), .Z(new_n323_));
  NAND3_X1  g122(.A1(new_n318_), .A2(KEYINPUT74), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT74), .B1(new_n318_), .B2(new_n323_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n310_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n326_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n309_), .ZN(new_n329_));
  XOR2_X1   g128(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n328_), .A2(new_n322_), .A3(new_n324_), .A4(new_n331_), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n327_), .A2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(KEYINPUT76), .B(KEYINPUT37), .Z(new_n334_));
  XNOR2_X1  g133(.A(new_n310_), .B(KEYINPUT75), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n332_), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n333_), .A2(new_n334_), .B1(new_n337_), .B2(KEYINPUT37), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G231gat), .A2(G233gat), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n234_), .A2(new_n233_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(new_n232_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G1gat), .B(G8gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  XOR2_X1   g144(.A(G15gat), .B(G22gat), .Z(new_n346_));
  NAND2_X1  g145(.A1(G1gat), .A2(G8gat), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n346_), .B1(KEYINPUT14), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n345_), .A2(new_n348_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n340_), .A2(new_n232_), .A3(new_n339_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n342_), .A2(new_n349_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n349_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n351_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n353_), .B1(new_n354_), .B2(new_n341_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT17), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n352_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G127gat), .B(G155gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT16), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G183gat), .B(G211gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT78), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n352_), .A2(new_n355_), .A3(new_n363_), .ZN(new_n364_));
  OR2_X1    g163(.A1(new_n361_), .A2(KEYINPUT17), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n362_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n364_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n338_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n304_), .A2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n371_), .A2(KEYINPUT79), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT23), .ZN(new_n374_));
  OR2_X1    g173(.A1(G169gat), .A2(G176gat), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n375_), .A2(KEYINPUT24), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(KEYINPUT24), .A3(new_n377_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n374_), .A2(new_n376_), .A3(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(KEYINPUT26), .B(G190gat), .Z(new_n380_));
  XOR2_X1   g179(.A(KEYINPUT25), .B(G183gat), .Z(new_n381_));
  OAI21_X1  g180(.A(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n382_), .A2(KEYINPUT92), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n374_), .B1(G183gat), .B2(G190gat), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT93), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n384_), .B(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT83), .B(G176gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT22), .B(G169gat), .ZN(new_n388_));
  AOI22_X1  g187(.A1(new_n387_), .A2(new_n388_), .B1(G169gat), .B2(G176gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n382_), .A2(KEYINPUT92), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n383_), .A2(new_n390_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G197gat), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(G204gat), .ZN(new_n394_));
  INV_X1    g193(.A(G204gat), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n395_), .A2(G197gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT21), .B1(new_n394_), .B2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G211gat), .B(G218gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT88), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n396_), .B1(new_n399_), .B2(new_n394_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n399_), .B2(new_n394_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n397_), .B(new_n398_), .C1(new_n401_), .C2(KEYINPUT21), .ZN(new_n402_));
  INV_X1    g201(.A(new_n398_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(KEYINPUT21), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n392_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G226gat), .A2(G233gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n407_), .B(KEYINPUT19), .Z(new_n408_));
  INV_X1    g207(.A(KEYINPUT20), .ZN(new_n409_));
  NOR2_X1   g208(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT82), .B(G183gat), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n410_), .B1(new_n411_), .B2(KEYINPUT25), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n379_), .B1(new_n380_), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n374_), .B1(G190gat), .B2(new_n411_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n389_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n409_), .B1(new_n416_), .B2(new_n405_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n406_), .A2(new_n408_), .A3(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n392_), .A2(new_n405_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n416_), .A2(new_n405_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n420_), .A2(new_n409_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n408_), .B(KEYINPUT91), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT18), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G64gat), .B(G92gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n426_), .B(new_n427_), .Z(new_n428_));
  NAND3_X1  g227(.A1(new_n418_), .A2(new_n424_), .A3(new_n428_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n402_), .A2(new_n404_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n390_), .A2(new_n430_), .A3(new_n382_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n408_), .B1(new_n431_), .B2(new_n417_), .ZN(new_n432_));
  OR2_X1    g231(.A1(new_n432_), .A2(KEYINPUT97), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(KEYINPUT97), .ZN(new_n434_));
  INV_X1    g233(.A(new_n423_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n419_), .A2(new_n435_), .A3(new_n421_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n428_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(KEYINPUT98), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT98), .B1(new_n437_), .B2(new_n438_), .ZN(new_n441_));
  OAI211_X1 g240(.A(KEYINPUT27), .B(new_n429_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n418_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n424_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n438_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n445_), .A2(KEYINPUT94), .A3(new_n429_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT27), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT94), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n448_), .B(new_n438_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n446_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n442_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI211_X1 g251(.A(G228gat), .B(G233gat), .C1(new_n430_), .C2(KEYINPUT89), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(G106gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(G141gat), .A2(G148gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT86), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G141gat), .A2(G148gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G155gat), .B(G162gat), .Z(new_n460_));
  INV_X1    g259(.A(KEYINPUT1), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT3), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n455_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT2), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n457_), .A2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n464_), .A2(new_n466_), .A3(new_n467_), .A4(new_n468_), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n459_), .A2(new_n462_), .B1(new_n460_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT29), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n405_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(G78gat), .ZN(new_n473_));
  XOR2_X1   g272(.A(new_n454_), .B(new_n473_), .Z(new_n474_));
  NAND2_X1  g273(.A1(new_n470_), .A2(new_n471_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G22gat), .B(G50gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT90), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n480_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n474_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n454_), .B(new_n473_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(new_n480_), .A3(new_n479_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G227gat), .A2(G233gat), .ZN(new_n487_));
  INV_X1    g286(.A(G15gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT30), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n416_), .B(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G127gat), .B(G134gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G113gat), .B(G120gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT84), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT85), .B1(new_n492_), .B2(new_n493_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n492_), .A2(new_n493_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT85), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n496_), .A2(new_n497_), .A3(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n491_), .B(new_n501_), .Z(new_n502_));
  XNOR2_X1  g301(.A(G71gat), .B(G99gat), .ZN(new_n503_));
  INV_X1    g302(.A(G43gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(KEYINPUT31), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n502_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n502_), .A2(new_n506_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G1gat), .B(G29gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(G85gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT0), .B(G57gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n512_), .B(new_n513_), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT4), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n501_), .A2(new_n470_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n494_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n470_), .B1(new_n518_), .B2(new_n498_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n516_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n520_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G225gat), .A2(G233gat), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n517_), .A2(new_n519_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(new_n522_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n515_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n524_), .A2(new_n515_), .A3(new_n526_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n510_), .A2(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n452_), .A2(KEYINPUT99), .A3(new_n486_), .A4(new_n531_), .ZN(new_n532_));
  NAND4_X1  g331(.A1(new_n531_), .A2(new_n486_), .A3(new_n442_), .A4(new_n450_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT99), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n446_), .A2(new_n449_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT95), .ZN(new_n537_));
  OR3_X1    g336(.A1(new_n527_), .A2(new_n537_), .A3(KEYINPUT33), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n517_), .A2(new_n519_), .A3(new_n523_), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n515_), .B(new_n539_), .C1(new_n521_), .C2(new_n523_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT33), .B1(new_n527_), .B2(new_n537_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n536_), .A2(new_n538_), .A3(new_n540_), .A4(new_n541_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n443_), .A2(new_n444_), .A3(KEYINPUT96), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n428_), .A2(KEYINPUT32), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n433_), .A2(new_n434_), .A3(new_n436_), .A4(new_n545_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n418_), .A2(new_n424_), .A3(KEYINPUT96), .ZN(new_n547_));
  OAI22_X1  g346(.A1(new_n543_), .A2(new_n546_), .B1(new_n545_), .B2(new_n547_), .ZN(new_n548_));
  AOI22_X1  g347(.A1(new_n548_), .A2(new_n530_), .B1(new_n483_), .B2(new_n485_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n509_), .B1(new_n542_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n486_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n451_), .B2(new_n530_), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n532_), .A2(new_n535_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  XOR2_X1   g352(.A(G113gat), .B(G141gat), .Z(new_n554_));
  XOR2_X1   g353(.A(G169gat), .B(G197gat), .Z(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  XOR2_X1   g355(.A(new_n556_), .B(KEYINPUT80), .Z(new_n557_));
  NAND2_X1  g356(.A1(new_n317_), .A2(new_n353_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n350_), .A2(new_n349_), .A3(new_n313_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n353_), .A2(new_n314_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n560_), .B1(new_n562_), .B2(new_n559_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n557_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT81), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n561_), .A2(new_n563_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(new_n556_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT81), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n568_), .B(new_n557_), .C1(new_n561_), .C2(new_n563_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n565_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n553_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n371_), .A2(KEYINPUT79), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n372_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n530_), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n574_), .A2(G1gat), .A3(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n577_));
  OR2_X1    g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n577_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n553_), .A2(new_n369_), .A3(new_n333_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n303_), .A2(new_n571_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(G1gat), .B1(new_n583_), .B2(new_n575_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n578_), .A2(new_n579_), .A3(new_n584_), .ZN(G1324gat));
  INV_X1    g384(.A(KEYINPUT39), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n451_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n586_), .B1(new_n587_), .B2(G8gat), .ZN(new_n588_));
  INV_X1    g387(.A(G8gat), .ZN(new_n589_));
  AOI211_X1 g388(.A(KEYINPUT39), .B(new_n589_), .C1(new_n582_), .C2(new_n451_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n451_), .A2(new_n589_), .ZN(new_n591_));
  OAI22_X1  g390(.A1(new_n588_), .A2(new_n590_), .B1(new_n574_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT40), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(G1325gat));
  AOI21_X1  g393(.A(new_n488_), .B1(new_n582_), .B2(new_n509_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(KEYINPUT41), .ZN(new_n596_));
  INV_X1    g395(.A(new_n574_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(new_n488_), .A3(new_n509_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(G1326gat));
  INV_X1    g398(.A(G22gat), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n582_), .B2(new_n551_), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT42), .Z(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(new_n600_), .A3(new_n551_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(G1327gat));
  INV_X1    g403(.A(new_n333_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n303_), .A2(new_n368_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n572_), .A2(new_n606_), .ZN(new_n607_));
  OR3_X1    g406(.A1(new_n607_), .A2(G29gat), .A3(new_n575_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n532_), .A2(new_n535_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n550_), .A2(new_n552_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(KEYINPUT101), .A2(KEYINPUT43), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n611_), .A2(new_n338_), .A3(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n338_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n612_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(KEYINPUT101), .A2(KEYINPUT43), .ZN(new_n616_));
  OAI22_X1  g415(.A1(new_n553_), .A2(new_n614_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n613_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n581_), .A2(new_n369_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(KEYINPUT44), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT44), .ZN(new_n622_));
  AOI211_X1 g421(.A(new_n622_), .B(new_n619_), .C1(new_n613_), .C2(new_n617_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n621_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(KEYINPUT102), .A3(new_n530_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G29gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT102), .B1(new_n624_), .B2(new_n530_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n608_), .B1(new_n626_), .B2(new_n627_), .ZN(G1328gat));
  XNOR2_X1  g427(.A(KEYINPUT104), .B(KEYINPUT46), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n452_), .A2(G36gat), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n572_), .A2(new_n606_), .A3(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT45), .Z(new_n633_));
  NAND2_X1  g432(.A1(new_n618_), .A2(new_n620_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n622_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n618_), .A2(KEYINPUT44), .A3(new_n620_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n635_), .A2(new_n451_), .A3(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n633_), .B1(new_n637_), .B2(G36gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n630_), .B1(new_n638_), .B2(KEYINPUT103), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT103), .ZN(new_n640_));
  INV_X1    g439(.A(G36gat), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n641_), .B1(new_n624_), .B2(new_n451_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n640_), .B(new_n629_), .C1(new_n642_), .C2(new_n633_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n639_), .A2(new_n643_), .ZN(G1329gat));
  NAND3_X1  g443(.A1(new_n624_), .A2(G43gat), .A3(new_n509_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n504_), .B1(new_n607_), .B2(new_n510_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n645_), .A2(KEYINPUT47), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT47), .B1(new_n645_), .B2(new_n646_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1330gat));
  INV_X1    g448(.A(new_n607_), .ZN(new_n650_));
  AOI21_X1  g449(.A(G50gat), .B1(new_n650_), .B2(new_n551_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n551_), .A2(G50gat), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n651_), .B1(new_n624_), .B2(new_n653_), .ZN(G1331gat));
  NOR2_X1   g453(.A1(new_n304_), .A2(new_n570_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n580_), .A2(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G57gat), .B1(new_n656_), .B2(new_n575_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n553_), .A2(new_n304_), .A3(new_n570_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n370_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n575_), .A2(G57gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n657_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT105), .ZN(G1332gat));
  OR3_X1    g461(.A1(new_n659_), .A2(G64gat), .A3(new_n452_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G64gat), .B1(new_n656_), .B2(new_n452_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n664_), .A2(KEYINPUT48), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(KEYINPUT48), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n663_), .B1(new_n665_), .B2(new_n666_), .ZN(G1333gat));
  OR3_X1    g466(.A1(new_n659_), .A2(G71gat), .A3(new_n510_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G71gat), .B1(new_n656_), .B2(new_n510_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(KEYINPUT49), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(KEYINPUT49), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n668_), .B1(new_n670_), .B2(new_n671_), .ZN(G1334gat));
  OAI21_X1  g471(.A(G78gat), .B1(new_n656_), .B2(new_n486_), .ZN(new_n673_));
  XOR2_X1   g472(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n673_), .A2(new_n675_), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n486_), .A2(G78gat), .ZN(new_n678_));
  OAI22_X1  g477(.A1(new_n676_), .A2(new_n677_), .B1(new_n659_), .B2(new_n678_), .ZN(G1335gat));
  NAND2_X1  g478(.A1(new_n655_), .A2(new_n369_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n613_), .B2(new_n617_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G85gat), .B1(new_n682_), .B2(new_n575_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n605_), .A2(new_n368_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n658_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n686_), .A2(new_n213_), .A3(new_n530_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n683_), .A2(new_n687_), .ZN(G1336gat));
  OAI21_X1  g487(.A(G92gat), .B1(new_n682_), .B2(new_n452_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n686_), .A2(new_n214_), .A3(new_n451_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1337gat));
  OR3_X1    g490(.A1(new_n685_), .A2(new_n226_), .A3(new_n510_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT107), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n243_), .B1(new_n681_), .B2(new_n509_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT51), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n692_), .B(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT51), .ZN(new_n698_));
  INV_X1    g497(.A(new_n694_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n695_), .A2(new_n700_), .ZN(G1338gat));
  INV_X1    g500(.A(KEYINPUT52), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n681_), .A2(new_n551_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(G106gat), .ZN(new_n704_));
  AOI211_X1 g503(.A(KEYINPUT52), .B(new_n222_), .C1(new_n681_), .C2(new_n551_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n551_), .A2(new_n222_), .ZN(new_n706_));
  OAI22_X1  g505(.A1(new_n704_), .A2(new_n705_), .B1(new_n685_), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g507(.A(KEYINPUT117), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n570_), .A2(new_n366_), .A3(new_n367_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n291_), .A2(new_n297_), .A3(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n338_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n291_), .A2(new_n297_), .A3(new_n710_), .A4(KEYINPUT108), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n713_), .A2(new_n714_), .A3(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n715_), .B(KEYINPUT110), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n718_), .A2(new_n721_), .A3(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n711_), .A2(new_n712_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n724_), .A2(new_n614_), .A3(new_n714_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n719_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n713_), .A2(new_n714_), .A3(new_n717_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT111), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n723_), .A2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(KEYINPUT55), .B(new_n282_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n273_), .A2(new_n277_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n733_), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(new_n282_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT55), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n285_), .A2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n257_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n260_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n732_), .A2(new_n734_), .A3(new_n736_), .A4(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(KEYINPUT56), .A3(new_n207_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n207_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT56), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n739_), .A2(KEYINPUT115), .A3(KEYINPUT56), .A4(new_n207_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n558_), .A2(G229gat), .A3(G233gat), .A4(new_n559_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n562_), .A2(new_n559_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n556_), .B1(new_n749_), .B2(new_n560_), .ZN(new_n750_));
  AOI22_X1  g549(.A1(new_n566_), .A2(new_n556_), .B1(new_n748_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n288_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT58), .B1(new_n747_), .B2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT116), .B1(new_n754_), .B2(new_n614_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT116), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT56), .B1(new_n739_), .B2(new_n207_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n741_), .B2(new_n740_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n752_), .B1(new_n758_), .B2(new_n746_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n756_), .B(new_n338_), .C1(new_n759_), .C2(KEYINPUT58), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n747_), .A2(KEYINPUT58), .A3(new_n753_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n755_), .A2(new_n760_), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT113), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT114), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT57), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n764_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n570_), .A2(new_n288_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n739_), .A2(KEYINPUT56), .A3(new_n207_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(new_n757_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n751_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n767_), .B1(new_n772_), .B2(new_n333_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n333_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n765_), .B1(new_n774_), .B2(new_n764_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n773_), .B1(new_n775_), .B2(KEYINPUT57), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n368_), .B1(new_n763_), .B2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n709_), .B1(new_n729_), .B2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n722_), .B1(new_n718_), .B2(new_n721_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n726_), .A2(KEYINPUT111), .A3(new_n727_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n754_), .A2(new_n614_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n761_), .B1(new_n782_), .B2(new_n756_), .ZN(new_n783_));
  AOI211_X1 g582(.A(KEYINPUT113), .B(new_n333_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n766_), .B1(new_n784_), .B2(new_n765_), .ZN(new_n785_));
  AOI22_X1  g584(.A1(new_n783_), .A2(new_n755_), .B1(new_n785_), .B2(new_n773_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n781_), .B(KEYINPUT117), .C1(new_n786_), .C2(new_n368_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n778_), .A2(new_n787_), .ZN(new_n788_));
  NOR4_X1   g587(.A1(new_n451_), .A2(new_n551_), .A3(new_n575_), .A4(new_n510_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT59), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n729_), .A2(new_n777_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n789_), .B1(KEYINPUT118), .B2(KEYINPUT59), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n793_), .B1(KEYINPUT118), .B2(new_n789_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n791_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(G113gat), .B1(new_n795_), .B2(new_n571_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n571_), .A2(G113gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n790_), .B2(new_n797_), .ZN(G1340gat));
  OAI21_X1  g597(.A(G120gat), .B1(new_n795_), .B2(new_n304_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n304_), .A2(KEYINPUT60), .ZN(new_n800_));
  MUX2_X1   g599(.A(new_n800_), .B(KEYINPUT60), .S(G120gat), .Z(new_n801_));
  NAND3_X1  g600(.A1(new_n788_), .A2(new_n789_), .A3(new_n801_), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n802_), .B(KEYINPUT119), .Z(new_n803_));
  NAND2_X1  g602(.A1(new_n799_), .A2(new_n803_), .ZN(G1341gat));
  OAI21_X1  g603(.A(G127gat), .B1(new_n795_), .B2(new_n369_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n369_), .A2(G127gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n790_), .B2(new_n806_), .ZN(G1342gat));
  OAI21_X1  g606(.A(G134gat), .B1(new_n795_), .B2(new_n614_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n605_), .A2(G134gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n808_), .B1(new_n790_), .B2(new_n809_), .ZN(G1343gat));
  NOR2_X1   g609(.A1(new_n486_), .A2(new_n509_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n812_), .A2(new_n451_), .A3(new_n575_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n778_), .B2(new_n787_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n570_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n303_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g618(.A1(new_n815_), .A2(new_n368_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT61), .B(G155gat), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n820_), .B(new_n821_), .ZN(G1346gat));
  NAND3_X1  g621(.A1(new_n815_), .A2(G162gat), .A3(new_n338_), .ZN(new_n823_));
  AOI211_X1 g622(.A(KEYINPUT120), .B(G162gat), .C1(new_n815_), .C2(new_n333_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n729_), .A2(new_n777_), .A3(new_n709_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n763_), .A2(new_n776_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n369_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT117), .B1(new_n828_), .B2(new_n781_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n333_), .B(new_n813_), .C1(new_n826_), .C2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(G162gat), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n825_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n823_), .B1(new_n824_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT121), .B(new_n823_), .C1(new_n824_), .C2(new_n832_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(G1347gat));
  AND2_X1   g636(.A1(new_n451_), .A2(new_n531_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n486_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n792_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(G169gat), .B1(new_n841_), .B2(new_n571_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT62), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n570_), .A2(new_n388_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n844_), .B(KEYINPUT122), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n843_), .B1(new_n841_), .B2(new_n845_), .ZN(G1348gat));
  NAND2_X1  g645(.A1(new_n788_), .A2(new_n486_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n788_), .A2(KEYINPUT123), .A3(new_n486_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n849_), .A2(new_n838_), .A3(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n303_), .A2(G176gat), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n840_), .A2(new_n303_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n851_), .A2(new_n852_), .B1(new_n387_), .B2(new_n853_), .ZN(G1349gat));
  AND3_X1   g653(.A1(new_n840_), .A2(new_n368_), .A3(new_n381_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n851_), .A2(new_n368_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n411_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(G1350gat));
  OR3_X1    g657(.A1(new_n841_), .A2(new_n605_), .A3(new_n380_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n840_), .A2(new_n338_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n860_), .A2(KEYINPUT124), .A3(G190gat), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT124), .B1(new_n860_), .B2(G190gat), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n859_), .B1(new_n861_), .B2(new_n862_), .ZN(G1351gat));
  NOR3_X1   g662(.A1(new_n812_), .A2(new_n452_), .A3(new_n530_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n788_), .A2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n571_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(new_n393_), .ZN(G1352gat));
  NOR2_X1   g666(.A1(new_n865_), .A2(new_n304_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n395_), .A2(KEYINPUT125), .ZN(new_n869_));
  AND2_X1   g668(.A1(new_n395_), .A2(KEYINPUT125), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n868_), .B2(new_n870_), .ZN(G1353gat));
  NOR2_X1   g671(.A1(new_n865_), .A2(new_n369_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n873_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n874_));
  XOR2_X1   g673(.A(KEYINPUT63), .B(G211gat), .Z(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n873_), .B2(new_n875_), .ZN(G1354gat));
  XNOR2_X1  g675(.A(KEYINPUT127), .B(G218gat), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n865_), .A2(new_n614_), .A3(new_n877_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n788_), .A2(new_n333_), .A3(new_n864_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT126), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n878_), .B1(new_n880_), .B2(new_n877_), .ZN(G1355gat));
endmodule


