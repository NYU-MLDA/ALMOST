//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n942_, new_n943_, new_n944_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT28), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(KEYINPUT88), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208_));
  AND3_X1   g007(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT89), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND4_X1  g013(.A1(KEYINPUT89), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G141gat), .ZN(new_n217_));
  INV_X1    g016(.A(G148gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(new_n218_), .A3(KEYINPUT3), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n211_), .A2(new_n216_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT90), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n211_), .A2(new_n216_), .A3(KEYINPUT90), .A4(new_n222_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n207_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G141gat), .A2(G148gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT87), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(KEYINPUT87), .A2(G141gat), .A3(G148gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n232_), .B1(G141gat), .B2(G148gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n206_), .B(KEYINPUT1), .Z(new_n234_));
  AOI21_X1  g033(.A(new_n233_), .B1(new_n205_), .B2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n227_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n203_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NOR4_X1   g038(.A1(new_n227_), .A2(KEYINPUT28), .A3(KEYINPUT29), .A4(new_n235_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G22gat), .B(G50gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n242_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT91), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G78gat), .B(G106gat), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT21), .ZN(new_n250_));
  INV_X1    g049(.A(G197gat), .ZN(new_n251_));
  INV_X1    g050(.A(G204gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT92), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT92), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G204gat), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n251_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(G197gat), .A2(G204gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n250_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(G218gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(G211gat), .ZN(new_n260_));
  INV_X1    g059(.A(G211gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(G218gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n253_), .A2(new_n255_), .A3(new_n251_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n250_), .B1(G197gat), .B2(G204gat), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n258_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT93), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n256_), .A2(new_n257_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n250_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n267_), .A2(new_n268_), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n268_), .B1(new_n267_), .B2(new_n271_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT29), .B1(new_n227_), .B2(new_n235_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G228gat), .A2(G233gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n267_), .A2(new_n271_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n276_), .B1(new_n275_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n249_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n275_), .A2(new_n279_), .ZN(new_n282_));
  OAI211_X1 g081(.A(new_n277_), .B(new_n248_), .C1(new_n282_), .C2(new_n276_), .ZN(new_n283_));
  NAND4_X1  g082(.A1(new_n246_), .A2(new_n247_), .A3(new_n281_), .A4(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(new_n283_), .A3(new_n247_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n244_), .A2(new_n245_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n284_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G226gat), .A2(G233gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT19), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT24), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(G169gat), .ZN(new_n299_));
  INV_X1    g098(.A(G176gat), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n301_), .A2(new_n295_), .A3(new_n294_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT25), .B(G183gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(KEYINPUT26), .B(G190gat), .ZN(new_n304_));
  AOI211_X1 g103(.A(new_n298_), .B(new_n302_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n297_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n306_), .A2(new_n292_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n307_), .B1(G183gat), .B2(G190gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT96), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT22), .B(G169gat), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n301_), .B1(new_n310_), .B2(new_n300_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT95), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n305_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n279_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT20), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n279_), .A2(KEYINPUT93), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n267_), .A2(new_n268_), .A3(new_n271_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT83), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n298_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(G190gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT81), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT81), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(G190gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n325_), .A3(KEYINPUT26), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT82), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT81), .B(G190gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT82), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(KEYINPUT26), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n322_), .A2(KEYINPUT26), .ZN(new_n332_));
  AND2_X1   g131(.A1(new_n303_), .A2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n302_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n301_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT84), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n299_), .A2(KEYINPUT22), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT22), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(G169gat), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n336_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n336_), .B1(new_n338_), .B2(G169gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(new_n300_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n335_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(G183gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n328_), .A2(new_n344_), .ZN(new_n345_));
  AOI22_X1  g144(.A1(new_n343_), .A2(KEYINPUT85), .B1(new_n307_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT85), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n347_), .B(new_n335_), .C1(new_n340_), .C2(new_n342_), .ZN(new_n348_));
  AOI22_X1  g147(.A1(new_n321_), .A2(new_n334_), .B1(new_n346_), .B2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n316_), .B1(new_n319_), .B2(new_n349_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n315_), .B1(new_n350_), .B2(KEYINPUT94), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n334_), .A2(new_n321_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n346_), .A2(new_n348_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n352_), .B(new_n353_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT94), .B1(new_n354_), .B2(KEYINPUT20), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n291_), .B1(new_n351_), .B2(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G8gat), .B(G36gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT18), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G64gat), .B(G92gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n359_), .B(new_n360_), .Z(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n316_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n352_), .A2(new_n353_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n274_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n365_), .A3(new_n291_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR3_X1   g166(.A1(new_n357_), .A2(new_n362_), .A3(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n361_), .B(KEYINPUT98), .Z(new_n369_));
  NAND3_X1  g168(.A1(new_n351_), .A2(new_n356_), .A3(new_n291_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n291_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT27), .ZN(new_n374_));
  NOR3_X1   g173(.A1(new_n368_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n362_), .B1(new_n357_), .B2(new_n367_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n354_), .A2(KEYINPUT94), .A3(KEYINPUT20), .ZN(new_n377_));
  OR2_X1    g176(.A1(new_n313_), .A2(new_n314_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n290_), .B1(new_n379_), .B2(new_n355_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(new_n361_), .A3(new_n366_), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT27), .B1(new_n376_), .B2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT99), .B1(new_n375_), .B2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n361_), .B1(new_n380_), .B2(new_n366_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n374_), .B1(new_n368_), .B2(new_n384_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n379_), .A2(new_n290_), .A3(new_n355_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n386_), .A2(new_n371_), .ZN(new_n387_));
  OAI211_X1 g186(.A(KEYINPUT27), .B(new_n381_), .C1(new_n387_), .C2(new_n369_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT99), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n288_), .B1(new_n383_), .B2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G71gat), .B(G99gat), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n392_), .B(G43gat), .Z(new_n393_));
  XNOR2_X1  g192(.A(new_n349_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G113gat), .B(G120gat), .ZN(new_n395_));
  XOR2_X1   g194(.A(G127gat), .B(G134gat), .Z(new_n396_));
  INV_X1    g195(.A(KEYINPUT86), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G127gat), .B(G134gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT86), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n395_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n398_), .A2(new_n400_), .A3(new_n395_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n394_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G227gat), .A2(G233gat), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n406_), .B(G15gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT30), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT31), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n394_), .A2(new_n404_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n405_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n409_), .B1(new_n405_), .B2(new_n410_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n207_), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n232_), .A2(new_n208_), .B1(new_n221_), .B2(new_n219_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT90), .B1(new_n415_), .B2(new_n216_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n226_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n414_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n235_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n404_), .A3(new_n419_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n398_), .A2(new_n400_), .A3(new_n395_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n421_), .A2(new_n401_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n422_), .B1(new_n227_), .B2(new_n235_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G225gat), .A2(G233gat), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n420_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G1gat), .B(G29gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(G85gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT0), .B(G57gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n427_), .B(new_n428_), .Z(new_n429_));
  AND3_X1   g228(.A1(new_n420_), .A2(new_n423_), .A3(KEYINPUT4), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n422_), .B(new_n431_), .C1(new_n227_), .C2(new_n235_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n424_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  OAI211_X1 g233(.A(new_n425_), .B(new_n429_), .C1(new_n430_), .C2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT97), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n425_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n429_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n420_), .A2(new_n423_), .A3(KEYINPUT4), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(new_n433_), .A3(new_n432_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT97), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n441_), .A2(new_n442_), .A3(new_n425_), .A4(new_n429_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n436_), .A2(new_n439_), .A3(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n413_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT33), .ZN(new_n446_));
  OR2_X1    g245(.A1(new_n435_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n440_), .A2(new_n424_), .A3(new_n432_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n420_), .A2(new_n423_), .A3(new_n433_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n449_), .A2(new_n438_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n435_), .A2(new_n446_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n376_), .A2(new_n381_), .A3(new_n447_), .A4(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n361_), .A2(KEYINPUT32), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n454_), .B1(new_n386_), .B2(new_n371_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n380_), .A2(new_n453_), .A3(new_n366_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n444_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n452_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n288_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n444_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n385_), .A3(new_n388_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n391_), .A2(new_n445_), .B1(new_n463_), .B2(new_n413_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G190gat), .B(G218gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G134gat), .B(G162gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT36), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT70), .ZN(new_n469_));
  OR2_X1    g268(.A1(G85gat), .A2(G92gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G85gat), .A2(G92gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT67), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT67), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(new_n474_), .A3(new_n471_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(G99gat), .A2(G106gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT7), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT6), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(G99gat), .A3(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n476_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n483_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT65), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT65), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n483_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n489_), .A3(new_n478_), .ZN(new_n490_));
  XOR2_X1   g289(.A(KEYINPUT66), .B(KEYINPUT8), .Z(new_n491_));
  AND3_X1   g290(.A1(new_n473_), .A2(new_n475_), .A3(new_n491_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n485_), .A2(KEYINPUT8), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n487_), .A2(new_n489_), .ZN(new_n494_));
  OR2_X1    g293(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT64), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n495_), .A2(KEYINPUT64), .A3(new_n496_), .ZN(new_n500_));
  AOI21_X1  g299(.A(G106gat), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n470_), .A2(KEYINPUT9), .A3(new_n471_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n502_), .B1(KEYINPUT9), .B2(new_n471_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n494_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n469_), .B1(new_n493_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n494_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n501_), .A2(new_n503_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n490_), .A2(new_n492_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT8), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n510_), .B1(new_n476_), .B2(new_n484_), .ZN(new_n511_));
  OAI211_X1 g310(.A(KEYINPUT70), .B(new_n508_), .C1(new_n509_), .C2(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G29gat), .B(G36gat), .Z(new_n513_));
  XOR2_X1   g312(.A(G43gat), .B(G50gat), .Z(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT15), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n505_), .A2(new_n512_), .A3(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G232gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(KEYINPUT74), .A3(KEYINPUT35), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n521_), .B1(KEYINPUT35), .B2(new_n520_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n485_), .A2(KEYINPUT8), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n490_), .A2(new_n492_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n504_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n522_), .B1(new_n525_), .B2(new_n515_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n520_), .A2(KEYINPUT35), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT74), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n517_), .A2(new_n526_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n529_), .B1(new_n517_), .B2(new_n526_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n467_), .A2(KEYINPUT36), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n531_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n533_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n517_), .A2(new_n526_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n529_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n535_), .B1(new_n538_), .B2(new_n530_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n468_), .B1(new_n534_), .B2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n464_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT71), .ZN(new_n542_));
  XOR2_X1   g341(.A(G71gat), .B(G78gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(G57gat), .B(G64gat), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n543_), .B1(KEYINPUT11), .B2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT68), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(KEYINPUT11), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n508_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n548_), .A2(new_n549_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT12), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n550_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n548_), .A2(new_n505_), .A3(KEYINPUT12), .A4(new_n512_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT69), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n548_), .A2(new_n557_), .A3(new_n549_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n555_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n550_), .A2(KEYINPUT69), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n558_), .B(new_n559_), .C1(new_n560_), .C2(new_n551_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G120gat), .B(G148gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT5), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G176gat), .B(G204gat), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n563_), .B(new_n564_), .Z(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n556_), .A2(new_n561_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n566_), .B1(new_n556_), .B2(new_n561_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n542_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n569_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(KEYINPUT71), .A3(new_n567_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT72), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n574_), .A2(KEYINPUT13), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(KEYINPUT13), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n573_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT13), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n570_), .A2(new_n572_), .A3(KEYINPUT72), .A4(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(KEYINPUT77), .B(G8gat), .Z(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT14), .B1(new_n582_), .B2(new_n202_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G15gat), .B(G22gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G1gat), .B(G8gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n515_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n586_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n585_), .B(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n515_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G229gat), .A2(G233gat), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n516_), .A2(new_n587_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n595_), .B1(new_n591_), .B2(new_n515_), .ZN(new_n597_));
  AOI22_X1  g396(.A1(new_n593_), .A2(new_n595_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G113gat), .B(G141gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G169gat), .B(G197gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT80), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(KEYINPUT80), .B1(new_n598_), .B2(new_n601_), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n598_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n601_), .B1(new_n607_), .B2(KEYINPUT79), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(KEYINPUT79), .B2(new_n607_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n548_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(new_n591_), .ZN(new_n614_));
  XOR2_X1   g413(.A(G127gat), .B(G155gat), .Z(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT17), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n614_), .A2(new_n621_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n620_), .A2(KEYINPUT17), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n614_), .A2(new_n621_), .A3(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n581_), .A2(new_n611_), .A3(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n541_), .A2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n202_), .B1(new_n627_), .B2(new_n444_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n385_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n389_), .B1(new_n385_), .B2(new_n388_), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n459_), .B(new_n445_), .C1(new_n629_), .C2(new_n630_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n461_), .A2(new_n385_), .A3(new_n388_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n288_), .B1(new_n452_), .B2(new_n457_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n413_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n610_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT100), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT37), .B1(new_n539_), .B2(KEYINPUT75), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT76), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n533_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n538_), .A2(new_n535_), .A3(new_n530_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n639_), .B1(new_n642_), .B2(new_n468_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n468_), .ZN(new_n644_));
  AOI211_X1 g443(.A(KEYINPUT76), .B(new_n644_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n638_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n540_), .A2(KEYINPUT76), .ZN(new_n647_));
  INV_X1    g446(.A(new_n638_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n642_), .A2(new_n639_), .A3(new_n468_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n646_), .A2(new_n650_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n581_), .A2(new_n651_), .A3(new_n625_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n637_), .A2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n444_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n653_), .A2(G1gat), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n628_), .B1(new_n655_), .B2(KEYINPUT38), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n655_), .A2(KEYINPUT38), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n657_), .A2(KEYINPUT101), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(KEYINPUT101), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n656_), .B1(new_n658_), .B2(new_n659_), .ZN(G1324gat));
  INV_X1    g459(.A(G8gat), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n629_), .A2(new_n630_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n627_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n637_), .A2(new_n662_), .A3(new_n582_), .A4(new_n652_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(G1325gat));
  INV_X1    g468(.A(new_n413_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n627_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G15gat), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT41), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n653_), .A2(G15gat), .A3(new_n413_), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1326gat));
  INV_X1    g474(.A(G22gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n627_), .B2(new_n288_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT42), .Z(new_n678_));
  NAND2_X1  g477(.A1(new_n288_), .A2(new_n676_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT103), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n678_), .B1(new_n653_), .B2(new_n680_), .ZN(G1327gat));
  NAND2_X1  g480(.A1(new_n625_), .A2(new_n540_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT106), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n578_), .A2(new_n580_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n637_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G29gat), .B1(new_n687_), .B2(new_n444_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n684_), .A2(new_n610_), .A3(new_n625_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n646_), .A2(new_n650_), .A3(KEYINPUT104), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n690_), .A2(KEYINPUT43), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n646_), .A2(new_n650_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n464_), .B2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(KEYINPUT43), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n635_), .A2(new_n651_), .A3(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n689_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n696_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n698_));
  INV_X1    g497(.A(new_n625_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n581_), .A2(new_n611_), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701_));
  AOI221_X4 g500(.A(new_n692_), .B1(new_n701_), .B2(KEYINPUT43), .C1(new_n631_), .C2(new_n634_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n694_), .B1(new_n635_), .B2(new_n651_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n700_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n698_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n697_), .A2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(KEYINPUT44), .B(new_n700_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n444_), .A2(G29gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n688_), .B1(new_n710_), .B2(new_n711_), .ZN(G1328gat));
  INV_X1    g511(.A(new_n662_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n713_), .A2(G36gat), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  OR3_X1    g514(.A1(new_n686_), .A2(KEYINPUT45), .A3(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT45), .B1(new_n686_), .B2(new_n715_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n708_), .A2(new_n662_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n720_), .B1(new_n697_), .B2(new_n706_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT107), .B1(new_n721_), .B2(G36gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT105), .B1(new_n696_), .B2(KEYINPUT44), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n704_), .A2(new_n698_), .A3(new_n705_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n719_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n726_));
  INV_X1    g525(.A(G36gat), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n718_), .B1(new_n722_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT46), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  OAI211_X1 g530(.A(KEYINPUT46), .B(new_n718_), .C1(new_n722_), .C2(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1329gat));
  XNOR2_X1  g532(.A(KEYINPUT108), .B(G43gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n687_), .B2(new_n670_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n670_), .A2(G43gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n710_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT47), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(G1330gat));
  NOR3_X1   g538(.A1(new_n707_), .A2(new_n459_), .A3(new_n709_), .ZN(new_n740_));
  INV_X1    g539(.A(G50gat), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n288_), .A2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT109), .ZN(new_n743_));
  OAI22_X1  g542(.A1(new_n740_), .A2(new_n741_), .B1(new_n686_), .B2(new_n743_), .ZN(G1331gat));
  NAND2_X1  g543(.A1(new_n581_), .A2(new_n611_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n745_), .A2(new_n625_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n541_), .ZN(new_n747_));
  INV_X1    g546(.A(G57gat), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n654_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n684_), .A2(new_n651_), .A3(new_n625_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n464_), .A2(new_n610_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n752_), .B2(new_n654_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n754_), .A2(KEYINPUT110), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(KEYINPUT110), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n749_), .B1(new_n755_), .B2(new_n756_), .ZN(G1332gat));
  OR3_X1    g556(.A1(new_n752_), .A2(G64gat), .A3(new_n713_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G64gat), .B1(new_n747_), .B2(new_n713_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(KEYINPUT48), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(KEYINPUT48), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n758_), .B1(new_n760_), .B2(new_n761_), .ZN(G1333gat));
  OR3_X1    g561(.A1(new_n752_), .A2(G71gat), .A3(new_n413_), .ZN(new_n763_));
  OAI21_X1  g562(.A(G71gat), .B1(new_n747_), .B2(new_n413_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n764_), .A2(KEYINPUT49), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n764_), .A2(KEYINPUT49), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n763_), .B1(new_n765_), .B2(new_n766_), .ZN(G1334gat));
  OR3_X1    g566(.A1(new_n752_), .A2(G78gat), .A3(new_n459_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G78gat), .B1(new_n747_), .B2(new_n459_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n769_), .A2(KEYINPUT50), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(KEYINPUT50), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n768_), .B1(new_n770_), .B2(new_n771_), .ZN(G1335gat));
  NAND2_X1  g571(.A1(new_n693_), .A2(new_n695_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n745_), .A2(new_n699_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G85gat), .B1(new_n775_), .B2(new_n654_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n751_), .A2(new_n581_), .A3(new_n683_), .ZN(new_n777_));
  INV_X1    g576(.A(G85gat), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n777_), .A2(new_n778_), .A3(new_n444_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(G1336gat));
  AOI21_X1  g579(.A(G92gat), .B1(new_n777_), .B2(new_n662_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n775_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n662_), .A2(G92gat), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT111), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n781_), .B1(new_n782_), .B2(new_n784_), .ZN(G1337gat));
  AOI21_X1  g584(.A(new_n413_), .B1(new_n500_), .B2(new_n499_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n777_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n782_), .A2(new_n670_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n788_), .A2(KEYINPUT112), .A3(G99gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT112), .B1(new_n788_), .B2(G99gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n787_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n791_), .B(new_n793_), .ZN(G1338gat));
  INV_X1    g593(.A(G106gat), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n777_), .A2(new_n795_), .A3(new_n288_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n782_), .A2(new_n288_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(G106gat), .ZN(new_n799_));
  AOI211_X1 g598(.A(KEYINPUT52), .B(new_n795_), .C1(new_n782_), .C2(new_n288_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g601(.A(new_n601_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n592_), .A2(new_n589_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n804_), .B2(new_n595_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT114), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n803_), .C1(new_n804_), .C2(new_n595_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n596_), .A2(new_n592_), .A3(new_n595_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n806_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n605_), .B2(new_n604_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT115), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT115), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n810_), .B(new_n813_), .C1(new_n605_), .C2(new_n604_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n568_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n555_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n556_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n553_), .A2(KEYINPUT55), .A3(new_n555_), .A4(new_n554_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT56), .B1(new_n820_), .B2(new_n565_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n822_), .B(new_n566_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n815_), .B1(new_n821_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT58), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n815_), .B(KEYINPUT58), .C1(new_n821_), .C2(new_n823_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n826_), .A2(new_n651_), .A3(new_n827_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n610_), .B(new_n567_), .C1(new_n821_), .C2(new_n823_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n812_), .A2(new_n814_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(new_n572_), .A3(new_n570_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n540_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  XOR2_X1   g631(.A(KEYINPUT116), .B(KEYINPUT57), .Z(new_n833_));
  OAI21_X1  g632(.A(new_n828_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n834_), .A2(new_n835_), .B1(KEYINPUT57), .B2(new_n832_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n699_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n651_), .A2(new_n625_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n684_), .A3(new_n611_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(KEYINPUT54), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT54), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n652_), .A2(new_n842_), .A3(new_n611_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n838_), .A2(new_n845_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n391_), .A2(new_n444_), .A3(new_n670_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n829_), .A2(new_n831_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n540_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(KEYINPUT57), .A3(new_n851_), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n828_), .B(new_n852_), .C1(new_n832_), .C2(new_n833_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n625_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n844_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n855_), .A2(new_n847_), .ZN(new_n856_));
  OAI22_X1  g655(.A1(new_n846_), .A2(new_n849_), .B1(new_n848_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(G113gat), .B1(new_n857_), .B2(new_n611_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n856_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n611_), .A2(G113gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n858_), .B1(new_n859_), .B2(new_n860_), .ZN(G1340gat));
  XNOR2_X1  g660(.A(KEYINPUT118), .B(G120gat), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n684_), .A2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n856_), .B1(KEYINPUT60), .B2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n581_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n863_), .B1(new_n866_), .B2(new_n857_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n867_), .B1(KEYINPUT60), .B2(new_n865_), .ZN(G1341gat));
  AOI21_X1  g667(.A(G127gat), .B1(new_n856_), .B2(new_n699_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n857_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n699_), .A2(G127gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT119), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n869_), .B1(new_n870_), .B2(new_n872_), .ZN(G1342gat));
  OAI21_X1  g672(.A(G134gat), .B1(new_n857_), .B2(new_n692_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n851_), .A2(G134gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n859_), .B2(new_n875_), .ZN(G1343gat));
  AOI21_X1  g675(.A(new_n670_), .B1(new_n854_), .B2(new_n844_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n877_), .A2(new_n444_), .A3(new_n288_), .A4(new_n713_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(new_n611_), .ZN(new_n879_));
  XOR2_X1   g678(.A(KEYINPUT120), .B(G141gat), .Z(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1344gat));
  NOR2_X1   g680(.A1(new_n878_), .A2(new_n684_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT121), .B(G148gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1345gat));
  NOR2_X1   g683(.A1(new_n878_), .A2(new_n625_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT61), .B(G155gat), .Z(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1346gat));
  OAI21_X1  g686(.A(G162gat), .B1(new_n878_), .B2(new_n692_), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n851_), .A2(G162gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n878_), .B2(new_n889_), .ZN(G1347gat));
  NAND2_X1  g689(.A1(new_n662_), .A2(new_n445_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n846_), .A2(new_n288_), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n610_), .A2(new_n310_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT123), .Z(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n891_), .A2(new_n288_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n610_), .B(new_n896_), .C1(new_n838_), .C2(new_n845_), .ZN(new_n897_));
  XOR2_X1   g696(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n898_));
  AND3_X1   g697(.A1(new_n897_), .A2(G169gat), .A3(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n897_), .B2(G169gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n895_), .B1(new_n899_), .B2(new_n900_), .ZN(G1348gat));
  NAND2_X1  g700(.A1(new_n855_), .A2(new_n459_), .ZN(new_n902_));
  NOR4_X1   g701(.A1(new_n902_), .A2(new_n300_), .A3(new_n684_), .A4(new_n891_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n892_), .A2(new_n581_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n300_), .ZN(G1349gat));
  NOR3_X1   g704(.A1(new_n902_), .A2(new_n625_), .A3(new_n891_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT124), .ZN(new_n907_));
  OR2_X1    g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  AOI21_X1  g707(.A(G183gat), .B1(new_n906_), .B2(new_n907_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n625_), .A2(new_n303_), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n908_), .A2(new_n909_), .B1(new_n892_), .B2(new_n910_), .ZN(G1350gat));
  NAND2_X1  g710(.A1(new_n892_), .A2(new_n651_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(G190gat), .ZN(new_n913_));
  NAND3_X1  g712(.A1(new_n892_), .A2(new_n304_), .A3(new_n540_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1351gat));
  AOI22_X1  g714(.A1(new_n853_), .A2(new_n625_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n662_), .A2(new_n461_), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n916_), .A2(new_n917_), .A3(new_n670_), .A4(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n918_), .ZN(new_n920_));
  AOI21_X1  g719(.A(KEYINPUT125), .B1(new_n877_), .B2(new_n920_), .ZN(new_n921_));
  OAI211_X1 g720(.A(G197gat), .B(new_n610_), .C1(new_n919_), .C2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT126), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n855_), .A2(new_n413_), .A3(new_n920_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n917_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n877_), .A2(KEYINPUT125), .A3(new_n920_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n928_), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n610_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n610_), .B1(new_n919_), .B2(new_n921_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(new_n251_), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n924_), .A2(new_n929_), .A3(new_n931_), .ZN(G1352gat));
  AOI21_X1  g731(.A(new_n684_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(G204gat), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n253_), .A2(new_n255_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n934_), .B1(new_n935_), .B2(new_n933_), .ZN(G1353gat));
  AOI211_X1 g735(.A(KEYINPUT63), .B(G211gat), .C1(new_n928_), .C2(new_n699_), .ZN(new_n937_));
  XOR2_X1   g736(.A(KEYINPUT63), .B(G211gat), .Z(new_n938_));
  NAND3_X1  g737(.A1(new_n928_), .A2(new_n699_), .A3(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n939_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n937_), .A2(new_n940_), .ZN(G1354gat));
  AOI21_X1  g740(.A(G218gat), .B1(new_n928_), .B2(new_n540_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n651_), .A2(G218gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(KEYINPUT127), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n942_), .B1(new_n928_), .B2(new_n944_), .ZN(G1355gat));
endmodule


