//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n613_, new_n614_, new_n615_, new_n617_, new_n618_,
    new_n619_, new_n620_, new_n621_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n844_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  AND2_X1   g005(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G226gat), .A2(G233gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT20), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G211gat), .B(G218gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT91), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n214_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G197gat), .A2(G204gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT88), .B(G197gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n218_), .B1(new_n219_), .B2(G204gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT21), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT92), .B1(new_n217_), .B2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n213_), .B(KEYINPUT91), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT92), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(KEYINPUT21), .A4(new_n220_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT21), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n227_), .B1(G197gat), .B2(G204gat), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n228_), .B1(new_n219_), .B2(G204gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT89), .ZN(new_n230_));
  INV_X1    g029(.A(new_n220_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT90), .B(KEYINPUT21), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n231_), .A2(new_n232_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n226_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G169gat), .ZN(new_n241_));
  INV_X1    g040(.A(G176gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n243_), .A2(KEYINPUT24), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(KEYINPUT24), .A3(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n240_), .A2(new_n244_), .A3(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT26), .B(G190gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT75), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT25), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(new_n250_), .B2(G183gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT25), .B(G183gat), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n248_), .B(new_n251_), .C1(new_n252_), .C2(new_n249_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n238_), .B(new_n239_), .C1(G183gat), .C2(G190gat), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n254_), .A2(new_n245_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT22), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT76), .B1(new_n256_), .B2(G169gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT22), .B(G169gat), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n242_), .B(new_n257_), .C1(new_n258_), .C2(KEYINPUT76), .ZN(new_n259_));
  AOI22_X1  g058(.A1(new_n247_), .A2(new_n253_), .B1(new_n255_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n212_), .B1(new_n235_), .B2(new_n261_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n222_), .A2(new_n225_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n258_), .A2(new_n242_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(new_n254_), .A3(new_n245_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n248_), .A2(new_n252_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n266_), .A2(new_n240_), .A3(new_n244_), .A4(new_n246_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n263_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n211_), .B1(new_n262_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n226_), .A2(new_n234_), .A3(new_n260_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT20), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n226_), .A2(new_n234_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n211_), .A3(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n207_), .B1(new_n270_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n267_), .A2(new_n265_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT97), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n212_), .B1(new_n280_), .B2(new_n263_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT98), .ZN(new_n282_));
  OAI22_X1  g081(.A1(new_n281_), .A2(new_n282_), .B1(new_n263_), .B2(new_n260_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n278_), .B(KEYINPUT97), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT20), .B1(new_n235_), .B2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n285_), .A2(KEYINPUT98), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n211_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n287_));
  NOR3_X1   g086(.A1(new_n272_), .A2(new_n211_), .A3(new_n274_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n277_), .B1(new_n290_), .B2(new_n207_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G1gat), .B(G29gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(G85gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT0), .B(G57gat), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n293_), .B(new_n294_), .Z(new_n295_));
  XNOR2_X1  g094(.A(G127gat), .B(G134gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT79), .ZN(new_n297_));
  XOR2_X1   g096(.A(G113gat), .B(G120gat), .Z(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT83), .ZN(new_n301_));
  INV_X1    g100(.A(G155gat), .ZN(new_n302_));
  INV_X1    g101(.A(G162gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G155gat), .A2(G162gat), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT86), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT85), .B1(G141gat), .B2(G148gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NOR3_X1   g111(.A1(KEYINPUT85), .A2(G141gat), .A3(G148gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n309_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT85), .ZN(new_n315_));
  INV_X1    g114(.A(G141gat), .ZN(new_n316_));
  INV_X1    g115(.A(G148gat), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  NAND4_X1  g117(.A1(new_n318_), .A2(KEYINPUT86), .A3(new_n311_), .A4(new_n310_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n314_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n321_), .A2(KEYINPUT2), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(KEYINPUT2), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n316_), .A2(new_n317_), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n322_), .A2(new_n323_), .B1(KEYINPUT3), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT87), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n320_), .A2(KEYINPUT87), .A3(new_n325_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n308_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n324_), .A2(new_n321_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n307_), .A2(KEYINPUT1), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n307_), .A2(KEYINPUT1), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n306_), .A2(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n332_), .B1(new_n334_), .B2(KEYINPUT84), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n306_), .A2(new_n333_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT84), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n331_), .B1(new_n335_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n300_), .B1(new_n330_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n308_), .ZN(new_n341_));
  AND3_X1   g140(.A1(new_n320_), .A2(KEYINPUT87), .A3(new_n325_), .ZN(new_n342_));
  AOI21_X1  g141(.A(KEYINPUT87), .B1(new_n320_), .B2(new_n325_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n341_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n339_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n344_), .A2(new_n345_), .A3(new_n299_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n340_), .A2(KEYINPUT4), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT94), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n340_), .A2(new_n346_), .A3(KEYINPUT94), .A4(KEYINPUT4), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT95), .B(KEYINPUT4), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT96), .B1(new_n340_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n344_), .A2(new_n345_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT96), .ZN(new_n356_));
  INV_X1    g155(.A(new_n353_), .ZN(new_n357_));
  NAND4_X1  g156(.A1(new_n355_), .A2(new_n356_), .A3(new_n300_), .A4(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n352_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n351_), .A2(new_n359_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n340_), .A2(new_n346_), .A3(new_n352_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n295_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n295_), .ZN(new_n364_));
  AOI211_X1 g163(.A(new_n361_), .B(new_n364_), .C1(new_n351_), .C2(new_n359_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n291_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT99), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT28), .B1(new_n355_), .B2(KEYINPUT29), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n263_), .B1(new_n355_), .B2(KEYINPUT29), .ZN(new_n370_));
  NOR3_X1   g169(.A1(new_n355_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n371_));
  OR3_X1    g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G228gat), .A2(G233gat), .ZN(new_n374_));
  INV_X1    g173(.A(G78gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(G106gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G22gat), .B(G50gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n372_), .A2(new_n373_), .A3(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n380_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n365_), .A2(KEYINPUT33), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n270_), .A2(new_n276_), .A3(new_n205_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n272_), .A2(new_n210_), .A3(new_n274_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n206_), .B1(new_n269_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n385_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n352_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n351_), .A2(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n340_), .A2(new_n346_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n295_), .B1(new_n392_), .B2(new_n389_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n388_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n360_), .A2(new_n362_), .A3(new_n295_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT33), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n384_), .A2(new_n394_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT99), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n291_), .B(new_n399_), .C1(new_n363_), .C2(new_n365_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n367_), .A2(new_n383_), .A3(new_n398_), .A4(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G227gat), .A2(G233gat), .ZN(new_n402_));
  INV_X1    g201(.A(G15gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G71gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(G99gat), .ZN(new_n406_));
  INV_X1    g205(.A(G71gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n404_), .B(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(G99gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n406_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT77), .B(KEYINPUT30), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n412_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n406_), .A2(new_n410_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT78), .B(G43gat), .Z(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n260_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n260_), .A2(new_n418_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n416_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n299_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n421_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n413_), .A2(new_n425_), .A3(new_n419_), .A4(new_n415_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT81), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n422_), .A2(new_n424_), .A3(new_n426_), .A4(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n422_), .A2(new_n427_), .A3(new_n426_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n424_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n427_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n428_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n363_), .A2(new_n365_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n285_), .A2(KEYINPUT98), .B1(new_n235_), .B2(new_n261_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n281_), .A2(new_n282_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n210_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n205_), .B1(new_n439_), .B2(new_n288_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n387_), .A2(KEYINPUT27), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT27), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n440_), .A2(new_n441_), .B1(new_n388_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n436_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n383_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n435_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n401_), .A2(new_n446_), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n381_), .A2(new_n382_), .A3(new_n433_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(new_n436_), .A3(new_n443_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(KEYINPUT70), .B(G1gat), .Z(new_n451_));
  INV_X1    g250(.A(G8gat), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT14), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G15gat), .B(G22gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G1gat), .B(G8gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(G29gat), .B(G36gat), .Z(new_n458_));
  XOR2_X1   g257(.A(G43gat), .B(G50gat), .Z(new_n459_));
  XOR2_X1   g258(.A(new_n458_), .B(new_n459_), .Z(new_n460_));
  XNOR2_X1  g259(.A(new_n457_), .B(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(G229gat), .A3(G233gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n460_), .B(KEYINPUT15), .Z(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n457_), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n457_), .A2(new_n460_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G229gat), .A2(G233gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n466_), .B(KEYINPUT72), .Z(new_n467_));
  NAND3_X1  g266(.A1(new_n464_), .A2(new_n465_), .A3(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n462_), .A2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(G113gat), .B(G141gat), .Z(new_n470_));
  XNOR2_X1  g269(.A(G169gat), .B(G197gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n469_), .A2(new_n472_), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT73), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n473_), .A2(KEYINPUT73), .A3(new_n474_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n478_), .B(KEYINPUT74), .Z(new_n479_));
  NAND2_X1  g278(.A1(new_n450_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT100), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT100), .B1(new_n450_), .B2(new_n479_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G85gat), .B(G92gat), .Z(new_n485_));
  NOR2_X1   g284(.A1(G99gat), .A2(G106gat), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT7), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G99gat), .A2(G106gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT6), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n489_), .B(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n485_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT10), .B(G99gat), .Z(new_n495_));
  AOI22_X1  g294(.A1(KEYINPUT9), .A2(new_n485_), .B1(new_n495_), .B2(new_n377_), .ZN(new_n496_));
  INV_X1    g295(.A(G85gat), .ZN(new_n497_));
  INV_X1    g296(.A(G92gat), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n497_), .A2(new_n498_), .A3(KEYINPUT9), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n491_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n494_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n485_), .A2(KEYINPUT8), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT64), .ZN(new_n504_));
  OR2_X1    g303(.A1(new_n488_), .A2(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n491_), .B1(new_n488_), .B2(new_n504_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n503_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n502_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n463_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G232gat), .A2(G233gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT34), .ZN(new_n512_));
  OAI221_X1 g311(.A(new_n510_), .B1(KEYINPUT35), .B2(new_n512_), .C1(new_n460_), .C2(new_n509_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(KEYINPUT35), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n514_), .B(KEYINPUT68), .Z(new_n515_));
  XOR2_X1   g314(.A(new_n513_), .B(new_n515_), .Z(new_n516_));
  XNOR2_X1  g315(.A(G190gat), .B(G218gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G134gat), .B(G162gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n519_), .B(KEYINPUT36), .Z(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n513_), .B(new_n515_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n519_), .A2(KEYINPUT36), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(KEYINPUT37), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT69), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n521_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n516_), .A2(KEYINPUT69), .A3(new_n520_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n528_), .A2(new_n524_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT37), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n526_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  XOR2_X1   g331(.A(G71gat), .B(G78gat), .Z(new_n533_));
  XNOR2_X1  g332(.A(G57gat), .B(G64gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n533_), .B1(KEYINPUT11), .B2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT65), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(KEYINPUT11), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G231gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(new_n457_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT71), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G127gat), .B(G155gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT16), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G183gat), .B(G211gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT17), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n543_), .B(new_n548_), .ZN(new_n549_));
  OR3_X1    g348(.A1(new_n541_), .A2(KEYINPUT17), .A3(new_n547_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT66), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n552_), .B1(new_n538_), .B2(new_n509_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n537_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n536_), .B(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n555_), .A2(KEYINPUT66), .A3(new_n508_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n553_), .B(new_n556_), .C1(new_n508_), .C2(new_n555_), .ZN(new_n557_));
  AND2_X1   g356(.A1(G230gat), .A2(G233gat), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT12), .B1(new_n555_), .B2(new_n508_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n538_), .A2(new_n509_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n558_), .B1(new_n555_), .B2(new_n508_), .ZN(new_n563_));
  AOI22_X1  g362(.A1(new_n557_), .A2(new_n558_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G120gat), .B(G148gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT5), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G176gat), .B(G204gat), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n566_), .B(new_n567_), .Z(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT67), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n564_), .A2(new_n569_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT13), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n570_), .A2(KEYINPUT13), .A3(new_n571_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n532_), .A2(new_n551_), .A3(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n484_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n436_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n579_), .A2(new_n451_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT38), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT102), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n577_), .A2(new_n478_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n585_), .A2(KEYINPUT101), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(KEYINPUT101), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n449_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n589_), .B1(new_n401_), .B2(new_n446_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n530_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n551_), .ZN(new_n594_));
  NOR3_X1   g393(.A1(new_n588_), .A2(new_n593_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(new_n580_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(G1gat), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n584_), .B(new_n597_), .C1(new_n582_), .C2(new_n581_), .ZN(G1324gat));
  INV_X1    g397(.A(new_n443_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n579_), .A2(new_n452_), .A3(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n595_), .A2(new_n599_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n601_), .B1(new_n602_), .B2(G8gat), .ZN(new_n603_));
  AOI211_X1 g402(.A(KEYINPUT39), .B(new_n452_), .C1(new_n595_), .C2(new_n599_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n600_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT104), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT104), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n607_), .B(new_n600_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n606_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n609_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(G1325gat));
  AOI21_X1  g411(.A(new_n403_), .B1(new_n595_), .B2(new_n435_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT41), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n579_), .A2(new_n403_), .A3(new_n435_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(G1326gat));
  INV_X1    g415(.A(G22gat), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n383_), .B(KEYINPUT105), .Z(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n595_), .B2(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT42), .Z(new_n620_));
  NAND3_X1  g419(.A1(new_n579_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(G1327gat));
  XNOR2_X1  g421(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n623_));
  OAI21_X1  g422(.A(KEYINPUT43), .B1(new_n590_), .B2(new_n532_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n590_), .A2(KEYINPUT43), .A3(new_n532_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n625_), .B2(KEYINPUT106), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT43), .ZN(new_n627_));
  INV_X1    g426(.A(new_n532_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n450_), .A2(KEYINPUT106), .A3(new_n627_), .A4(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n626_), .A2(new_n630_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n586_), .A2(new_n594_), .A3(new_n587_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n623_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT44), .ZN(new_n635_));
  OAI211_X1 g434(.A(new_n635_), .B(new_n632_), .C1(new_n626_), .C2(new_n630_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n436_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(G29gat), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n594_), .A2(new_n591_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n639_), .A2(new_n576_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT108), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI211_X1 g442(.A(KEYINPUT108), .B(new_n640_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n580_), .A2(new_n638_), .ZN(new_n646_));
  OAI22_X1  g445(.A1(new_n637_), .A2(new_n638_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT109), .Z(G1328gat));
  NOR2_X1   g447(.A1(new_n443_), .A2(G36gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n643_), .A2(new_n644_), .A3(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT45), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT45), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n643_), .A2(new_n652_), .A3(new_n644_), .A4(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT110), .ZN(new_n656_));
  INV_X1    g455(.A(new_n636_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n623_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n450_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n629_), .A3(new_n624_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n658_), .B1(new_n662_), .B2(new_n632_), .ZN(new_n663_));
  OAI211_X1 g462(.A(new_n656_), .B(new_n599_), .C1(new_n657_), .C2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G36gat), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n634_), .A2(new_n636_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n656_), .B1(new_n666_), .B2(new_n599_), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n654_), .B(new_n655_), .C1(new_n665_), .C2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n599_), .B1(new_n657_), .B2(new_n663_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT110), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(G36gat), .A3(new_n664_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n655_), .B1(new_n672_), .B2(new_n654_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n669_), .A2(new_n673_), .ZN(G1329gat));
  AOI21_X1  g473(.A(new_n433_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n675_));
  INV_X1    g474(.A(G43gat), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n435_), .A2(new_n676_), .ZN(new_n677_));
  OAI22_X1  g476(.A1(new_n675_), .A2(new_n676_), .B1(new_n645_), .B2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n678_), .B(new_n679_), .Z(G1330gat));
  INV_X1    g479(.A(G50gat), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n383_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n643_), .A2(new_n618_), .A3(new_n644_), .ZN(new_n683_));
  AOI22_X1  g482(.A1(new_n666_), .A2(new_n682_), .B1(new_n683_), .B2(new_n681_), .ZN(G1331gat));
  NAND3_X1  g483(.A1(new_n532_), .A2(new_n551_), .A3(new_n576_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT113), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n590_), .A2(new_n478_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(G57gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n688_), .A2(new_n689_), .A3(new_n580_), .ZN(new_n690_));
  NOR4_X1   g489(.A1(new_n593_), .A2(new_n479_), .A3(new_n594_), .A4(new_n577_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n691_), .A2(new_n580_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n690_), .B1(new_n692_), .B2(new_n689_), .ZN(G1332gat));
  INV_X1    g492(.A(G64gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n691_), .B2(new_n599_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT48), .Z(new_n696_));
  NAND3_X1  g495(.A1(new_n688_), .A2(new_n694_), .A3(new_n599_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1333gat));
  AOI21_X1  g497(.A(new_n407_), .B1(new_n691_), .B2(new_n435_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT49), .Z(new_n700_));
  NAND3_X1  g499(.A1(new_n688_), .A2(new_n407_), .A3(new_n435_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(G1334gat));
  AOI21_X1  g501(.A(new_n375_), .B1(new_n691_), .B2(new_n618_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT50), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n688_), .A2(new_n375_), .A3(new_n618_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1335gat));
  NAND4_X1  g505(.A1(new_n687_), .A2(new_n591_), .A3(new_n594_), .A4(new_n576_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n497_), .B1(new_n707_), .B2(new_n436_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT114), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n577_), .A2(new_n551_), .A3(new_n478_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n662_), .A2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n436_), .A2(new_n497_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT115), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n709_), .B1(new_n711_), .B2(new_n713_), .ZN(G1336gat));
  INV_X1    g513(.A(new_n707_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n498_), .A3(new_n599_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n711_), .A2(new_n599_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n718_), .B2(new_n498_), .ZN(G1337gat));
  INV_X1    g518(.A(new_n433_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n715_), .A2(new_n720_), .A3(new_n495_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n711_), .A2(new_n435_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(G99gat), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT118), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT117), .B(KEYINPUT51), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n723_), .A2(new_n724_), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n724_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT116), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n723_), .A2(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT51), .B1(new_n723_), .B2(new_n728_), .ZN(new_n730_));
  OAI22_X1  g529(.A1(new_n726_), .A2(new_n727_), .B1(new_n729_), .B2(new_n730_), .ZN(G1338gat));
  NAND3_X1  g530(.A1(new_n715_), .A2(new_n377_), .A3(new_n445_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT52), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n711_), .A2(new_n445_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(G106gat), .ZN(new_n735_));
  AOI211_X1 g534(.A(KEYINPUT52), .B(new_n377_), .C1(new_n711_), .C2(new_n445_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g537(.A1(new_n599_), .A2(new_n436_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n720_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n568_), .ZN(new_n742_));
  AOI22_X1  g541(.A1(new_n476_), .A2(new_n477_), .B1(new_n564_), .B2(new_n742_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n555_), .A2(KEYINPUT12), .A3(new_n508_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n560_), .B1(new_n538_), .B2(new_n509_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n553_), .A2(new_n556_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n558_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT55), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n749_), .B(new_n563_), .C1(new_n744_), .C2(new_n745_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT119), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n562_), .A2(new_n563_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT55), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(new_n750_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT119), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(new_n758_), .A3(new_n748_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n742_), .B1(new_n754_), .B2(new_n759_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(KEYINPUT56), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  AOI211_X1 g561(.A(new_n762_), .B(new_n742_), .C1(new_n754_), .C2(new_n759_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n743_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n472_), .B1(new_n461_), .B2(new_n467_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n467_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n464_), .A2(new_n465_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n474_), .A2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n769_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n764_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT57), .B1(new_n772_), .B2(new_n530_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n774_), .B(new_n591_), .C1(new_n764_), .C2(new_n771_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n753_), .A2(KEYINPUT119), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n758_), .B1(new_n757_), .B2(new_n748_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n568_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n779_), .A2(KEYINPUT120), .A3(new_n762_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT120), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n760_), .B2(KEYINPUT56), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n760_), .A2(KEYINPUT56), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n780_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n769_), .B1(new_n564_), .B2(new_n742_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n784_), .A2(KEYINPUT58), .A3(new_n785_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n788_), .A2(new_n628_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n551_), .B1(new_n776_), .B2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n578_), .A2(new_n479_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT54), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n383_), .B(new_n741_), .C1(new_n791_), .C2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(G113gat), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(new_n478_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n479_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT121), .ZN(new_n799_));
  INV_X1    g598(.A(new_n789_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT58), .B1(new_n784_), .B2(new_n785_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n532_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n564_), .A2(new_n742_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n477_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n804_), .B2(new_n475_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n779_), .A2(new_n762_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n783_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n530_), .B1(new_n807_), .B2(new_n770_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n774_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n772_), .A2(KEYINPUT57), .A3(new_n530_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n594_), .B1(new_n802_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n792_), .B(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n445_), .B1(new_n812_), .B2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(KEYINPUT59), .B1(new_n815_), .B2(new_n741_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT59), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n794_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n799_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n815_), .A2(KEYINPUT59), .A3(new_n741_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n794_), .A2(new_n817_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(KEYINPUT121), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n798_), .B1(new_n819_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n797_), .B1(new_n823_), .B2(new_n796_), .ZN(G1340gat));
  AOI21_X1  g623(.A(new_n577_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n825_));
  INV_X1    g624(.A(G120gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n577_), .B2(KEYINPUT60), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(KEYINPUT60), .B2(new_n826_), .ZN(new_n828_));
  OAI22_X1  g627(.A1(new_n825_), .A2(new_n826_), .B1(new_n794_), .B2(new_n828_), .ZN(G1341gat));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n795_), .A2(new_n830_), .A3(new_n551_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n594_), .B1(new_n819_), .B2(new_n822_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n830_), .ZN(G1342gat));
  INV_X1    g632(.A(G134gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n795_), .A2(new_n834_), .A3(new_n591_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n532_), .B1(new_n819_), .B2(new_n822_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n834_), .ZN(G1343gat));
  NAND2_X1  g636(.A1(new_n812_), .A2(new_n814_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n435_), .A2(new_n383_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n739_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n478_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g642(.A1(new_n840_), .A2(new_n577_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT122), .B(G148gat), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1345gat));
  OR3_X1    g645(.A1(new_n840_), .A2(KEYINPUT123), .A3(new_n594_), .ZN(new_n847_));
  OAI21_X1  g646(.A(KEYINPUT123), .B1(new_n840_), .B2(new_n594_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT61), .B(G155gat), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n847_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1346gat));
  OAI21_X1  g651(.A(G162gat), .B1(new_n840_), .B2(new_n532_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n591_), .A2(new_n303_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n840_), .B2(new_n854_), .ZN(G1347gat));
  INV_X1    g654(.A(KEYINPUT62), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n435_), .A2(new_n599_), .A3(new_n436_), .ZN(new_n857_));
  XOR2_X1   g656(.A(new_n857_), .B(KEYINPUT124), .Z(new_n858_));
  NOR2_X1   g657(.A1(new_n858_), .A2(new_n618_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n838_), .A2(new_n478_), .A3(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n861_));
  OAI21_X1  g660(.A(G169gat), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n861_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n856_), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n864_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n866_), .A2(new_n862_), .A3(KEYINPUT62), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n838_), .A2(new_n859_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n478_), .A2(new_n258_), .ZN(new_n869_));
  XOR2_X1   g668(.A(new_n869_), .B(KEYINPUT126), .Z(new_n870_));
  OAI22_X1  g669(.A1(new_n865_), .A2(new_n867_), .B1(new_n868_), .B2(new_n870_), .ZN(G1348gat));
  INV_X1    g670(.A(new_n815_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n872_), .A2(new_n577_), .A3(new_n858_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n576_), .A2(new_n242_), .ZN(new_n874_));
  OAI22_X1  g673(.A1(new_n873_), .A2(new_n242_), .B1(new_n868_), .B2(new_n874_), .ZN(G1349gat));
  NOR3_X1   g674(.A1(new_n868_), .A2(new_n252_), .A3(new_n594_), .ZN(new_n876_));
  OR3_X1    g675(.A1(new_n872_), .A2(new_n594_), .A3(new_n858_), .ZN(new_n877_));
  INV_X1    g676(.A(G183gat), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n877_), .B2(new_n878_), .ZN(G1350gat));
  OAI21_X1  g678(.A(G190gat), .B1(new_n868_), .B2(new_n532_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n591_), .A2(new_n248_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n868_), .B2(new_n881_), .ZN(G1351gat));
  NAND2_X1  g681(.A1(new_n839_), .A2(new_n436_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n599_), .B1(new_n883_), .B2(KEYINPUT127), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n884_), .B1(KEYINPUT127), .B2(new_n883_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n838_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n478_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n576_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g689(.A1(new_n886_), .A2(new_n551_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n892_));
  AND2_X1   g691(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n891_), .A2(new_n892_), .A3(new_n893_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n891_), .B2(new_n892_), .ZN(G1354gat));
  INV_X1    g694(.A(G218gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n886_), .A2(new_n896_), .A3(new_n591_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n886_), .A2(new_n628_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n896_), .ZN(G1355gat));
endmodule


