//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n203_), .B(KEYINPUT96), .Z(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(G169gat), .ZN(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT23), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT87), .ZN(new_n211_));
  NOR3_X1   g010(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT23), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n207_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(KEYINPUT97), .B(KEYINPUT24), .Z(new_n216_));
  INV_X1    g015(.A(G169gat), .ZN(new_n217_));
  INV_X1    g016(.A(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n212_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(new_n210_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT25), .B(G183gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(KEYINPUT26), .B(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G169gat), .B(G176gat), .Z(new_n226_));
  NAND2_X1  g025(.A1(new_n216_), .A2(new_n226_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n220_), .A2(new_n222_), .A3(new_n225_), .A4(new_n227_), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n215_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT21), .ZN(new_n230_));
  INV_X1    g029(.A(G197gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G204gat), .ZN(new_n232_));
  INV_X1    g031(.A(G204gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G197gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n230_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT91), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G211gat), .B(G218gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT92), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(new_n233_), .B2(G197gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n231_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n239_), .A2(new_n234_), .A3(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n237_), .B1(new_n241_), .B2(KEYINPUT21), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n236_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n237_), .A2(new_n230_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n244_), .A2(new_n241_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n229_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT20), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n222_), .B1(G183gat), .B2(G190gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n207_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(new_n226_), .B2(KEYINPUT24), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n225_), .B(new_n252_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n250_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n248_), .B1(new_n255_), .B2(new_n246_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n205_), .B1(new_n247_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n248_), .B1(new_n229_), .B2(new_n246_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n203_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n254_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(G8gat), .B(G36gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT18), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G64gat), .B(G92gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n264_), .B(new_n265_), .Z(new_n266_));
  NAND3_X1  g065(.A1(new_n258_), .A2(new_n262_), .A3(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n266_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n268_), .B1(new_n269_), .B2(new_n257_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT27), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT102), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT102), .ZN(new_n274_));
  AOI211_X1 g073(.A(new_n274_), .B(KEYINPUT27), .C1(new_n267_), .C2(new_n270_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n247_), .A2(new_n205_), .A3(new_n256_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n260_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n268_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n267_), .A2(new_n279_), .A3(KEYINPUT27), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT103), .B1(new_n276_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT103), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n283_), .B(new_n280_), .C1(new_n273_), .C2(new_n275_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT95), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G228gat), .A2(G233gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n287_), .B(KEYINPUT90), .Z(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(new_n289_), .A2(KEYINPUT93), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  NOR2_X1   g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n294_), .B(KEYINPUT3), .Z(new_n295_));
  NAND2_X1  g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n296_), .B(KEYINPUT2), .Z(new_n297_));
  OAI211_X1 g096(.A(new_n291_), .B(new_n293_), .C1(new_n295_), .C2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n292_), .B1(KEYINPUT1), .B2(new_n291_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n299_), .B1(KEYINPUT1), .B2(new_n291_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n294_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n296_), .A3(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n298_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n290_), .B1(new_n305_), .B2(new_n246_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(G78gat), .ZN(new_n307_));
  INV_X1    g106(.A(G78gat), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n308_), .B(new_n290_), .C1(new_n305_), .C2(new_n246_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n289_), .A2(KEYINPUT93), .ZN(new_n311_));
  INV_X1    g110(.A(G106gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n307_), .A2(new_n309_), .A3(new_n313_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(G22gat), .B(G50gat), .Z(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n303_), .A2(new_n304_), .A3(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n321_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n319_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n303_), .A2(new_n304_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n320_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n303_), .A2(new_n304_), .A3(new_n321_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n318_), .A3(new_n327_), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n324_), .A2(new_n328_), .A3(KEYINPUT89), .ZN(new_n329_));
  AOI21_X1  g128(.A(KEYINPUT89), .B1(new_n324_), .B2(new_n328_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n317_), .A2(KEYINPUT94), .A3(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n324_), .A2(new_n328_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n315_), .A2(new_n316_), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(KEYINPUT94), .B1(new_n317_), .B2(new_n331_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n286_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n317_), .A2(new_n331_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT94), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n340_), .A2(KEYINPUT95), .A3(new_n332_), .A4(new_n334_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G225gat), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G127gat), .B(G134gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G113gat), .B(G120gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n303_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n303_), .A2(new_n347_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(KEYINPUT4), .A3(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n303_), .A2(new_n347_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT100), .ZN(new_n352_));
  XOR2_X1   g151(.A(KEYINPUT99), .B(KEYINPUT4), .Z(new_n353_));
  AND3_X1   g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n352_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n344_), .B(new_n350_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n348_), .A2(new_n349_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n343_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360_));
  INV_X1    g159(.A(G85gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT0), .B(G57gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n359_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n356_), .A2(new_n364_), .A3(new_n358_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G71gat), .B(G99gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G43gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n254_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(new_n347_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G227gat), .A2(G233gat), .ZN(new_n374_));
  INV_X1    g173(.A(G15gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT30), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT31), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n373_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n369_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n285_), .A2(new_n342_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n271_), .A2(KEYINPUT98), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT98), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n267_), .A2(new_n270_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n364_), .B1(new_n357_), .B2(new_n344_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n350_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n386_), .B1(new_n387_), .B2(new_n344_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n367_), .A2(KEYINPUT33), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n383_), .A2(new_n385_), .A3(new_n388_), .A4(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT33), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n366_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT101), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n266_), .A2(KEYINPUT32), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n258_), .A2(new_n262_), .A3(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n277_), .A2(new_n278_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n395_), .B1(new_n396_), .B2(new_n394_), .ZN(new_n397_));
  OAI22_X1  g196(.A1(new_n390_), .A2(new_n393_), .B1(new_n368_), .B2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n369_), .B1(new_n337_), .B2(new_n341_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n276_), .A2(new_n281_), .ZN(new_n400_));
  AOI22_X1  g199(.A1(new_n342_), .A2(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n382_), .B1(new_n401_), .B2(new_n379_), .ZN(new_n402_));
  INV_X1    g201(.A(G230gat), .ZN(new_n403_));
  INV_X1    g202(.A(G233gat), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(G99gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n406_), .A2(new_n312_), .A3(KEYINPUT65), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT65), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(G99gat), .B2(G106gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT7), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT66), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT66), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT7), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n407_), .A2(new_n409_), .A3(new_n411_), .A4(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT64), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OAI211_X1 g216(.A(KEYINPUT64), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G99gat), .A2(G106gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT6), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(G99gat), .A3(G106gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n414_), .A2(new_n419_), .A3(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT67), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT8), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT67), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n414_), .A2(new_n419_), .A3(new_n428_), .A4(new_n424_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G85gat), .B(G92gat), .Z(new_n430_));
  NAND4_X1  g229(.A1(new_n426_), .A2(new_n427_), .A3(new_n429_), .A4(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n422_), .B1(G99gat), .B2(G106gat), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n420_), .A2(KEYINPUT6), .ZN(new_n433_));
  OAI21_X1  g232(.A(KEYINPUT68), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT68), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n421_), .A2(new_n423_), .A3(new_n435_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n434_), .A2(new_n419_), .A3(new_n414_), .A4(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT69), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(new_n430_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT8), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n438_), .B1(new_n437_), .B2(new_n430_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n431_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G57gat), .B(G64gat), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n443_), .A2(KEYINPUT11), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(KEYINPUT11), .ZN(new_n445_));
  XOR2_X1   g244(.A(G71gat), .B(G78gat), .Z(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  OR2_X1    g246(.A1(new_n445_), .A2(new_n446_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  XOR2_X1   g248(.A(KEYINPUT10), .B(G99gat), .Z(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n312_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n430_), .A2(KEYINPUT9), .ZN(new_n452_));
  INV_X1    g251(.A(G92gat), .ZN(new_n453_));
  OR3_X1    g252(.A1(new_n361_), .A2(new_n453_), .A3(KEYINPUT9), .ZN(new_n454_));
  NAND4_X1  g253(.A1(new_n451_), .A2(new_n452_), .A3(new_n424_), .A4(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n442_), .A2(new_n449_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT70), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n442_), .A2(new_n455_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n449_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n456_), .A2(new_n457_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n405_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT12), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n405_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n456_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n455_), .B(KEYINPUT71), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n442_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(KEYINPUT12), .A3(new_n460_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n466_), .A2(new_n468_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n464_), .A2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G176gat), .B(G204gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT74), .ZN(new_n475_));
  XOR2_X1   g274(.A(G120gat), .B(G148gat), .Z(new_n476_));
  XOR2_X1   g275(.A(new_n475_), .B(new_n476_), .Z(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n477_), .B(new_n478_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n479_), .A2(KEYINPUT72), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n473_), .B(new_n480_), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n481_), .A2(KEYINPUT13), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(KEYINPUT13), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G229gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G29gat), .B(G36gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G43gat), .B(G50gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT15), .ZN(new_n489_));
  OR2_X1    g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G15gat), .B(G22gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G1gat), .B(G8gat), .ZN(new_n492_));
  INV_X1    g291(.A(G1gat), .ZN(new_n493_));
  OR2_X1    g292(.A1(KEYINPUT81), .A2(G8gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(KEYINPUT81), .A2(G8gat), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT14), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n491_), .B(new_n492_), .C1(new_n496_), .C2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n491_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n492_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n488_), .A2(new_n489_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n490_), .A2(new_n498_), .A3(new_n501_), .A4(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n498_), .ZN(new_n504_));
  AND2_X1   g303(.A1(KEYINPUT81), .A2(G8gat), .ZN(new_n505_));
  NOR2_X1   g304(.A1(KEYINPUT81), .A2(G8gat), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT14), .B1(new_n507_), .B2(new_n493_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n492_), .B1(new_n508_), .B2(new_n491_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n488_), .B1(new_n504_), .B2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(KEYINPUT85), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT85), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n501_), .A2(new_n498_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n512_), .B1(new_n513_), .B2(new_n488_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n485_), .B(new_n503_), .C1(new_n511_), .C2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G113gat), .B(G141gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G169gat), .B(G197gat), .ZN(new_n517_));
  XOR2_X1   g316(.A(new_n516_), .B(new_n517_), .Z(new_n518_));
  NOR2_X1   g317(.A1(new_n513_), .A2(new_n488_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n510_), .A2(KEYINPUT85), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n513_), .A2(new_n512_), .A3(new_n488_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n515_), .B(new_n518_), .C1(new_n485_), .C2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT86), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n485_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n511_), .A2(new_n514_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n526_), .B1(new_n527_), .B2(new_n519_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n528_), .A2(KEYINPUT86), .A3(new_n515_), .A4(new_n518_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n528_), .A2(new_n515_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n518_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n484_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT84), .ZN(new_n537_));
  XOR2_X1   g336(.A(G127gat), .B(G155gat), .Z(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT16), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G183gat), .B(G211gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT17), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n537_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(new_n460_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(new_n513_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT82), .B(KEYINPUT83), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G231gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n548_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n541_), .A2(new_n542_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G190gat), .B(G218gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT77), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G134gat), .B(G162gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n558_), .A2(KEYINPUT36), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n442_), .A2(new_n488_), .A3(new_n455_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G232gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT35), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT71), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n455_), .B(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n437_), .A2(new_n430_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT69), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT8), .A3(new_n439_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n568_), .B1(new_n571_), .B2(new_n431_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n490_), .A2(new_n502_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n560_), .B(new_n566_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT76), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n564_), .A2(new_n565_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n573_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n470_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT76), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n578_), .A2(new_n579_), .A3(new_n560_), .A4(new_n566_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n575_), .A2(new_n576_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n576_), .B1(new_n575_), .B2(new_n580_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n559_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n576_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n580_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n470_), .A2(new_n577_), .B1(new_n565_), .B2(new_n564_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n579_), .B1(new_n586_), .B2(new_n560_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n584_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n575_), .A2(new_n576_), .A3(new_n580_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n557_), .B(KEYINPUT36), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n583_), .A2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT80), .B1(new_n592_), .B2(KEYINPUT37), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT80), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT37), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n583_), .A2(new_n591_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n590_), .B(KEYINPUT78), .Z(new_n598_));
  NAND3_X1  g397(.A1(new_n588_), .A2(new_n589_), .A3(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n583_), .A2(new_n599_), .A3(KEYINPUT79), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n600_), .B(KEYINPUT37), .C1(KEYINPUT79), .C2(new_n599_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n553_), .B1(new_n597_), .B2(new_n601_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n402_), .A2(new_n536_), .A3(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n493_), .A3(new_n369_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT38), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n342_), .A2(new_n398_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n399_), .A2(new_n400_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n337_), .A2(new_n341_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n610_));
  AOI22_X1  g409(.A1(new_n608_), .A2(new_n380_), .B1(new_n610_), .B2(new_n381_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n592_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n611_), .A2(new_n553_), .A3(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n536_), .B(KEYINPUT104), .Z(new_n614_));
  AND2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G1gat), .B1(new_n616_), .B2(new_n368_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n605_), .A2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT105), .Z(G1324gat));
  INV_X1    g418(.A(new_n285_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n603_), .A2(new_n507_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n615_), .A2(new_n620_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n622_), .A2(new_n623_), .A3(G8gat), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n623_), .B1(new_n622_), .B2(G8gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n621_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(KEYINPUT40), .B(new_n621_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1325gat));
  AOI21_X1  g429(.A(new_n375_), .B1(new_n615_), .B2(new_n379_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT41), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n603_), .A2(new_n375_), .A3(new_n379_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1326gat));
  INV_X1    g433(.A(G22gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n615_), .B2(new_n609_), .ZN(new_n636_));
  XOR2_X1   g435(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n603_), .A2(new_n635_), .A3(new_n609_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(G1327gat));
  NOR2_X1   g439(.A1(new_n552_), .A2(new_n592_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n402_), .A2(new_n536_), .A3(new_n641_), .ZN(new_n642_));
  OR3_X1    g441(.A1(new_n642_), .A2(G29gat), .A3(new_n368_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n597_), .A2(new_n601_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n402_), .A2(KEYINPUT107), .A3(KEYINPUT43), .A4(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n646_), .A2(new_n553_), .ZN(new_n647_));
  OR2_X1    g446(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n648_));
  NAND2_X1  g447(.A1(KEYINPUT107), .A2(KEYINPUT43), .ZN(new_n649_));
  OAI211_X1 g448(.A(new_n648_), .B(new_n649_), .C1(new_n611_), .C2(new_n644_), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n647_), .A2(KEYINPUT44), .A3(new_n614_), .A4(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n650_), .A2(new_n646_), .A3(new_n614_), .A4(new_n553_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n651_), .A2(new_n654_), .A3(new_n369_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n655_), .A2(KEYINPUT108), .A3(G29gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(KEYINPUT108), .B1(new_n655_), .B2(G29gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n643_), .B1(new_n656_), .B2(new_n657_), .ZN(G1328gat));
  NAND3_X1  g457(.A1(new_n651_), .A2(new_n654_), .A3(new_n620_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G36gat), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n642_), .A2(G36gat), .A3(new_n285_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n660_), .A2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n660_), .A2(new_n663_), .A3(new_n665_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(G1329gat));
  INV_X1    g468(.A(G43gat), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n380_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n651_), .A2(new_n654_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(KEYINPUT111), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT111), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n651_), .A2(new_n654_), .A3(new_n674_), .A4(new_n671_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n670_), .B1(new_n642_), .B2(new_n380_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n673_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(KEYINPUT47), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT47), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n673_), .A2(new_n679_), .A3(new_n675_), .A4(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1330gat));
  NAND4_X1  g480(.A1(new_n651_), .A2(new_n654_), .A3(G50gat), .A4(new_n609_), .ZN(new_n682_));
  INV_X1    g481(.A(G50gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n683_), .B1(new_n642_), .B2(new_n342_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n682_), .A2(new_n684_), .ZN(G1331gat));
  INV_X1    g484(.A(new_n484_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(new_n534_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n402_), .A2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(new_n602_), .ZN(new_n689_));
  INV_X1    g488(.A(G57gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n690_), .A3(new_n369_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n613_), .A2(new_n687_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G57gat), .B1(new_n692_), .B2(new_n368_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1332gat));
  OAI21_X1  g493(.A(G64gat), .B1(new_n692_), .B2(new_n285_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT48), .ZN(new_n696_));
  INV_X1    g495(.A(G64gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n689_), .A2(new_n697_), .A3(new_n620_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT112), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n696_), .A2(KEYINPUT112), .A3(new_n698_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1333gat));
  OAI21_X1  g502(.A(G71gat), .B1(new_n692_), .B2(new_n380_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT49), .ZN(new_n705_));
  INV_X1    g504(.A(G71gat), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n689_), .A2(new_n706_), .A3(new_n379_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1334gat));
  OAI21_X1  g507(.A(G78gat), .B1(new_n692_), .B2(new_n342_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT50), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n689_), .A2(new_n308_), .A3(new_n609_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1335gat));
  NAND2_X1  g511(.A1(new_n688_), .A2(new_n641_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(new_n361_), .A3(new_n369_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n650_), .A2(new_n646_), .A3(new_n553_), .A4(new_n687_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n716_), .A2(KEYINPUT113), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(KEYINPUT113), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n717_), .A2(new_n369_), .A3(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n715_), .B1(new_n719_), .B2(new_n361_), .ZN(G1336gat));
  NAND3_X1  g519(.A1(new_n714_), .A2(new_n453_), .A3(new_n620_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n717_), .A2(new_n620_), .A3(new_n718_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(new_n453_), .ZN(G1337gat));
  OAI21_X1  g522(.A(G99gat), .B1(new_n716_), .B2(new_n380_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n714_), .A2(new_n450_), .A3(new_n379_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(KEYINPUT114), .A2(KEYINPUT51), .ZN(new_n727_));
  XOR2_X1   g526(.A(new_n726_), .B(new_n727_), .Z(G1338gat));
  NAND3_X1  g527(.A1(new_n714_), .A2(new_n312_), .A3(new_n609_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n716_), .A2(new_n342_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n731_), .B2(G106gat), .ZN(new_n732_));
  OAI211_X1 g531(.A(G106gat), .B(new_n730_), .C1(new_n716_), .C2(new_n342_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n729_), .B1(new_n732_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT53), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n737_), .B(new_n729_), .C1(new_n732_), .C2(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1339gat));
  INV_X1    g538(.A(KEYINPUT119), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n464_), .A2(new_n472_), .A3(new_n479_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n503_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n527_), .A2(new_n742_), .A3(new_n485_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n532_), .B1(new_n522_), .B2(new_n526_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n525_), .B2(new_n529_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n741_), .A2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n449_), .B1(new_n442_), .B2(new_n455_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n460_), .A2(KEYINPUT12), .ZN(new_n749_));
  OAI22_X1  g548(.A1(new_n748_), .A2(KEYINPUT12), .B1(new_n572_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n456_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n405_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n456_), .A2(new_n467_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n750_), .B2(new_n754_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n466_), .A2(new_n468_), .A3(KEYINPUT55), .A4(new_n471_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n752_), .A2(new_n755_), .A3(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n479_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(KEYINPUT56), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT56), .B1(new_n757_), .B2(new_n758_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n747_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT58), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n747_), .B(KEYINPUT58), .C1(new_n760_), .C2(new_n761_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n597_), .A2(new_n764_), .A3(new_n601_), .A4(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n746_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n481_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n757_), .A2(new_n758_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT56), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n761_), .A2(KEYINPUT117), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n759_), .ZN(new_n776_));
  AND3_X1   g575(.A1(new_n741_), .A2(new_n534_), .A3(KEYINPUT116), .ZN(new_n777_));
  AOI21_X1  g576(.A(KEYINPUT116), .B1(new_n741_), .B2(new_n534_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n769_), .B1(new_n776_), .B2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT57), .B1(new_n780_), .B2(new_n612_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n759_), .B1(new_n761_), .B2(KEYINPUT117), .ZN(new_n782_));
  AOI211_X1 g581(.A(new_n773_), .B(KEYINPUT56), .C1(new_n757_), .C2(new_n758_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n481_), .A2(new_n768_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT57), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n786_), .A2(new_n787_), .A3(new_n592_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n767_), .B1(new_n781_), .B2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n740_), .B1(new_n789_), .B2(new_n552_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT54), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n484_), .A2(new_n534_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n792_), .B2(new_n602_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n602_), .A3(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n787_), .B1(new_n786_), .B2(new_n592_), .ZN(new_n797_));
  AOI211_X1 g596(.A(KEYINPUT57), .B(new_n612_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n766_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(KEYINPUT119), .A3(new_n553_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n790_), .A2(new_n796_), .A3(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n610_), .A2(new_n369_), .A3(new_n379_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n802_), .A2(KEYINPUT59), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n799_), .A2(KEYINPUT118), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT118), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n806_), .B(new_n766_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n805_), .A2(new_n553_), .A3(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n802_), .B1(new_n808_), .B2(new_n796_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT59), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n804_), .B(new_n534_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G113gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n553_), .B1(new_n789_), .B2(new_n806_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n807_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n796_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n802_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OR3_X1    g616(.A1(new_n817_), .A2(G113gat), .A3(new_n535_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n812_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT120), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n812_), .A2(new_n821_), .A3(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(G1340gat));
  NAND2_X1  g622(.A1(new_n817_), .A2(KEYINPUT59), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n804_), .ZN(new_n825_));
  OAI21_X1  g624(.A(G120gat), .B1(new_n825_), .B2(new_n686_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT60), .ZN(new_n827_));
  AOI21_X1  g626(.A(G120gat), .B1(new_n484_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT121), .B1(new_n827_), .B2(G120gat), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n828_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n826_), .B1(new_n817_), .B2(new_n832_), .ZN(G1341gat));
  AOI21_X1  g632(.A(G127gat), .B1(new_n809_), .B2(new_n552_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n825_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n552_), .A2(G127gat), .ZN(new_n836_));
  XOR2_X1   g635(.A(new_n836_), .B(KEYINPUT122), .Z(new_n837_));
  AOI21_X1  g636(.A(new_n834_), .B1(new_n835_), .B2(new_n837_), .ZN(G1342gat));
  OAI21_X1  g637(.A(G134gat), .B1(new_n825_), .B2(new_n644_), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n592_), .A2(G134gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n817_), .B2(new_n840_), .ZN(G1343gat));
  AOI21_X1  g640(.A(new_n552_), .B1(new_n799_), .B2(KEYINPUT118), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n842_), .A2(new_n807_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n342_), .A2(new_n368_), .A3(new_n379_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n285_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT123), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT123), .ZN(new_n847_));
  INV_X1    g646(.A(new_n845_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n815_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n846_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n534_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n484_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g653(.A(KEYINPUT61), .B(G155gat), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT124), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n850_), .B2(new_n552_), .ZN(new_n858_));
  AOI211_X1 g657(.A(KEYINPUT124), .B(new_n553_), .C1(new_n846_), .C2(new_n849_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n856_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n847_), .B1(new_n815_), .B2(new_n848_), .ZN(new_n861_));
  AOI211_X1 g660(.A(KEYINPUT123), .B(new_n845_), .C1(new_n808_), .C2(new_n796_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n552_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT124), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n850_), .A2(new_n857_), .A3(new_n552_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n864_), .A2(new_n865_), .A3(new_n855_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n860_), .A2(new_n866_), .ZN(G1346gat));
  AND3_X1   g666(.A1(new_n850_), .A2(G162gat), .A3(new_n645_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G162gat), .B1(new_n850_), .B2(new_n612_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT125), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT125), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n592_), .B1(new_n846_), .B2(new_n849_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(G162gat), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n868_), .B1(new_n870_), .B2(new_n873_), .ZN(G1347gat));
  AND2_X1   g673(.A1(new_n801_), .A2(new_n342_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n620_), .A2(new_n381_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(new_n534_), .A3(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT62), .B1(new_n878_), .B2(KEYINPUT22), .ZN(new_n879_));
  OAI21_X1  g678(.A(G169gat), .B1(new_n878_), .B2(KEYINPUT62), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n217_), .B2(new_n879_), .ZN(G1348gat));
  AND2_X1   g681(.A1(new_n875_), .A2(new_n877_), .ZN(new_n883_));
  AOI21_X1  g682(.A(G176gat), .B1(new_n883_), .B2(new_n484_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n843_), .A2(new_n609_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n876_), .A2(new_n218_), .A3(new_n686_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n885_), .B2(new_n886_), .ZN(G1349gat));
  NOR2_X1   g686(.A1(new_n876_), .A2(new_n553_), .ZN(new_n888_));
  AOI21_X1  g687(.A(G183gat), .B1(new_n885_), .B2(new_n888_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n876_), .A2(new_n223_), .A3(new_n553_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n875_), .B2(new_n890_), .ZN(G1350gat));
  NAND3_X1  g690(.A1(new_n883_), .A2(new_n224_), .A3(new_n612_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n875_), .A2(new_n645_), .A3(new_n877_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT126), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n893_), .A2(new_n894_), .A3(G190gat), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n893_), .B2(G190gat), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n892_), .B1(new_n895_), .B2(new_n896_), .ZN(G1351gat));
  NAND3_X1  g696(.A1(new_n620_), .A2(new_n399_), .A3(new_n380_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n843_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n534_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n484_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g702(.A1(new_n843_), .A2(new_n553_), .A3(new_n898_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  AND2_X1   g704(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n904_), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n907_), .B1(new_n904_), .B2(new_n905_), .ZN(G1354gat));
  AOI21_X1  g707(.A(G218gat), .B1(new_n899_), .B2(new_n612_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n645_), .A2(G218gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT127), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n899_), .B2(new_n911_), .ZN(G1355gat));
endmodule


