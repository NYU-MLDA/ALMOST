//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n582_, new_n583_, new_n584_, new_n585_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n785_, new_n786_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n805_,
    new_n806_, new_n808_, new_n809_, new_n810_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n827_,
    new_n828_, new_n829_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_;
  XOR2_X1   g000(.A(G64gat), .B(G92gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT19), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G211gat), .B(G218gat), .Z(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G197gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(new_n213_), .A2(G204gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(G204gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT21), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  OR3_X1    g015(.A1(new_n213_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n214_), .A2(KEYINPUT91), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n217_), .B1(new_n218_), .B2(new_n215_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n212_), .B(new_n216_), .C1(new_n219_), .C2(KEYINPUT21), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(KEYINPUT21), .A3(new_n211_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT23), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n224_), .B1(G183gat), .B2(G190gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G169gat), .A2(G176gat), .ZN(new_n226_));
  INV_X1    g025(.A(G169gat), .ZN(new_n227_));
  OR3_X1    g026(.A1(new_n227_), .A2(KEYINPUT84), .A3(KEYINPUT22), .ZN(new_n228_));
  INV_X1    g027(.A(G176gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT22), .B1(new_n227_), .B2(KEYINPUT84), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n225_), .A2(new_n226_), .A3(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT25), .B(G183gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT26), .B(G190gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n227_), .A2(new_n229_), .ZN(new_n236_));
  OR2_X1    g035(.A1(new_n236_), .A2(KEYINPUT24), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(KEYINPUT24), .A3(new_n226_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n235_), .A2(new_n224_), .A3(new_n237_), .A4(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n232_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n222_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT95), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n222_), .A2(KEYINPUT95), .A3(new_n240_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(KEYINPUT22), .B(G169gat), .Z(new_n246_));
  OAI211_X1 g045(.A(new_n225_), .B(new_n226_), .C1(G176gat), .C2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n239_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n222_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT20), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n210_), .B1(new_n245_), .B2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n250_), .B1(new_n222_), .B2(new_n248_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n240_), .B2(new_n222_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n254_), .A2(new_n209_), .ZN(new_n255_));
  OAI211_X1 g054(.A(KEYINPUT32), .B(new_n207_), .C1(new_n252_), .C2(new_n255_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n251_), .A2(new_n243_), .A3(new_n210_), .A4(new_n244_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n254_), .A2(new_n209_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n207_), .A2(KEYINPUT32), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n257_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G1gat), .B(G29gat), .ZN(new_n261_));
  INV_X1    g060(.A(G85gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n261_), .B(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT0), .B(G57gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G225gat), .A2(G233gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G155gat), .B(G162gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT89), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G141gat), .A2(G148gat), .ZN(new_n272_));
  AND2_X1   g071(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n273_));
  NOR2_X1   g072(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n272_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT87), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT87), .ZN(new_n277_));
  OAI211_X1 g076(.A(new_n277_), .B(new_n272_), .C1(new_n273_), .C2(new_n274_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n271_), .B1(new_n276_), .B2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT88), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n268_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n268_), .A2(KEYINPUT2), .ZN(new_n283_));
  AND2_X1   g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n272_), .B1(new_n284_), .B2(KEYINPUT1), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n285_), .B1(new_n268_), .B2(KEYINPUT1), .ZN(new_n286_));
  AOI22_X1  g085(.A1(new_n283_), .A2(new_n286_), .B1(G141gat), .B2(G148gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n282_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G113gat), .B(G120gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(G134gat), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT85), .B(G127gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n290_), .B(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n290_), .B(new_n291_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n295_), .B1(new_n282_), .B2(new_n287_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n294_), .A2(KEYINPUT97), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT97), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n288_), .A2(new_n298_), .A3(new_n293_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n267_), .B1(new_n297_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT98), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n299_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT4), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n296_), .A2(KEYINPUT4), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n267_), .A3(new_n305_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n265_), .B1(new_n302_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n303_), .A2(new_n266_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n301_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n300_), .A2(KEYINPUT98), .ZN(new_n310_));
  NAND4_X1  g109(.A1(new_n306_), .A2(new_n309_), .A3(new_n265_), .A4(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n256_), .B(new_n260_), .C1(new_n307_), .C2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n257_), .A2(new_n258_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n206_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n257_), .A2(new_n258_), .A3(new_n207_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n304_), .A2(new_n266_), .A3(new_n305_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n265_), .B1(new_n303_), .B2(new_n267_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n317_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT33), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n311_), .A2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n302_), .A2(KEYINPUT33), .A3(new_n265_), .A4(new_n306_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n320_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n313_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G227gat), .A2(G233gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n326_), .B(KEYINPUT31), .Z(new_n327_));
  XNOR2_X1  g126(.A(new_n295_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(new_n240_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G71gat), .B(G99gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n330_), .B(G43gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT30), .B(G15gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n329_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT29), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n222_), .B1(new_n288_), .B2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(G228gat), .A3(G233gat), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n337_), .A2(KEYINPUT93), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(KEYINPUT93), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G228gat), .A2(G233gat), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n340_), .B(new_n222_), .C1(new_n288_), .C2(new_n335_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n341_), .A2(KEYINPUT92), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(KEYINPUT92), .ZN(new_n343_));
  AOI22_X1  g142(.A1(new_n338_), .A2(new_n339_), .B1(new_n342_), .B2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G78gat), .B(G106gat), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(G22gat), .B(G50gat), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n288_), .A2(new_n335_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n350_), .B1(new_n288_), .B2(new_n335_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n348_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n353_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(new_n347_), .A3(new_n351_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n346_), .B1(new_n357_), .B2(KEYINPUT94), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n345_), .B1(new_n354_), .B2(new_n356_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n344_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n344_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n334_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n325_), .A2(new_n364_), .ZN(new_n365_));
  OR3_X1    g164(.A1(new_n344_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n334_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n360_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n206_), .B1(new_n252_), .B2(new_n255_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(KEYINPUT27), .A3(new_n316_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT99), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n369_), .A2(KEYINPUT99), .A3(KEYINPUT27), .A4(new_n316_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT27), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n317_), .A2(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n372_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n307_), .A2(new_n312_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n368_), .A2(new_n376_), .A3(new_n363_), .A4(new_n377_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n365_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G230gat), .A2(G233gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT8), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT7), .ZN(new_n382_));
  INV_X1    g181(.A(G99gat), .ZN(new_n383_));
  INV_X1    g182(.A(G106gat), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G99gat), .A2(G106gat), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n385_), .A2(new_n388_), .A3(new_n389_), .A4(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G85gat), .B(G92gat), .Z(new_n392_));
  AOI21_X1  g191(.A(new_n381_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n385_), .A2(new_n390_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n397_));
  NOR3_X1   g196(.A1(new_n396_), .A2(new_n397_), .A3(KEYINPUT65), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT65), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n399_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n395_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT66), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT8), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n392_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT65), .B1(new_n396_), .B2(new_n397_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n388_), .A2(new_n399_), .A3(new_n389_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n394_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n407_), .B2(KEYINPUT66), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n393_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT64), .ZN(new_n410_));
  INV_X1    g209(.A(G92gat), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n410_), .B1(new_n262_), .B2(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(new_n412_), .A2(KEYINPUT9), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(KEYINPUT9), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n413_), .B(new_n414_), .C1(G85gat), .C2(G92gat), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n405_), .A2(new_n406_), .ZN(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT10), .B(G99gat), .Z(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(new_n384_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT67), .B1(new_n409_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n393_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n416_), .A2(KEYINPUT66), .A3(new_n395_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n392_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n381_), .B1(new_n407_), .B2(KEYINPUT66), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n422_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT67), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n419_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n421_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G71gat), .B(G78gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G57gat), .B(G64gat), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n431_), .A2(KEYINPUT11), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(KEYINPUT11), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n430_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n433_), .A2(new_n430_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n429_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n436_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n421_), .A2(new_n438_), .A3(new_n428_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n380_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT12), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  AOI211_X1 g241(.A(new_n441_), .B(new_n436_), .C1(new_n426_), .C2(new_n419_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n442_), .A2(new_n437_), .A3(new_n380_), .A4(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(KEYINPUT68), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n443_), .B1(new_n429_), .B2(new_n436_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT68), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(new_n442_), .A4(new_n380_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n440_), .B1(new_n446_), .B2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT5), .B(G176gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(G204gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G120gat), .B(G148gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n450_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(KEYINPUT69), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n455_), .B1(new_n450_), .B2(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT13), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  XOR2_X1   g258(.A(G15gat), .B(G22gat), .Z(new_n460_));
  XOR2_X1   g259(.A(KEYINPUT76), .B(G1gat), .Z(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(G8gat), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n460_), .B1(new_n462_), .B2(KEYINPUT14), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G1gat), .B(G8gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G29gat), .B(G36gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G43gat), .B(G50gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n468_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n466_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n465_), .B(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G229gat), .A2(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n473_), .A2(KEYINPUT80), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n475_), .ZN(new_n477_));
  XOR2_X1   g276(.A(new_n463_), .B(new_n464_), .Z(new_n478_));
  AND3_X1   g277(.A1(new_n469_), .A2(new_n471_), .A3(KEYINPUT15), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT15), .B1(new_n469_), .B2(new_n471_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n478_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n465_), .A2(new_n472_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT80), .B1(new_n485_), .B2(new_n475_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n476_), .B1(new_n477_), .B2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G113gat), .B(G141gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT82), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G169gat), .B(G197gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT81), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n487_), .B(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(new_n493_), .B(KEYINPUT83), .Z(new_n494_));
  NOR3_X1   g293(.A1(new_n379_), .A2(new_n459_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT71), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT70), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n426_), .A2(new_n419_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n497_), .B1(new_n498_), .B2(new_n482_), .ZN(new_n499_));
  AOI211_X1 g298(.A(KEYINPUT70), .B(new_n481_), .C1(new_n426_), .C2(new_n419_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n496_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n409_), .A2(new_n420_), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT70), .B1(new_n502_), .B2(new_n481_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n498_), .A2(new_n497_), .A3(new_n482_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(KEYINPUT71), .A3(new_n504_), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT72), .B1(new_n429_), .B2(new_n472_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT72), .ZN(new_n507_));
  INV_X1    g306(.A(new_n472_), .ZN(new_n508_));
  AOI211_X1 g307(.A(new_n507_), .B(new_n508_), .C1(new_n421_), .C2(new_n428_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n501_), .B(new_n505_), .C1(new_n506_), .C2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G232gat), .A2(G233gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT34), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n512_), .A2(KEYINPUT35), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n512_), .A2(KEYINPUT35), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  OAI221_X1 g315(.A(new_n516_), .B1(new_n499_), .B2(new_n500_), .C1(new_n506_), .C2(new_n509_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G190gat), .B(G218gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G134gat), .B(G162gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n519_), .B(new_n520_), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT36), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n521_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n524_), .A2(KEYINPUT36), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n514_), .A2(new_n525_), .A3(new_n517_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n523_), .A2(KEYINPUT73), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT73), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n514_), .A2(new_n528_), .A3(new_n525_), .A4(new_n517_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n529_), .A2(KEYINPUT37), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT74), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT37), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n518_), .A2(KEYINPUT75), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n522_), .B1(new_n518_), .B2(KEYINPUT75), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n533_), .B(new_n526_), .C1(new_n534_), .C2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT74), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n527_), .A2(new_n530_), .A3(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n532_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G231gat), .A2(G233gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(new_n540_), .B(KEYINPUT77), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n465_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(new_n438_), .ZN(new_n543_));
  XOR2_X1   g342(.A(G127gat), .B(G155gat), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(G211gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(KEYINPUT16), .B(G183gat), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n547_), .A2(KEYINPUT17), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(KEYINPUT17), .ZN(new_n549_));
  AND3_X1   g348(.A1(new_n543_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT78), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT78), .B1(new_n543_), .B2(new_n549_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n552_), .B1(new_n553_), .B2(new_n550_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT79), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n539_), .A2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n495_), .A2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n377_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n461_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n561_), .B(KEYINPUT38), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n526_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n379_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n493_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n459_), .A2(new_n566_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n565_), .A2(new_n567_), .A3(new_n555_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(new_n559_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(G1gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n562_), .A2(new_n570_), .ZN(G1324gat));
  INV_X1    g370(.A(G8gat), .ZN(new_n572_));
  INV_X1    g371(.A(new_n376_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(new_n568_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT39), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n574_), .B1(KEYINPUT100), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(KEYINPUT100), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n558_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g380(.A(G15gat), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(new_n568_), .B2(new_n367_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT41), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n558_), .A2(new_n582_), .A3(new_n367_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(G1326gat));
  INV_X1    g385(.A(G22gat), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n361_), .A2(new_n362_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n587_), .B1(new_n568_), .B2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT101), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT42), .Z(new_n591_));
  NAND3_X1  g390(.A1(new_n558_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(G1327gat));
  NAND2_X1  g392(.A1(new_n556_), .A2(new_n564_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n495_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(G29gat), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n597_), .A3(new_n559_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT43), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n365_), .A2(new_n378_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n539_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n532_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n602_));
  OAI21_X1  g401(.A(KEYINPUT43), .B1(new_n379_), .B2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n555_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n567_), .ZN(new_n605_));
  XOR2_X1   g404(.A(KEYINPUT102), .B(KEYINPUT44), .Z(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(new_n604_), .B(new_n567_), .C1(KEYINPUT102), .C2(KEYINPUT44), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(new_n559_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n598_), .B1(new_n613_), .B2(new_n597_), .ZN(G1328gat));
  OAI21_X1  g413(.A(KEYINPUT103), .B1(new_n610_), .B2(new_n376_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT103), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n608_), .A2(new_n616_), .A3(new_n609_), .A4(new_n573_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n615_), .A2(G36gat), .A3(new_n617_), .ZN(new_n618_));
  OR2_X1    g417(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n619_));
  INV_X1    g418(.A(G36gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n596_), .A2(new_n620_), .A3(new_n573_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT45), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n618_), .A2(new_n619_), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT104), .ZN(new_n624_));
  OAI21_X1  g423(.A(KEYINPUT105), .B1(new_n624_), .B2(KEYINPUT46), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n623_), .B(new_n625_), .ZN(G1329gat));
  OAI21_X1  g425(.A(G43gat), .B1(new_n610_), .B2(new_n334_), .ZN(new_n627_));
  INV_X1    g426(.A(G43gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n596_), .A2(new_n628_), .A3(new_n367_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n630_), .B(new_n631_), .Z(G1330gat));
  NAND2_X1  g431(.A1(new_n611_), .A2(new_n588_), .ZN(new_n633_));
  OR2_X1    g432(.A1(new_n633_), .A2(KEYINPUT107), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(KEYINPUT107), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(G50gat), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(G50gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n596_), .A2(new_n637_), .A3(new_n588_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(G1331gat));
  NOR3_X1   g438(.A1(new_n379_), .A2(new_n493_), .A3(new_n458_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n640_), .A2(new_n557_), .ZN(new_n641_));
  AOI21_X1  g440(.A(G57gat), .B1(new_n641_), .B2(new_n559_), .ZN(new_n642_));
  AND4_X1   g441(.A1(new_n555_), .A2(new_n565_), .A3(new_n459_), .A4(new_n494_), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n643_), .A2(new_n559_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n642_), .B1(new_n644_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g444(.A(G64gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n643_), .B2(new_n573_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT48), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n641_), .A2(new_n646_), .A3(new_n573_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(G1333gat));
  INV_X1    g449(.A(G71gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n643_), .B2(new_n367_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT49), .Z(new_n653_));
  NAND3_X1  g452(.A1(new_n641_), .A2(new_n651_), .A3(new_n367_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1334gat));
  INV_X1    g454(.A(G78gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n643_), .B2(new_n588_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT108), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT50), .Z(new_n659_));
  NAND3_X1  g458(.A1(new_n641_), .A2(new_n656_), .A3(new_n588_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1335gat));
  AND2_X1   g460(.A1(new_n640_), .A2(new_n595_), .ZN(new_n662_));
  AOI21_X1  g461(.A(G85gat), .B1(new_n662_), .B2(new_n559_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n458_), .A2(new_n493_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n604_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT109), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n604_), .A2(KEYINPUT109), .A3(new_n664_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n559_), .A2(G85gat), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT110), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n663_), .B1(new_n669_), .B2(new_n671_), .ZN(G1336gat));
  AOI21_X1  g471(.A(G92gat), .B1(new_n662_), .B2(new_n573_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n376_), .A2(new_n411_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n669_), .B2(new_n674_), .ZN(G1337gat));
  NAND3_X1  g474(.A1(new_n667_), .A2(new_n367_), .A3(new_n668_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(G99gat), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT51), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n662_), .A2(new_n417_), .A3(new_n367_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT112), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT111), .B1(new_n677_), .B2(new_n679_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT111), .ZN(new_n684_));
  INV_X1    g483(.A(new_n679_), .ZN(new_n685_));
  AOI211_X1 g484(.A(new_n684_), .B(new_n685_), .C1(new_n676_), .C2(G99gat), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n683_), .A2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n682_), .B1(new_n687_), .B2(KEYINPUT51), .ZN(new_n688_));
  NOR4_X1   g487(.A1(new_n683_), .A2(new_n686_), .A3(new_n681_), .A4(new_n678_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1338gat));
  INV_X1    g489(.A(new_n588_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G106gat), .B1(new_n665_), .B2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT52), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n662_), .A2(new_n384_), .A3(new_n588_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g495(.A(new_n455_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n566_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n446_), .A2(new_n449_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT55), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n447_), .A2(KEYINPUT55), .A3(new_n442_), .A4(new_n380_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT116), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n447_), .A2(new_n442_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT115), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT115), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n447_), .A2(new_n707_), .A3(new_n442_), .ZN(new_n708_));
  NAND4_X1  g507(.A1(new_n706_), .A2(G230gat), .A3(G233gat), .A4(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n701_), .A2(new_n704_), .A3(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n456_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(KEYINPUT56), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT56), .B1(new_n710_), .B2(new_n711_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n698_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(KEYINPUT117), .ZN(new_n715_));
  INV_X1    g514(.A(new_n491_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n487_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n485_), .B(KEYINPUT118), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(new_n474_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT119), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n720_), .A2(new_n721_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n717_), .B1(new_n722_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n457_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT117), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n698_), .B(new_n727_), .C1(new_n712_), .C2(new_n713_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n715_), .A2(new_n726_), .A3(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n563_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT57), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n729_), .A2(KEYINPUT57), .A3(new_n563_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT121), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n710_), .A2(new_n711_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT56), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n710_), .A2(KEYINPUT56), .A3(new_n711_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n724_), .A2(new_n697_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n736_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n734_), .B1(new_n743_), .B2(new_n602_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n742_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n735_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n539_), .A2(new_n746_), .A3(KEYINPUT121), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n741_), .A2(KEYINPUT58), .A3(new_n742_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n744_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n732_), .A2(new_n733_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n556_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n602_), .A2(new_n555_), .A3(new_n458_), .A4(new_n494_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n752_), .A2(KEYINPUT114), .A3(KEYINPUT54), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT114), .B1(new_n752_), .B2(KEYINPUT54), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT113), .B1(new_n752_), .B2(KEYINPUT54), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n602_), .A2(new_n555_), .A3(new_n494_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT113), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .A4(new_n458_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n755_), .A2(new_n756_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n751_), .A2(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n573_), .A2(new_n377_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n367_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n762_), .A2(new_n691_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(G113gat), .B1(new_n767_), .B2(new_n493_), .ZN(new_n768_));
  XOR2_X1   g567(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n769_));
  NAND4_X1  g568(.A1(new_n762_), .A2(new_n691_), .A3(new_n765_), .A4(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(KEYINPUT123), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n766_), .A2(KEYINPUT59), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n588_), .B1(new_n751_), .B2(new_n761_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT123), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(new_n765_), .A4(new_n769_), .ZN(new_n775_));
  AND4_X1   g574(.A1(G113gat), .A2(new_n771_), .A3(new_n772_), .A4(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n494_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n768_), .B1(new_n776_), .B2(new_n777_), .ZN(G1340gat));
  NAND4_X1  g577(.A1(new_n771_), .A2(new_n772_), .A3(new_n459_), .A4(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(G120gat), .ZN(new_n780_));
  INV_X1    g579(.A(G120gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n458_), .B2(KEYINPUT60), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n767_), .B(new_n782_), .C1(KEYINPUT60), .C2(new_n781_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n780_), .A2(new_n783_), .ZN(G1341gat));
  AOI21_X1  g583(.A(G127gat), .B1(new_n767_), .B2(new_n555_), .ZN(new_n785_));
  AND4_X1   g584(.A1(new_n555_), .A2(new_n771_), .A3(new_n772_), .A4(new_n775_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n786_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g586(.A(G134gat), .B1(new_n767_), .B2(new_n564_), .ZN(new_n788_));
  AND4_X1   g587(.A1(G134gat), .A2(new_n771_), .A3(new_n772_), .A4(new_n775_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n789_), .B2(new_n539_), .ZN(G1343gat));
  AND2_X1   g589(.A1(new_n760_), .A2(new_n756_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n556_), .A2(new_n750_), .B1(new_n791_), .B2(new_n755_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n792_), .A2(new_n367_), .A3(new_n691_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(new_n763_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n493_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(G141gat), .ZN(new_n796_));
  INV_X1    g595(.A(G141gat), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n794_), .A2(new_n797_), .A3(new_n493_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n796_), .A2(new_n798_), .ZN(G1344gat));
  NAND2_X1  g598(.A1(new_n794_), .A2(new_n459_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(G148gat), .ZN(new_n801_));
  INV_X1    g600(.A(G148gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n794_), .A2(new_n802_), .A3(new_n459_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1345gat));
  NAND3_X1  g603(.A1(new_n793_), .A2(new_n555_), .A3(new_n763_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(KEYINPUT61), .B(G155gat), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1346gat));
  NAND2_X1  g606(.A1(new_n794_), .A2(new_n564_), .ZN(new_n808_));
  INV_X1    g607(.A(G162gat), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n602_), .A2(new_n809_), .ZN(new_n810_));
  AOI22_X1  g609(.A1(new_n808_), .A2(new_n809_), .B1(new_n794_), .B2(new_n810_), .ZN(G1347gat));
  NOR2_X1   g610(.A1(new_n559_), .A2(new_n376_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n773_), .A2(new_n367_), .A3(new_n493_), .A4(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT62), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n813_), .A2(new_n814_), .A3(G169gat), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n814_), .B1(new_n813_), .B2(G169gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n773_), .A2(new_n367_), .A3(new_n812_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n566_), .A2(new_n246_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT124), .ZN(new_n819_));
  OAI22_X1  g618(.A1(new_n815_), .A2(new_n816_), .B1(new_n817_), .B2(new_n819_), .ZN(G1348gat));
  OAI22_X1  g619(.A1(new_n817_), .A2(new_n458_), .B1(KEYINPUT125), .B2(new_n229_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n812_), .ZN(new_n822_));
  NOR4_X1   g621(.A1(new_n792_), .A2(new_n334_), .A3(new_n588_), .A4(new_n822_), .ZN(new_n823_));
  XOR2_X1   g622(.A(KEYINPUT125), .B(G176gat), .Z(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n459_), .A3(new_n824_), .ZN(new_n825_));
  AND2_X1   g624(.A1(new_n821_), .A2(new_n825_), .ZN(G1349gat));
  NAND2_X1  g625(.A1(new_n823_), .A2(new_n555_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(G183gat), .ZN(new_n828_));
  INV_X1    g627(.A(new_n233_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(new_n827_), .ZN(G1350gat));
  INV_X1    g629(.A(G190gat), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n831_), .B1(new_n823_), .B2(new_n539_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n234_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n817_), .A2(new_n563_), .A3(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT126), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n823_), .A2(new_n564_), .A3(new_n234_), .ZN(new_n836_));
  OAI21_X1  g635(.A(G190gat), .B1(new_n817_), .B2(new_n602_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT126), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n836_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n835_), .A2(new_n839_), .ZN(G1351gat));
  NAND3_X1  g639(.A1(new_n793_), .A2(new_n493_), .A3(new_n812_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT127), .B1(new_n841_), .B2(new_n213_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n213_), .ZN(new_n843_));
  NOR4_X1   g642(.A1(new_n792_), .A2(new_n367_), .A3(new_n691_), .A4(new_n822_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT127), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(G197gat), .A4(new_n493_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n842_), .A2(new_n843_), .A3(new_n846_), .ZN(G1352gat));
  NAND2_X1  g646(.A1(new_n844_), .A2(new_n459_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g648(.A(KEYINPUT63), .B(G211gat), .C1(new_n844_), .C2(new_n555_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n844_), .A2(new_n555_), .ZN(new_n851_));
  XOR2_X1   g650(.A(KEYINPUT63), .B(G211gat), .Z(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(G1354gat));
  AOI21_X1  g652(.A(G218gat), .B1(new_n844_), .B2(new_n564_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n539_), .A2(G218gat), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n844_), .B2(new_n855_), .ZN(G1355gat));
endmodule


