//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n933_, new_n934_,
    new_n935_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203_));
  INV_X1    g002(.A(G8gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G1gat), .B(G8gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(new_n206_), .B(new_n207_), .Z(new_n208_));
  NAND2_X1  g007(.A1(G231gat), .A2(G233gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G71gat), .B(G78gat), .Z(new_n211_));
  XNOR2_X1  g010(.A(G57gat), .B(G64gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n211_), .B1(KEYINPUT11), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(KEYINPUT11), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n210_), .B(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G127gat), .B(G155gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT16), .ZN(new_n219_));
  INV_X1    g018(.A(G183gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(G211gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n222_), .A2(new_n223_), .ZN(new_n225_));
  OR3_X1    g024(.A1(new_n217_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n217_), .A2(new_n225_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(KEYINPUT89), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G141gat), .A2(G148gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT3), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G141gat), .A2(G148gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(KEYINPUT85), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n230_), .B(new_n232_), .C1(KEYINPUT2), .C2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G155gat), .A2(G162gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT86), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n235_), .B(new_n238_), .C1(G155gat), .C2(G162gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT90), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n234_), .A2(new_n231_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n236_), .B(KEYINPUT86), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n243_));
  OAI22_X1  g042(.A1(new_n242_), .A2(new_n243_), .B1(G155gat), .B2(G162gat), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT87), .ZN(new_n245_));
  OAI22_X1  g044(.A1(new_n244_), .A2(new_n245_), .B1(KEYINPUT1), .B2(new_n238_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  OAI211_X1 g046(.A(KEYINPUT88), .B(new_n241_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n241_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT88), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n240_), .A2(new_n248_), .A3(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G127gat), .B(G134gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G113gat), .B(G120gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n253_), .B(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n255_), .B(KEYINPUT84), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT4), .B1(new_n252_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n252_), .A2(new_n256_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n239_), .A2(KEYINPUT90), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n239_), .A2(KEYINPUT90), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n259_), .A2(new_n260_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n261_), .A2(new_n255_), .A3(new_n248_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n258_), .A2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n257_), .B1(new_n263_), .B2(KEYINPUT4), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G225gat), .A2(G233gat), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G1gat), .B(G29gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT0), .ZN(new_n269_));
  INV_X1    g068(.A(G57gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(G85gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n263_), .A2(new_n265_), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n267_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n273_), .B1(new_n267_), .B2(new_n274_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G64gat), .B(G92gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G8gat), .B(G36gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT100), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n280_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT19), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G211gat), .B(G218gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(KEYINPUT92), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT21), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G197gat), .B(G204gat), .Z(new_n291_));
  OAI21_X1  g090(.A(new_n291_), .B1(KEYINPUT21), .B2(new_n287_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n290_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT93), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OR3_X1    g097(.A1(new_n296_), .A2(KEYINPUT82), .A3(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT82), .B1(new_n296_), .B2(new_n298_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n299_), .B(new_n300_), .C1(KEYINPUT23), .C2(new_n297_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT80), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT24), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT25), .B(G183gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT26), .B(G190gat), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n303_), .A2(new_n304_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT24), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n301_), .B(new_n307_), .C1(new_n303_), .C2(new_n309_), .ZN(new_n310_));
  MUX2_X1   g109(.A(KEYINPUT23), .B(new_n296_), .S(new_n298_), .Z(new_n311_));
  OAI21_X1  g110(.A(new_n311_), .B1(G183gat), .B2(G190gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT22), .B(G169gat), .ZN(new_n313_));
  INV_X1    g112(.A(G176gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n308_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n310_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT93), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n293_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n295_), .A2(new_n317_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n301_), .B1(G183gat), .B2(G190gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n315_), .A2(new_n308_), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n323_), .B(KEYINPUT97), .Z(new_n324_));
  AND2_X1   g123(.A1(new_n307_), .A2(new_n311_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n303_), .B1(KEYINPUT96), .B2(new_n309_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(KEYINPUT96), .B2(new_n309_), .ZN(new_n327_));
  AOI22_X1  g126(.A1(new_n322_), .A2(new_n324_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT103), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n294_), .B1(new_n328_), .B2(KEYINPUT103), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT20), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n321_), .B1(new_n332_), .B2(KEYINPUT104), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT104), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n334_), .B(KEYINPUT20), .C1(new_n330_), .C2(new_n331_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n286_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  OR2_X1    g135(.A1(new_n328_), .A2(new_n294_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n293_), .B(new_n318_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n317_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n337_), .A2(new_n340_), .A3(KEYINPUT20), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n341_), .A2(new_n285_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n283_), .B1(new_n336_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n285_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n286_), .A2(KEYINPUT20), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT98), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n328_), .A2(new_n346_), .A3(new_n294_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n346_), .B1(new_n328_), .B2(new_n294_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n320_), .B(new_n345_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n283_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n344_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n351_), .A2(KEYINPUT27), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n343_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT27), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n350_), .B1(new_n344_), .B2(new_n349_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT101), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n351_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  AOI211_X1 g156(.A(KEYINPUT101), .B(new_n350_), .C1(new_n344_), .C2(new_n349_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n354_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n277_), .A2(new_n353_), .A3(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G15gat), .B(G43gat), .ZN(new_n361_));
  INV_X1    g160(.A(G227gat), .ZN(new_n362_));
  INV_X1    g161(.A(G233gat), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n310_), .A2(KEYINPUT30), .A3(new_n316_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT30), .B1(new_n310_), .B2(new_n316_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n364_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT30), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n317_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n364_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n365_), .A3(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G71gat), .B(G99gat), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n368_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(new_n368_), .B2(new_n372_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n361_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n256_), .B(KEYINPUT31), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT83), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n368_), .A2(new_n372_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n373_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n361_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n383_), .A3(new_n374_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n377_), .A2(new_n379_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n379_), .B1(new_n377_), .B2(new_n384_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G78gat), .B(G106gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n390_), .A2(KEYINPUT94), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(new_n252_), .B2(KEYINPUT29), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G22gat), .B(G50gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396_));
  INV_X1    g195(.A(new_n392_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n261_), .A2(new_n396_), .A3(new_n248_), .A4(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n393_), .A2(new_n395_), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n395_), .B1(new_n393_), .B2(new_n398_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n391_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n401_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n403_), .A2(new_n390_), .A3(new_n399_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT95), .ZN(new_n406_));
  INV_X1    g205(.A(G228gat), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n407_), .A2(new_n363_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n252_), .A2(KEYINPUT29), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n410_), .B2(new_n293_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n338_), .A2(new_n408_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n406_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n414_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n416_), .A2(new_n411_), .A3(KEYINPUT95), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n405_), .A2(new_n418_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n402_), .B(new_n404_), .C1(new_n415_), .C2(new_n417_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n388_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n387_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n419_), .A2(new_n420_), .B1(new_n385_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n360_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT102), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n425_), .A2(KEYINPUT33), .ZN(new_n426_));
  INV_X1    g225(.A(new_n274_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n427_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(new_n428_), .B2(new_n273_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n357_), .A2(new_n358_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n267_), .A2(new_n274_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n273_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n426_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n263_), .A2(new_n265_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n435_), .A2(new_n432_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n436_), .B1(new_n266_), .B2(new_n264_), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n429_), .A2(new_n430_), .A3(new_n434_), .A4(new_n437_), .ZN(new_n438_));
  OAI211_X1 g237(.A(KEYINPUT32), .B(new_n350_), .C1(new_n336_), .C2(new_n342_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n350_), .A2(KEYINPUT32), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n344_), .A2(new_n349_), .A3(new_n440_), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n439_), .B(new_n441_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n438_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n422_), .A2(new_n385_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n444_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n228_), .B1(new_n424_), .B2(new_n446_), .ZN(new_n447_));
  XOR2_X1   g246(.A(KEYINPUT10), .B(G99gat), .Z(new_n448_));
  INV_X1    g247(.A(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(G92gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n272_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G85gat), .A2(G92gat), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(KEYINPUT9), .A3(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n453_), .A2(KEYINPUT9), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n450_), .A2(new_n454_), .A3(new_n455_), .A4(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT66), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT65), .ZN(new_n463_));
  AND2_X1   g262(.A1(G85gat), .A2(G92gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(G85gat), .A2(G92gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n452_), .A2(KEYINPUT65), .A3(new_n453_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT8), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT64), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT64), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT8), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n466_), .A2(new_n467_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT7), .ZN(new_n474_));
  INV_X1    g273(.A(G99gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n449_), .ZN(new_n476_));
  OAI21_X1  g275(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n477_));
  AND4_X1   g276(.A1(new_n458_), .A2(new_n476_), .A3(new_n459_), .A4(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n462_), .B1(new_n473_), .B2(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n466_), .A2(new_n467_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n476_), .A2(new_n458_), .A3(new_n459_), .A4(new_n477_), .ZN(new_n481_));
  NAND4_X1  g280(.A1(new_n480_), .A2(KEYINPUT66), .A3(new_n481_), .A4(new_n472_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n477_), .ZN(new_n483_));
  NOR3_X1   g282(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT67), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n476_), .A2(new_n486_), .A3(new_n477_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n460_), .A3(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n468_), .B1(new_n488_), .B2(new_n480_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT68), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n479_), .B(new_n482_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n466_), .A2(new_n467_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n458_), .A2(new_n459_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n476_), .A2(new_n477_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n494_), .B2(KEYINPUT67), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n492_), .B1(new_n495_), .B2(new_n487_), .ZN(new_n496_));
  NOR3_X1   g295(.A1(new_n496_), .A2(KEYINPUT68), .A3(new_n468_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n461_), .B1(new_n491_), .B2(new_n497_), .ZN(new_n498_));
  XOR2_X1   g297(.A(G29gat), .B(G36gat), .Z(new_n499_));
  XOR2_X1   g298(.A(G43gat), .B(G50gat), .Z(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT15), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n498_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT72), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G232gat), .A2(G233gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT34), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT35), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n461_), .B(new_n501_), .C1(new_n491_), .C2(new_n497_), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n505_), .A2(new_n506_), .A3(new_n511_), .A4(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n512_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT68), .B1(new_n496_), .B2(new_n468_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n482_), .A2(new_n479_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n489_), .A2(new_n490_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n503_), .B1(new_n518_), .B2(new_n461_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n508_), .A2(KEYINPUT35), .ZN(new_n520_));
  NOR3_X1   g319(.A1(new_n514_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n511_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n505_), .B2(KEYINPUT72), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n513_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G190gat), .B(G218gat), .Z(new_n525_));
  XNOR2_X1  g324(.A(G134gat), .B(G162gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT36), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT73), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT74), .B1(new_n524_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n524_), .A2(KEYINPUT74), .A3(new_n530_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n524_), .A2(KEYINPUT76), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n527_), .B(KEYINPUT36), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n511_), .B1(new_n519_), .B2(new_n506_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n505_), .A2(new_n512_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n537_), .B1(new_n538_), .B2(new_n520_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT76), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n513_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n535_), .A2(new_n536_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n534_), .A2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(new_n447_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT13), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n498_), .A2(new_n215_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n216_), .B(new_n461_), .C1(new_n491_), .C2(new_n497_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n546_), .A2(KEYINPUT69), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G230gat), .A2(G233gat), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT69), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n498_), .A2(new_n551_), .A3(new_n215_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT70), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n548_), .A2(KEYINPUT70), .A3(new_n550_), .A4(new_n552_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n547_), .A2(KEYINPUT12), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n216_), .B1(new_n518_), .B2(new_n461_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n498_), .A2(new_n560_), .A3(new_n215_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n549_), .B1(new_n559_), .B2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n555_), .A2(new_n556_), .A3(new_n563_), .ZN(new_n564_));
  XOR2_X1   g363(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n565_));
  XNOR2_X1  g364(.A(G120gat), .B(G148gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(G176gat), .B(G204gat), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n567_), .B(new_n568_), .Z(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n564_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n546_), .A2(KEYINPUT12), .A3(new_n547_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n561_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n553_), .A2(new_n554_), .B1(new_n573_), .B2(new_n549_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n569_), .B1(new_n574_), .B2(new_n556_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n545_), .B1(new_n571_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n564_), .A2(new_n570_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n574_), .A2(new_n556_), .A3(new_n569_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(KEYINPUT13), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n208_), .A2(new_n501_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT78), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n208_), .A2(new_n501_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(G229gat), .A3(G233gat), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n503_), .A2(new_n208_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G229gat), .A2(G233gat), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n586_), .A2(new_n587_), .A3(new_n581_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(G169gat), .ZN(new_n590_));
  INV_X1    g389(.A(G197gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n585_), .A2(new_n588_), .A3(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n593_), .A2(KEYINPUT79), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(KEYINPUT79), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n585_), .A2(new_n588_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n592_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n580_), .A2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n544_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n277_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n202_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT37), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n524_), .A2(KEYINPUT74), .A3(new_n530_), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n542_), .B(new_n606_), .C1(new_n531_), .C2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT77), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT77), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n534_), .A2(new_n610_), .A3(new_n606_), .A4(new_n542_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n539_), .A2(new_n513_), .A3(new_n536_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT75), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n534_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT37), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n612_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n447_), .A2(new_n602_), .A3(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT105), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n619_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n277_), .A2(G1gat), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n620_), .A2(new_n621_), .A3(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT106), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT106), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n620_), .A2(new_n626_), .A3(new_n621_), .A4(new_n622_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n605_), .B1(new_n629_), .B2(KEYINPUT38), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT38), .B1(new_n624_), .B2(new_n627_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n631_), .A2(KEYINPUT107), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(KEYINPUT107), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n630_), .A2(new_n632_), .A3(new_n633_), .ZN(G1324gat));
  AND2_X1   g433(.A1(new_n353_), .A2(new_n359_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n620_), .A2(new_n204_), .A3(new_n636_), .A4(new_n621_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT39), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n447_), .A2(new_n636_), .A3(new_n602_), .A4(new_n543_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(G8gat), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n639_), .A2(new_n638_), .A3(G8gat), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n637_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT108), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT108), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n637_), .B(new_n644_), .C1(new_n640_), .C2(new_n641_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n643_), .A2(KEYINPUT40), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT40), .B1(new_n643_), .B2(new_n645_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1325gat));
  INV_X1    g447(.A(G15gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n649_), .B1(new_n603_), .B2(new_n444_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT41), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n620_), .A2(new_n621_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n649_), .A3(new_n444_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1326gat));
  INV_X1    g453(.A(G22gat), .ZN(new_n655_));
  INV_X1    g454(.A(new_n419_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n420_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n655_), .B1(new_n603_), .B2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(KEYINPUT109), .B(KEYINPUT42), .Z(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n652_), .A2(new_n655_), .A3(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1327gat));
  NAND2_X1  g462(.A1(new_n424_), .A2(new_n446_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n543_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n602_), .A2(new_n228_), .ZN(new_n667_));
  OR3_X1    g466(.A1(new_n666_), .A2(KEYINPUT111), .A3(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT111), .B1(new_n666_), .B2(new_n667_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(G29gat), .B1(new_n670_), .B2(new_n604_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  AOI22_X1  g471(.A1(new_n609_), .A2(new_n611_), .B1(KEYINPUT37), .B2(new_n615_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n664_), .B2(new_n673_), .ZN(new_n674_));
  AOI211_X1 g473(.A(KEYINPUT43), .B(new_n617_), .C1(new_n424_), .C2(new_n446_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n667_), .B(KEYINPUT110), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(KEYINPUT44), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n676_), .A2(KEYINPUT44), .A3(new_n677_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n681_), .A2(G29gat), .A3(new_n604_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n671_), .B1(new_n680_), .B2(new_n682_), .ZN(G1328gat));
  NAND2_X1  g482(.A1(new_n681_), .A2(new_n636_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G36gat), .B1(new_n679_), .B2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n635_), .A2(G36gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n668_), .A2(new_n669_), .A3(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT45), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT46), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n685_), .A2(new_n688_), .A3(KEYINPUT46), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1329gat));
  AND2_X1   g492(.A1(new_n670_), .A2(new_n444_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n681_), .A2(G43gat), .A3(new_n444_), .ZN(new_n695_));
  OAI22_X1  g494(.A1(new_n694_), .A2(G43gat), .B1(new_n679_), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g496(.A(G50gat), .B1(new_n670_), .B2(new_n658_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n681_), .A2(G50gat), .A3(new_n658_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n680_), .B2(new_n699_), .ZN(G1331gat));
  INV_X1    g499(.A(new_n580_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(new_n600_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n544_), .A2(new_n702_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G57gat), .B1(new_n703_), .B2(new_n277_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n600_), .B1(new_n612_), .B2(new_n616_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n447_), .A2(new_n580_), .A3(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(new_n270_), .A3(new_n604_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n707_), .ZN(G1332gat));
  INV_X1    g507(.A(G64gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n706_), .A2(new_n709_), .A3(new_n636_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n703_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n709_), .B1(new_n711_), .B2(new_n636_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n712_), .A2(new_n714_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n710_), .B1(new_n715_), .B2(new_n716_), .ZN(G1333gat));
  OAI21_X1  g516(.A(G71gat), .B1(new_n703_), .B2(new_n388_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT49), .ZN(new_n719_));
  INV_X1    g518(.A(G71gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n706_), .A2(new_n720_), .A3(new_n444_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1334gat));
  INV_X1    g521(.A(G78gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n706_), .A2(new_n723_), .A3(new_n658_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT50), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n711_), .A2(new_n658_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(G78gat), .ZN(new_n727_));
  AOI211_X1 g526(.A(KEYINPUT50), .B(new_n723_), .C1(new_n711_), .C2(new_n658_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT113), .ZN(G1335gat));
  INV_X1    g529(.A(new_n228_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n701_), .A2(new_n731_), .A3(new_n600_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n676_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G85gat), .B1(new_n734_), .B2(new_n277_), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n664_), .A2(new_n665_), .A3(new_n732_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n272_), .A3(new_n604_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1336gat));
  OAI21_X1  g537(.A(G92gat), .B1(new_n734_), .B2(new_n635_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n736_), .A2(new_n451_), .A3(new_n636_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(G1337gat));
  AND3_X1   g540(.A1(new_n736_), .A2(new_n444_), .A3(new_n448_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n733_), .A2(new_n444_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n743_), .B2(G99gat), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT51), .Z(G1338gat));
  OAI211_X1 g544(.A(new_n658_), .B(new_n732_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G106gat), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT52), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n746_), .A2(new_n749_), .A3(G106gat), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n736_), .A2(new_n449_), .A3(new_n658_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT114), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n755_));
  AND3_X1   g554(.A1(new_n746_), .A2(new_n749_), .A3(G106gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n749_), .B1(new_n746_), .B2(G106gat), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n755_), .B(new_n752_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n754_), .A2(KEYINPUT53), .A3(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT53), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n755_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n758_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n759_), .A2(new_n763_), .ZN(G1339gat));
  NOR2_X1   g563(.A1(new_n636_), .A2(new_n277_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n572_), .A2(new_n550_), .A3(new_n561_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT115), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT115), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n572_), .A2(new_n769_), .A3(new_n550_), .A4(new_n561_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n563_), .A2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n573_), .A2(KEYINPUT55), .A3(new_n549_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n569_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT118), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n768_), .A2(new_n770_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n773_), .A2(new_n774_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n570_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n776_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n777_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT55), .B1(new_n573_), .B2(new_n549_), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n772_), .B(new_n550_), .C1(new_n572_), .C2(new_n561_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n784_), .B1(new_n787_), .B2(new_n771_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n779_), .A2(new_n783_), .A3(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT119), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n792_), .A2(KEYINPUT58), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n584_), .A2(new_n587_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n598_), .ZN(new_n796_));
  OR2_X1    g595(.A1(new_n796_), .A2(KEYINPUT117), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n587_), .B1(new_n208_), .B2(new_n501_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n796_), .A2(KEYINPUT117), .B1(new_n586_), .B2(new_n798_), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n594_), .A2(new_n595_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n578_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n791_), .A2(new_n794_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(new_n673_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n794_), .B1(new_n791_), .B2(new_n802_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n577_), .A2(new_n578_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n800_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n569_), .B1(new_n787_), .B2(new_n771_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(KEYINPUT56), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n782_), .A2(KEYINPUT116), .A3(new_n776_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n778_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n600_), .A2(new_n578_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n808_), .B1(new_n813_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT57), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n665_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  OAI22_X1  g618(.A1(new_n804_), .A2(new_n805_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT56), .B1(new_n775_), .B2(new_n570_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n778_), .B1(new_n821_), .B2(KEYINPUT116), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n810_), .A2(new_n809_), .A3(KEYINPUT56), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n815_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n807_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT57), .B1(new_n825_), .B2(new_n543_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n228_), .B1(new_n820_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n576_), .A2(new_n731_), .A3(new_n579_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n705_), .B2(new_n830_), .ZN(new_n831_));
  NOR4_X1   g630(.A1(new_n673_), .A2(KEYINPUT54), .A3(new_n829_), .A4(new_n600_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n766_), .B1(new_n827_), .B2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n423_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(G113gat), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n600_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n835_), .B2(new_n423_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n817_), .B1(new_n816_), .B2(new_n665_), .ZN(new_n842_));
  AOI211_X1 g641(.A(KEYINPUT118), .B(new_n784_), .C1(new_n787_), .C2(new_n771_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n789_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n844_));
  NOR3_X1   g643(.A1(new_n821_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n793_), .B1(new_n845_), .B2(new_n801_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n673_), .A3(new_n803_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n788_), .B1(new_n783_), .B2(new_n809_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n814_), .B1(new_n848_), .B2(new_n812_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n818_), .B1(new_n849_), .B2(new_n808_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n842_), .A2(new_n847_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n833_), .B1(new_n851_), .B2(new_n228_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n423_), .ZN(new_n853_));
  NOR4_X1   g652(.A1(new_n852_), .A2(KEYINPUT59), .A3(new_n853_), .A4(new_n766_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n841_), .A2(new_n854_), .A3(new_n601_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n839_), .B1(new_n855_), .B2(new_n838_), .ZN(G1340gat));
  NOR2_X1   g655(.A1(new_n841_), .A2(new_n854_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n701_), .A2(G120gat), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n835_), .B(new_n423_), .C1(KEYINPUT60), .C2(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n857_), .A2(new_n859_), .A3(new_n580_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G120gat), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(KEYINPUT60), .B2(new_n859_), .ZN(G1341gat));
  INV_X1    g661(.A(G127gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n863_), .B1(new_n857_), .B2(new_n731_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n836_), .A2(G127gat), .A3(new_n228_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT120), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n865_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT120), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n841_), .A2(new_n854_), .A3(new_n228_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n867_), .B(new_n868_), .C1(new_n869_), .C2(new_n863_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n866_), .A2(new_n870_), .ZN(G1342gat));
  INV_X1    g670(.A(G134gat), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n837_), .A2(new_n872_), .A3(new_n665_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n841_), .A2(new_n854_), .A3(new_n617_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n873_), .B1(new_n874_), .B2(new_n872_), .ZN(G1343gat));
  NAND3_X1  g674(.A1(new_n835_), .A2(KEYINPUT121), .A3(new_n421_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(KEYINPUT121), .B1(new_n835_), .B2(new_n421_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n600_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT122), .B(G141gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1344gat));
  OAI21_X1  g680(.A(new_n580_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g682(.A(new_n731_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(KEYINPUT61), .B(G155gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1346gat));
  INV_X1    g685(.A(G162gat), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n887_), .B(new_n665_), .C1(new_n877_), .C2(new_n878_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n878_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n617_), .B1(new_n889_), .B2(new_n876_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n888_), .B1(new_n890_), .B2(new_n887_), .ZN(G1347gat));
  NAND2_X1  g690(.A1(new_n827_), .A2(new_n834_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n635_), .A2(new_n604_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n894_), .A2(new_n895_), .A3(new_n388_), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT123), .B1(new_n893_), .B2(new_n444_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n896_), .A2(new_n658_), .A3(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n892_), .A2(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(G169gat), .B1(new_n899_), .B2(new_n601_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(KEYINPUT62), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n899_), .A2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n892_), .A2(KEYINPUT124), .A3(new_n898_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n600_), .A2(new_n313_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(KEYINPUT125), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n901_), .B1(new_n905_), .B2(new_n907_), .ZN(G1348gat));
  NOR3_X1   g707(.A1(new_n899_), .A2(new_n314_), .A3(new_n701_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n905_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n580_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n911_), .B2(new_n314_), .ZN(G1349gat));
  OAI21_X1  g711(.A(new_n220_), .B1(new_n899_), .B2(new_n228_), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n228_), .A2(new_n305_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n905_), .B2(new_n914_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT126), .ZN(G1350gat));
  OAI21_X1  g715(.A(G190gat), .B1(new_n905_), .B2(new_n617_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n665_), .A2(new_n306_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n905_), .B2(new_n918_), .ZN(G1351gat));
  AND3_X1   g718(.A1(new_n892_), .A2(new_n421_), .A3(new_n893_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n920_), .A2(G197gat), .A3(new_n600_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n921_), .A2(KEYINPUT127), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n921_), .A2(KEYINPUT127), .ZN(new_n923_));
  AOI21_X1  g722(.A(G197gat), .B1(new_n920_), .B2(new_n600_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n922_), .A2(new_n923_), .A3(new_n924_), .ZN(G1352gat));
  NAND2_X1  g724(.A1(new_n920_), .A2(new_n580_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g726(.A1(new_n920_), .A2(new_n731_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  AND2_X1   g728(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n928_), .A2(new_n929_), .A3(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n931_), .B1(new_n928_), .B2(new_n929_), .ZN(G1354gat));
  INV_X1    g731(.A(G218gat), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n920_), .A2(new_n933_), .A3(new_n665_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n920_), .A2(new_n673_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n935_), .B2(new_n933_), .ZN(G1355gat));
endmodule


