//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_;
  INV_X1    g000(.A(KEYINPUT37), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G190gat), .B(G218gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  NAND2_X1  g004(.A1(G232gat), .A2(G233gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n206_), .B(KEYINPUT34), .Z(new_n207_));
  INV_X1    g006(.A(KEYINPUT35), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT79), .ZN(new_n210_));
  INV_X1    g009(.A(new_n207_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n210_), .B1(KEYINPUT35), .B2(new_n211_), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT67), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT67), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(KEYINPUT6), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(new_n215_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n217_), .B1(new_n218_), .B2(new_n213_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G92gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(G85gat), .ZN(new_n222_));
  INV_X1    g021(.A(G85gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(G92gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT9), .ZN(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT10), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n228_), .A2(G99gat), .ZN(new_n229_));
  INV_X1    g028(.A(G99gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(KEYINPUT10), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n227_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT9), .ZN(new_n234_));
  NAND2_X1  g033(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(G85gat), .A4(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n226_), .A2(new_n232_), .A3(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT7), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n238_), .A2(new_n230_), .A3(new_n227_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT8), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n220_), .B1(new_n237_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n225_), .A2(KEYINPUT8), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n214_), .A2(new_n215_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(KEYINPUT68), .A2(KEYINPUT6), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n241_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n214_), .A2(new_n215_), .A3(new_n249_), .A4(new_n250_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n246_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n225_), .A2(KEYINPUT8), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n245_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G29gat), .B(G36gat), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(G50gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(G43gat), .ZN(new_n260_));
  INV_X1    g059(.A(G43gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(G50gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT74), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n260_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n258_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n260_), .A2(new_n262_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT74), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n260_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(new_n257_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT15), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n266_), .A2(new_n270_), .A3(KEYINPUT15), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT75), .B1(new_n256_), .B2(new_n275_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n266_), .A2(new_n270_), .A3(KEYINPUT15), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT15), .B1(new_n266_), .B2(new_n270_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT75), .ZN(new_n280_));
  INV_X1    g079(.A(new_n250_), .ZN(new_n281_));
  OAI22_X1  g080(.A1(new_n218_), .A2(new_n213_), .B1(new_n281_), .B2(new_n248_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n253_), .A2(new_n242_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n246_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n255_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n241_), .A2(KEYINPUT8), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n234_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n230_), .A2(KEYINPUT10), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n228_), .A2(G99gat), .ZN(new_n290_));
  AOI21_X1  g089(.A(G106gat), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n287_), .B1(new_n292_), .B2(new_n236_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n285_), .B(new_n286_), .C1(new_n293_), .C2(new_n220_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n279_), .A2(new_n280_), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n212_), .B1(new_n276_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT77), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(KEYINPUT69), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n237_), .A2(new_n244_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n220_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT69), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n301_), .A2(new_n302_), .A3(new_n285_), .A4(new_n286_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n303_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n297_), .B1(new_n304_), .B2(new_n271_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n271_), .ZN(new_n306_));
  AOI211_X1 g105(.A(KEYINPUT77), .B(new_n306_), .C1(new_n298_), .C2(new_n303_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n296_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT80), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(KEYINPUT80), .B(new_n296_), .C1(new_n305_), .C2(new_n307_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT76), .ZN(new_n312_));
  INV_X1    g111(.A(new_n295_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n280_), .B1(new_n279_), .B2(new_n294_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n276_), .A2(KEYINPUT76), .A3(new_n295_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n315_), .B(new_n316_), .C1(new_n305_), .C2(new_n307_), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n310_), .A2(new_n311_), .B1(new_n209_), .B2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n205_), .B1(new_n318_), .B2(KEYINPUT81), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n209_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n303_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n255_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n302_), .B1(new_n322_), .B2(new_n285_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n271_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT77), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n304_), .A2(new_n297_), .A3(new_n271_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT80), .B1(new_n327_), .B2(new_n296_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n311_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n320_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT81), .ZN(new_n331_));
  INV_X1    g130(.A(new_n205_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT78), .B(KEYINPUT36), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n319_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n318_), .A2(KEYINPUT36), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n319_), .B2(new_n333_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n202_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n319_), .A2(new_n333_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n334_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n342_), .A2(KEYINPUT37), .A3(new_n336_), .A4(new_n335_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n339_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G15gat), .B(G22gat), .ZN(new_n346_));
  INV_X1    g145(.A(G1gat), .ZN(new_n347_));
  INV_X1    g146(.A(G8gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT14), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G1gat), .B(G8gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G231gat), .A2(G233gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n352_), .B(new_n353_), .Z(new_n354_));
  NOR2_X1   g153(.A1(KEYINPUT70), .A2(G71gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G78gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(KEYINPUT70), .A2(G71gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n356_), .A2(new_n357_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n358_), .ZN(new_n360_));
  OAI21_X1  g159(.A(G78gat), .B1(new_n360_), .B2(new_n355_), .ZN(new_n361_));
  INV_X1    g160(.A(G57gat), .ZN(new_n362_));
  INV_X1    g161(.A(G64gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G57gat), .A2(G64gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n359_), .A2(new_n361_), .A3(KEYINPUT11), .A4(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n359_), .A2(new_n361_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(KEYINPUT11), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT11), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n364_), .A2(new_n370_), .A3(new_n365_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n369_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n367_), .B1(new_n368_), .B2(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n354_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n354_), .A2(new_n373_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G127gat), .B(G155gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G211gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT16), .B(G183gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT17), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n379_), .A2(KEYINPUT17), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n374_), .A2(new_n375_), .A3(new_n380_), .A4(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT82), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n373_), .A2(KEYINPUT71), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT71), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n385_), .B(new_n367_), .C1(new_n368_), .C2(new_n372_), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n380_), .B1(new_n354_), .B2(new_n387_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n388_), .B1(new_n354_), .B2(new_n387_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n383_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT101), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G211gat), .B(G218gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT95), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G197gat), .A2(G204gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT94), .B(G204gat), .ZN(new_n396_));
  OAI211_X1 g195(.A(KEYINPUT21), .B(new_n395_), .C1(new_n396_), .C2(G197gat), .ZN(new_n397_));
  INV_X1    g196(.A(G197gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G204gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n394_), .B(new_n397_), .C1(KEYINPUT21), .C2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n392_), .B(KEYINPUT95), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(KEYINPUT21), .A3(new_n400_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT90), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT85), .B(G183gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT25), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT86), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(G183gat), .B1(KEYINPUT87), .B2(KEYINPUT25), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(KEYINPUT87), .B2(KEYINPUT25), .ZN(new_n412_));
  XOR2_X1   g211(.A(KEYINPUT26), .B(G190gat), .Z(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n407_), .A2(KEYINPUT86), .A3(KEYINPUT25), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n410_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(G169gat), .A2(G176gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT88), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT88), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n419_), .B1(G169gat), .B2(G176gat), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT24), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G183gat), .A2(G190gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT23), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G169gat), .A2(G176gat), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n418_), .A2(new_n420_), .A3(KEYINPUT24), .A4(new_n426_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n416_), .A2(new_n425_), .A3(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G190gat), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n407_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT22), .B(G169gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT89), .ZN(new_n432_));
  INV_X1    g231(.A(G176gat), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n432_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n436_));
  OAI221_X1 g235(.A(new_n426_), .B1(new_n430_), .B2(new_n424_), .C1(new_n435_), .C2(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n406_), .B1(new_n428_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n428_), .A2(new_n437_), .A3(new_n406_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n405_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G226gat), .A2(G233gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT19), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT20), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(KEYINPUT25), .B(G183gat), .Z(new_n446_));
  OAI21_X1  g245(.A(new_n427_), .B1(new_n413_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n425_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n447_), .B1(new_n448_), .B2(KEYINPUT99), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT99), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n425_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n431_), .B(KEYINPUT100), .Z(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n433_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(G183gat), .A2(G190gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n424_), .A2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n456_), .B1(G169gat), .B2(G176gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n452_), .A2(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n445_), .B1(new_n459_), .B2(new_n404_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n391_), .B1(new_n441_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n440_), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n462_), .A2(new_n404_), .A3(new_n438_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n449_), .A2(new_n451_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT20), .B1(new_n464_), .B2(new_n405_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n443_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n404_), .B1(new_n462_), .B2(new_n438_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n405_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n467_), .A2(KEYINPUT101), .A3(new_n468_), .A4(new_n445_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n461_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G64gat), .B(G92gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(G8gat), .B(G36gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT102), .B(KEYINPUT18), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n470_), .A2(new_n476_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n461_), .A2(new_n466_), .A3(new_n475_), .A4(new_n469_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT27), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT96), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n401_), .A2(new_n481_), .A3(new_n403_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n481_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT20), .B1(new_n484_), .B2(new_n459_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n443_), .B1(new_n485_), .B2(new_n441_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n465_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n443_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n439_), .A2(new_n440_), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n487_), .B(new_n488_), .C1(new_n489_), .C2(new_n404_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n486_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n480_), .B1(new_n491_), .B2(new_n476_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n479_), .A2(new_n480_), .B1(new_n492_), .B2(new_n478_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G22gat), .B(G50gat), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(G155gat), .ZN(new_n496_));
  INV_X1    g295(.A(G162gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(G155gat), .A2(G162gat), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G141gat), .A2(G148gat), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n501_), .B(KEYINPUT2), .Z(new_n502_));
  NOR2_X1   g301(.A1(G141gat), .A2(G148gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT3), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT3), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n503_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n500_), .B1(new_n502_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT1), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n499_), .B1(new_n498_), .B2(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT1), .B1(new_n496_), .B2(new_n497_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n504_), .A2(new_n501_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n509_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT28), .B1(new_n516_), .B2(KEYINPUT29), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n516_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n495_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n519_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(new_n517_), .A3(new_n494_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(G78gat), .B(G106gat), .Z(new_n525_));
  XOR2_X1   g324(.A(new_n525_), .B(KEYINPUT97), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n516_), .A2(KEYINPUT29), .ZN(new_n528_));
  INV_X1    g327(.A(G228gat), .ZN(new_n529_));
  INV_X1    g328(.A(G233gat), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n404_), .A2(new_n528_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n528_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n482_), .A2(new_n534_), .A3(new_n483_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n527_), .B(new_n533_), .C1(new_n535_), .C2(new_n532_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n524_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n484_), .A2(new_n528_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(new_n531_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n525_), .B1(new_n539_), .B2(new_n533_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT98), .B1(new_n537_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n525_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n535_), .A2(new_n532_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n533_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n542_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT98), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(new_n536_), .A4(new_n524_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n526_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n536_), .ZN(new_n549_));
  AOI22_X1  g348(.A1(new_n541_), .A2(new_n547_), .B1(new_n549_), .B2(new_n523_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G127gat), .B(G134gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G113gat), .B(G120gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(new_n516_), .B2(KEYINPUT103), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT103), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n509_), .A2(new_n515_), .A3(new_n553_), .A4(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(KEYINPUT4), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G225gat), .A2(G233gat), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n559_), .B(KEYINPUT104), .Z(new_n560_));
  INV_X1    g359(.A(KEYINPUT4), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n516_), .A2(new_n561_), .A3(new_n554_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n558_), .A2(new_n560_), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n560_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n555_), .A2(new_n564_), .A3(new_n557_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G1gat), .B(G29gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(G85gat), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT0), .B(G57gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n570_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n563_), .A2(new_n572_), .A3(new_n565_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G71gat), .B(G99gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT30), .B(G43gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n554_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n489_), .B(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(KEYINPUT93), .B(KEYINPUT31), .Z(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT92), .B(G15gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G227gat), .A2(G233gat), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT91), .Z(new_n585_));
  XNOR2_X1  g384(.A(new_n583_), .B(new_n585_), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n580_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n580_), .A2(new_n586_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n493_), .A2(new_n550_), .A3(new_n575_), .A4(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n541_), .A2(new_n547_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n549_), .A2(new_n523_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n574_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT105), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n573_), .A2(new_n594_), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n558_), .A2(new_n564_), .A3(new_n562_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT106), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n555_), .A2(new_n560_), .A3(new_n557_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n598_), .B2(new_n570_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n596_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n597_), .A3(new_n570_), .ZN(new_n601_));
  AOI22_X1  g400(.A1(new_n595_), .A2(KEYINPUT33), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n573_), .A2(new_n594_), .A3(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n477_), .A2(new_n602_), .A3(new_n478_), .A4(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n475_), .A2(KEYINPUT32), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n491_), .A2(new_n607_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n461_), .A2(new_n466_), .A3(new_n606_), .A4(new_n469_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n574_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n605_), .A2(new_n610_), .ZN(new_n611_));
  AOI22_X1  g410(.A1(new_n593_), .A2(new_n493_), .B1(new_n611_), .B2(new_n550_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n590_), .B1(new_n612_), .B2(new_n589_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n373_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n298_), .A2(new_n615_), .A3(new_n303_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT12), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n304_), .A2(new_n373_), .ZN(new_n619_));
  AND4_X1   g418(.A1(KEYINPUT12), .A2(new_n294_), .A3(new_n386_), .A4(new_n384_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G230gat), .A2(G233gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n618_), .A2(new_n619_), .A3(new_n621_), .A4(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n616_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n615_), .B1(new_n298_), .B2(new_n303_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n624_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(G176gat), .B(G204gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n626_), .A2(new_n629_), .A3(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT73), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT73), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n626_), .A2(new_n629_), .A3(new_n637_), .A4(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n626_), .A2(new_n629_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n634_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT13), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n279_), .A2(new_n352_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G229gat), .A2(G233gat), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n306_), .A2(new_n352_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n352_), .B(new_n271_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n648_), .B1(new_n649_), .B2(new_n646_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(G113gat), .B(G141gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G169gat), .B(G197gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT83), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n650_), .B(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT84), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n644_), .A2(new_n656_), .ZN(new_n657_));
  NOR4_X1   g456(.A1(new_n345_), .A2(new_n390_), .A3(new_n614_), .A4(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n347_), .A3(new_n574_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT38), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n655_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n644_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT107), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n664_), .A2(new_n390_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n342_), .A2(new_n336_), .A3(new_n335_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n614_), .A2(new_n666_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n347_), .B1(new_n668_), .B2(new_n574_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n661_), .A2(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n670_), .B1(new_n660_), .B2(new_n659_), .ZN(G1324gat));
  INV_X1    g470(.A(new_n493_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n658_), .A2(new_n348_), .A3(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n665_), .A2(new_n672_), .A3(new_n667_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT39), .ZN(new_n675_));
  AND3_X1   g474(.A1(new_n674_), .A2(new_n675_), .A3(G8gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n674_), .B2(G8gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n678_), .B(new_n680_), .ZN(G1325gat));
  INV_X1    g480(.A(G15gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n658_), .A2(new_n682_), .A3(new_n589_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n668_), .A2(new_n589_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G15gat), .ZN(new_n685_));
  XOR2_X1   g484(.A(KEYINPUT109), .B(KEYINPUT41), .Z(new_n686_));
  AND2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n685_), .A2(new_n686_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n683_), .B1(new_n687_), .B2(new_n688_), .ZN(G1326gat));
  INV_X1    g488(.A(G22gat), .ZN(new_n690_));
  INV_X1    g489(.A(new_n550_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n658_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n665_), .A2(new_n691_), .A3(new_n667_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n693_), .A2(new_n694_), .A3(G22gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n693_), .B2(G22gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(G1327gat));
  NAND2_X1  g498(.A1(new_n666_), .A2(new_n390_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n614_), .A2(new_n700_), .A3(new_n657_), .ZN(new_n701_));
  AOI21_X1  g500(.A(G29gat), .B1(new_n701_), .B2(new_n574_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n339_), .A2(new_n613_), .A3(new_n343_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n339_), .A2(new_n613_), .A3(KEYINPUT43), .A4(new_n343_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n705_), .A2(new_n390_), .A3(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT111), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n664_), .A2(KEYINPUT111), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n708_), .A2(new_n709_), .A3(new_n710_), .ZN(new_n711_));
  OAI211_X1 g510(.A(KEYINPUT111), .B(KEYINPUT44), .C1(new_n707_), .C2(new_n664_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n574_), .A2(G29gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n702_), .B1(new_n713_), .B2(new_n714_), .ZN(G1328gat));
  INV_X1    g514(.A(G36gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n701_), .A2(new_n716_), .A3(new_n672_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT45), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n493_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(new_n716_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT46), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  OAI211_X1 g521(.A(KEYINPUT46), .B(new_n718_), .C1(new_n719_), .C2(new_n716_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(G1329gat));
  NAND3_X1  g523(.A1(new_n713_), .A2(G43gat), .A3(new_n589_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n701_), .A2(new_n589_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n725_), .B(new_n726_), .C1(G43gat), .C2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n589_), .ZN(new_n729_));
  AOI211_X1 g528(.A(new_n261_), .B(new_n729_), .C1(new_n711_), .C2(new_n712_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n727_), .A2(G43gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT47), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n728_), .A2(new_n732_), .ZN(G1330gat));
  AOI21_X1  g532(.A(G50gat), .B1(new_n701_), .B2(new_n691_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n550_), .A2(new_n259_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n713_), .B2(new_n735_), .ZN(G1331gat));
  NOR2_X1   g535(.A1(new_n644_), .A2(new_n662_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NOR4_X1   g537(.A1(new_n345_), .A2(new_n390_), .A3(new_n614_), .A4(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G57gat), .B1(new_n739_), .B2(new_n574_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n656_), .A2(new_n390_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NOR4_X1   g541(.A1(new_n614_), .A2(new_n666_), .A3(new_n644_), .A4(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n575_), .A2(new_n362_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1332gat));
  NAND3_X1  g544(.A1(new_n739_), .A2(new_n363_), .A3(new_n672_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n672_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G64gat), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(KEYINPUT48), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(KEYINPUT48), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(G1333gat));
  INV_X1    g550(.A(G71gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n739_), .A2(new_n752_), .A3(new_n589_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n743_), .A2(new_n589_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G71gat), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(KEYINPUT49), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(KEYINPUT49), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(G1334gat));
  NAND3_X1  g557(.A1(new_n739_), .A2(new_n357_), .A3(new_n691_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n743_), .A2(new_n691_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G78gat), .ZN(new_n761_));
  XOR2_X1   g560(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n762_));
  AND2_X1   g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n761_), .A2(new_n762_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n759_), .B1(new_n763_), .B2(new_n764_), .ZN(G1335gat));
  NOR3_X1   g564(.A1(new_n614_), .A2(new_n738_), .A3(new_n700_), .ZN(new_n766_));
  AOI21_X1  g565(.A(G85gat), .B1(new_n766_), .B2(new_n574_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n707_), .A2(new_n738_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n575_), .A2(new_n223_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n767_), .B1(new_n768_), .B2(new_n769_), .ZN(G1336gat));
  AOI21_X1  g569(.A(G92gat), .B1(new_n766_), .B2(new_n672_), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n672_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n768_), .B2(new_n772_), .ZN(G1337gat));
  OAI211_X1 g572(.A(new_n766_), .B(new_n589_), .C1(new_n229_), .C2(new_n231_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n707_), .A2(new_n729_), .A3(new_n738_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n230_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n766_), .A2(new_n227_), .A3(new_n691_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n390_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n780_), .A2(new_n691_), .A3(new_n706_), .A4(new_n737_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n781_), .A2(new_n782_), .A3(G106gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n781_), .B2(G106gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n778_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g585(.A(G113gat), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n646_), .B1(new_n645_), .B2(new_n647_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n649_), .A2(new_n646_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n653_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n653_), .B2(new_n650_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n639_), .B2(new_n642_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n628_), .A2(new_n620_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n625_), .B1(new_n795_), .B2(new_n618_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n626_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n795_), .A2(KEYINPUT55), .A3(new_n625_), .A4(new_n618_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  AND4_X1   g599(.A1(new_n794_), .A2(new_n800_), .A3(KEYINPUT56), .A4(new_n641_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT114), .B1(new_n639_), .B2(new_n662_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT114), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n803_), .B(new_n655_), .C1(new_n636_), .C2(new_n638_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n801_), .A2(new_n802_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n800_), .A2(new_n641_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT56), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n800_), .A2(KEYINPUT56), .A3(new_n641_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(KEYINPUT115), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n793_), .B1(new_n805_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n788_), .B1(new_n811_), .B2(new_n666_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n808_), .A2(new_n809_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n792_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT58), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n813_), .A2(KEYINPUT58), .A3(new_n814_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n339_), .A2(new_n343_), .A3(new_n817_), .A4(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n337_), .A2(new_n338_), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n807_), .B(new_n634_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n794_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n639_), .A2(new_n662_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n803_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n639_), .A2(KEYINPUT114), .A3(new_n662_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n822_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT56), .B1(new_n800_), .B2(new_n641_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n827_), .A2(new_n821_), .A3(new_n794_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n820_), .B(KEYINPUT57), .C1(new_n829_), .C2(new_n793_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n812_), .A2(new_n819_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n390_), .ZN(new_n832_));
  XOR2_X1   g631(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n833_));
  NAND2_X1  g632(.A1(new_n643_), .A2(KEYINPUT13), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n643_), .A2(KEYINPUT13), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n741_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n833_), .B1(new_n344_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n833_), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n837_), .B(new_n840_), .C1(new_n339_), .C2(new_n343_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n839_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n691_), .B1(new_n832_), .B2(new_n842_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n672_), .A2(new_n575_), .A3(new_n729_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n787_), .B1(new_n845_), .B2(new_n655_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n845_), .A2(KEYINPUT59), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n843_), .A2(new_n850_), .A3(new_n844_), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n849_), .A2(G113gat), .A3(new_n656_), .A4(new_n851_), .ZN(new_n852_));
  OAI211_X1 g651(.A(KEYINPUT116), .B(new_n787_), .C1(new_n845_), .C2(new_n655_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n848_), .A2(new_n852_), .A3(new_n853_), .ZN(G1340gat));
  INV_X1    g653(.A(new_n644_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n849_), .A2(new_n855_), .A3(new_n851_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(G120gat), .ZN(new_n857_));
  INV_X1    g656(.A(new_n845_), .ZN(new_n858_));
  INV_X1    g657(.A(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n644_), .B2(KEYINPUT60), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n858_), .B(new_n860_), .C1(KEYINPUT60), .C2(new_n859_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n857_), .A2(new_n861_), .ZN(G1341gat));
  AOI21_X1  g661(.A(G127gat), .B1(new_n858_), .B2(new_n779_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n849_), .A2(new_n851_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n779_), .A2(G127gat), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(KEYINPUT117), .Z(new_n866_));
  AOI21_X1  g665(.A(new_n863_), .B1(new_n864_), .B2(new_n866_), .ZN(G1342gat));
  AOI21_X1  g666(.A(G134gat), .B1(new_n858_), .B2(new_n666_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT118), .B(G134gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n344_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n868_), .B1(new_n864_), .B2(new_n870_), .ZN(G1343gat));
  NAND2_X1  g670(.A1(new_n832_), .A2(new_n842_), .ZN(new_n872_));
  NOR4_X1   g671(.A1(new_n672_), .A2(new_n550_), .A3(new_n575_), .A4(new_n589_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n662_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g675(.A1(new_n872_), .A2(new_n873_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n644_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT119), .B(G148gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1345gat));
  XNOR2_X1  g679(.A(KEYINPUT61), .B(G155gat), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n874_), .A2(new_n779_), .A3(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n881_), .B1(new_n877_), .B2(new_n390_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT120), .B(KEYINPUT121), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n883_), .A2(new_n886_), .A3(new_n884_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1346gat));
  AOI21_X1  g689(.A(G162gat), .B1(new_n874_), .B2(new_n666_), .ZN(new_n891_));
  NOR3_X1   g690(.A1(new_n877_), .A2(new_n497_), .A3(new_n344_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(G1347gat));
  NOR3_X1   g692(.A1(new_n493_), .A2(new_n574_), .A3(new_n729_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n872_), .A2(new_n550_), .A3(new_n662_), .A4(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n895_), .A2(new_n896_), .A3(G169gat), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT122), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n895_), .A2(G169gat), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(KEYINPUT62), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n895_), .A2(KEYINPUT122), .A3(new_n896_), .A4(G169gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n899_), .A2(new_n901_), .A3(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n872_), .A2(new_n550_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n894_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n906_), .A2(new_n453_), .A3(new_n662_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n903_), .A2(new_n907_), .ZN(G1348gat));
  AOI21_X1  g707(.A(G176gat), .B1(new_n906_), .B2(new_n855_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n904_), .A2(KEYINPUT123), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n843_), .A2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n905_), .B1(new_n910_), .B2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n644_), .A2(new_n433_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n909_), .B1(new_n913_), .B2(new_n914_), .ZN(G1349gat));
  AND3_X1   g714(.A1(new_n906_), .A2(new_n779_), .A3(new_n446_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n913_), .A2(new_n779_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n407_), .ZN(G1350gat));
  INV_X1    g717(.A(new_n906_), .ZN(new_n919_));
  OAI21_X1  g718(.A(G190gat), .B1(new_n919_), .B2(new_n344_), .ZN(new_n920_));
  OR2_X1    g719(.A1(new_n820_), .A2(new_n413_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n919_), .B2(new_n921_), .ZN(G1351gat));
  NOR4_X1   g721(.A1(new_n493_), .A2(new_n550_), .A3(new_n574_), .A4(new_n589_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n872_), .A2(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n655_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(KEYINPUT124), .B(G197gat), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n925_), .B(new_n926_), .ZN(G1352gat));
  AND2_X1   g726(.A1(new_n872_), .A2(new_n923_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n855_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(G204gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n930_), .B1(new_n396_), .B2(new_n929_), .ZN(G1353gat));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n390_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n933_));
  AND3_X1   g732(.A1(new_n928_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n932_), .B1(new_n928_), .B2(new_n933_), .ZN(new_n935_));
  OAI22_X1  g734(.A1(new_n934_), .A2(new_n935_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n928_), .A2(new_n933_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(KEYINPUT125), .ZN(new_n938_));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n928_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n938_), .A2(new_n939_), .A3(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n936_), .A2(new_n941_), .ZN(G1354gat));
  XOR2_X1   g741(.A(KEYINPUT127), .B(G218gat), .Z(new_n943_));
  AND3_X1   g742(.A1(new_n928_), .A2(new_n345_), .A3(new_n943_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n924_), .A2(new_n820_), .ZN(new_n945_));
  OR2_X1    g744(.A1(new_n945_), .A2(KEYINPUT126), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n943_), .B1(new_n945_), .B2(KEYINPUT126), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n944_), .B1(new_n946_), .B2(new_n947_), .ZN(G1355gat));
endmodule


