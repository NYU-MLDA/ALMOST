//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n910_, new_n911_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G71gat), .B(G99gat), .Z(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  AND2_X1   g008(.A1(KEYINPUT78), .A2(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT22), .ZN(new_n211_));
  AOI21_X1  g010(.A(G176gat), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(KEYINPUT78), .A2(G169gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT22), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n209_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(G183gat), .B2(G190gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n216_), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT79), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT79), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n220_), .A2(new_n216_), .A3(G183gat), .A4(G190gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n217_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n215_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT25), .B(G183gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT26), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n226_), .A2(KEYINPUT77), .A3(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT77), .ZN(new_n228_));
  INV_X1    g027(.A(G190gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT26), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n225_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n208_), .A2(KEYINPUT24), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G183gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT23), .B1(new_n237_), .B2(new_n229_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(new_n218_), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n231_), .A2(new_n234_), .A3(new_n236_), .A4(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n224_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT30), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT80), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT30), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n224_), .A2(new_n244_), .A3(new_n240_), .ZN(new_n245_));
  AND3_X1   g044(.A1(new_n242_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n243_), .B1(new_n242_), .B2(new_n245_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n207_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G127gat), .B(G134gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G113gat), .B(G120gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT31), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT81), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n242_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n206_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n248_), .A2(new_n253_), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n248_), .B2(new_n255_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(G78gat), .B(G106gat), .Z(new_n259_));
  NAND2_X1  g058(.A1(G228gat), .A2(G233gat), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT88), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G141gat), .B(G148gat), .Z(new_n263_));
  OR2_X1    g062(.A1(G155gat), .A2(G162gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G155gat), .A2(G162gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT82), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT82), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(G155gat), .A3(G162gat), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT83), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n264_), .B(new_n270_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  AOI211_X1 g072(.A(KEYINPUT83), .B(new_n269_), .C1(new_n266_), .C2(new_n268_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n263_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT84), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G141gat), .A2(G148gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT2), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT2), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(G141gat), .A3(G148gat), .ZN(new_n280_));
  AND2_X1   g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT3), .ZN(new_n282_));
  INV_X1    g081(.A(G141gat), .ZN(new_n283_));
  INV_X1    g082(.A(G148gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n282_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n276_), .B1(new_n281_), .B2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n267_), .B1(G155gat), .B2(G162gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n265_), .A2(KEYINPUT82), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n264_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT85), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT85), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n293_), .B(new_n264_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n278_), .A2(new_n280_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n295_), .A2(KEYINPUT84), .A3(new_n286_), .A4(new_n285_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n288_), .A2(new_n292_), .A3(new_n294_), .A4(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n275_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT29), .ZN(new_n299_));
  INV_X1    g098(.A(G204gat), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(KEYINPUT86), .A3(G197gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(G197gat), .ZN(new_n302_));
  INV_X1    g101(.A(G197gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(G204gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  OAI211_X1 g104(.A(KEYINPUT21), .B(new_n301_), .C1(new_n305_), .C2(KEYINPUT86), .ZN(new_n306_));
  AND2_X1   g105(.A1(KEYINPUT87), .A2(KEYINPUT21), .ZN(new_n307_));
  NOR2_X1   g106(.A1(KEYINPUT87), .A2(KEYINPUT21), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G197gat), .B(G204gat), .ZN(new_n310_));
  INV_X1    g109(.A(G211gat), .ZN(new_n311_));
  INV_X1    g110(.A(G218gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G211gat), .A2(G218gat), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n309_), .A2(new_n310_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n313_), .A2(KEYINPUT21), .A3(new_n314_), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n306_), .A2(new_n315_), .B1(new_n305_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n262_), .B1(new_n299_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT29), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n320_), .B1(new_n275_), .B2(new_n297_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n260_), .B(KEYINPUT88), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NOR3_X1   g122(.A1(new_n321_), .A2(new_n317_), .A3(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n259_), .B1(new_n319_), .B2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n299_), .A2(new_n318_), .A3(new_n322_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n259_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n262_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n328_), .B1(new_n321_), .B2(new_n317_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n326_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n275_), .A2(new_n297_), .A3(new_n320_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT28), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT28), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n275_), .A2(new_n297_), .A3(new_n333_), .A4(new_n320_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G22gat), .B(G50gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n332_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n334_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n335_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n325_), .A2(new_n330_), .A3(new_n336_), .A4(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n330_), .A2(KEYINPUT89), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n327_), .B1(new_n326_), .B2(new_n329_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n339_), .A2(new_n336_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT89), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n346_), .B(new_n259_), .C1(new_n319_), .C2(new_n324_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT90), .B1(new_n344_), .B2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n325_), .A2(KEYINPUT89), .A3(new_n330_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT90), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(new_n345_), .A4(new_n347_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n341_), .B1(new_n349_), .B2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n275_), .A2(new_n297_), .A3(KEYINPUT93), .ZN(new_n354_));
  INV_X1    g153(.A(new_n251_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n275_), .A2(new_n297_), .A3(KEYINPUT93), .A4(new_n251_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(KEYINPUT4), .A3(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G225gat), .A2(G233gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT4), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n298_), .A2(new_n361_), .A3(new_n355_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(new_n360_), .A3(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n356_), .A2(new_n359_), .A3(new_n357_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G1gat), .B(G29gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT94), .B(G85gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT0), .B(G57gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n365_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n363_), .A2(new_n364_), .A3(new_n370_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT96), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G8gat), .B(G36gat), .ZN(new_n376_));
  INV_X1    g175(.A(G92gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT18), .B(G64gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT20), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n236_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n222_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n226_), .A2(new_n229_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n385_), .A2(KEYINPUT91), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT91), .B1(new_n385_), .B2(new_n386_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n225_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n239_), .B1(G183gat), .B2(G190gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT22), .B(G169gat), .ZN(new_n391_));
  INV_X1    g190(.A(G176gat), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n209_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n384_), .A2(new_n389_), .B1(new_n390_), .B2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n382_), .B1(new_n394_), .B2(new_n317_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G226gat), .A2(G233gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT19), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n318_), .A2(new_n241_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n395_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n317_), .A2(new_n224_), .A3(new_n240_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n401_), .B(KEYINPUT20), .C1(new_n394_), .C2(new_n317_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n402_), .A2(KEYINPUT92), .A3(new_n397_), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT92), .B1(new_n402_), .B2(new_n397_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n381_), .B(new_n400_), .C1(new_n403_), .C2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n399_), .B1(new_n395_), .B2(KEYINPUT95), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT95), .ZN(new_n408_));
  AOI211_X1 g207(.A(new_n408_), .B(new_n382_), .C1(new_n394_), .C2(new_n317_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n397_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n402_), .A2(new_n397_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n381_), .B1(new_n410_), .B2(new_n412_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n406_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n363_), .A2(KEYINPUT96), .A3(new_n364_), .A4(new_n370_), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n375_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n400_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n380_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n380_), .B(new_n400_), .C1(new_n403_), .C2(new_n404_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n358_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n356_), .A2(new_n360_), .A3(new_n357_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n371_), .A3(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n419_), .A2(new_n420_), .A3(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n373_), .A2(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n373_), .A2(new_n425_), .ZN(new_n427_));
  NOR3_X1   g226(.A1(new_n424_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n353_), .B1(new_n416_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n352_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n345_), .A2(new_n347_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n351_), .B1(new_n431_), .B2(new_n350_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n340_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n375_), .A2(new_n415_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n419_), .A2(new_n420_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT27), .ZN(new_n436_));
  INV_X1    g235(.A(new_n400_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n402_), .A2(new_n397_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT92), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n402_), .A2(KEYINPUT92), .A3(new_n397_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n437_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n436_), .B1(new_n442_), .B2(new_n380_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n410_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n418_), .B1(new_n444_), .B2(new_n411_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n435_), .A2(new_n436_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n433_), .A2(new_n434_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n429_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n258_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n353_), .A2(new_n449_), .A3(new_n446_), .A4(new_n434_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT97), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  AOI211_X1 g251(.A(new_n258_), .B(new_n341_), .C1(new_n349_), .C2(new_n352_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n453_), .A2(KEYINPUT97), .A3(new_n434_), .A4(new_n446_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n258_), .A2(new_n448_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT76), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G1gat), .B(G8gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT73), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G15gat), .B(G22gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G1gat), .A2(G8gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(KEYINPUT14), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n458_), .A2(new_n462_), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n457_), .A2(KEYINPUT73), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n457_), .A2(KEYINPUT73), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n464_), .A2(new_n461_), .A3(new_n459_), .A4(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G29gat), .B(G36gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G43gat), .B(G50gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n470_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n468_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n467_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n473_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n475_), .B1(new_n463_), .B2(new_n466_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n476_), .A2(KEYINPUT75), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n474_), .B(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G229gat), .A2(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT15), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n475_), .B(new_n482_), .ZN(new_n483_));
  AND2_X1   g282(.A1(new_n463_), .A2(new_n466_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n476_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n479_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G113gat), .B(G141gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G169gat), .B(G197gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n481_), .A2(new_n486_), .A3(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n490_), .B1(new_n481_), .B2(new_n486_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n456_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n493_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(KEYINPUT76), .A3(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n455_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT98), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G120gat), .B(G148gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(new_n300_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT5), .B(G176gat), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n502_), .B(new_n503_), .Z(new_n504_));
  XNOR2_X1  g303(.A(G57gat), .B(G64gat), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n505_), .A2(KEYINPUT11), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(KEYINPUT11), .ZN(new_n507_));
  XOR2_X1   g306(.A(G71gat), .B(G78gat), .Z(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  OR2_X1    g308(.A1(new_n507_), .A2(new_n508_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT7), .ZN(new_n513_));
  INV_X1    g312(.A(G99gat), .ZN(new_n514_));
  INV_X1    g313(.A(G106gat), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G99gat), .A2(G106gat), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n516_), .A2(new_n519_), .A3(new_n520_), .A4(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G85gat), .B(G92gat), .Z(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT8), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT8), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n522_), .A2(new_n526_), .A3(new_n523_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  XOR2_X1   g328(.A(KEYINPUT10), .B(G99gat), .Z(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(new_n515_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n531_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n532_));
  INV_X1    g331(.A(G85gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n377_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT65), .B(G85gat), .ZN(new_n537_));
  AOI21_X1  g336(.A(KEYINPUT9), .B1(new_n537_), .B2(G92gat), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT66), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n536_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n533_), .A2(KEYINPUT65), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT65), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(G85gat), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n543_), .A3(G92gat), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT9), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT66), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n532_), .B1(new_n540_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n512_), .B1(new_n529_), .B2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n544_), .A2(new_n539_), .A3(new_n545_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n536_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n547_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n531_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n553_));
  AOI22_X1  g352(.A1(new_n552_), .A2(new_n553_), .B1(new_n525_), .B2(new_n527_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(new_n511_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n549_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G230gat), .A2(G233gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT64), .Z(new_n558_));
  NAND2_X1  g357(.A1(new_n556_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT67), .B(KEYINPUT12), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n560_), .B1(new_n554_), .B2(new_n511_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(KEYINPUT67), .A2(KEYINPUT12), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n512_), .B(new_n563_), .C1(new_n529_), .C2(new_n548_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n558_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n561_), .A2(new_n564_), .A3(new_n565_), .A4(new_n555_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n504_), .B1(new_n559_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n559_), .A2(new_n566_), .A3(new_n504_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT69), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(KEYINPUT68), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n569_), .B2(KEYINPUT68), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n568_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n573_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(new_n567_), .A3(new_n571_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n577_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT70), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT13), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n574_), .A2(new_n576_), .A3(new_n582_), .A4(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n581_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G231gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n467_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(new_n511_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G127gat), .B(G155gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(new_n311_), .ZN(new_n590_));
  XOR2_X1   g389(.A(KEYINPUT16), .B(G183gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT17), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n588_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n588_), .A2(KEYINPUT17), .A3(new_n592_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT74), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n596_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n594_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  NAND2_X1  g403(.A1(new_n554_), .A2(new_n475_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n605_), .B1(new_n554_), .B2(new_n483_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT72), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n609_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n606_), .A2(new_n607_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT34), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n606_), .A2(new_n615_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n610_), .A2(new_n612_), .A3(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n614_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n601_), .B(new_n604_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n612_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n611_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n615_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n610_), .A2(new_n612_), .A3(new_n616_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n604_), .A2(new_n601_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n604_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT36), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .A4(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n619_), .A2(KEYINPUT37), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(KEYINPUT37), .B1(new_n619_), .B2(new_n627_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n600_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n585_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n500_), .A2(new_n631_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n632_), .A2(G1gat), .A3(new_n434_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(KEYINPUT38), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n635_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n638_));
  INV_X1    g437(.A(new_n455_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n619_), .A2(new_n627_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT100), .Z(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT101), .ZN(new_n643_));
  INV_X1    g442(.A(new_n585_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n644_), .A2(new_n498_), .A3(new_n600_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n434_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n638_), .B1(new_n649_), .B2(G1gat), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n636_), .B(new_n637_), .C1(new_n650_), .C2(new_n633_), .ZN(G1324gat));
  OR3_X1    g450(.A1(new_n632_), .A2(G8gat), .A3(new_n446_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n446_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n643_), .A2(new_n653_), .A3(new_n645_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT39), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n654_), .A2(new_n655_), .A3(G8gat), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n655_), .B1(new_n654_), .B2(G8gat), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n652_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g458(.A(G15gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n647_), .B2(new_n449_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n662_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n449_), .A2(new_n660_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n663_), .B(new_n664_), .C1(new_n632_), .C2(new_n665_), .ZN(G1326gat));
  OR3_X1    g465(.A1(new_n632_), .A2(G22gat), .A3(new_n353_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n647_), .A2(new_n433_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n668_), .A2(new_n669_), .A3(G22gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n668_), .B2(G22gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n667_), .B1(new_n670_), .B2(new_n671_), .ZN(G1327gat));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n581_), .A2(new_n497_), .A3(new_n584_), .A4(new_n600_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT102), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n628_), .A2(new_n629_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT43), .B1(new_n677_), .B2(KEYINPUT103), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n679_), .B1(new_n455_), .B2(new_n677_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n677_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n452_), .A2(new_n454_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n449_), .B1(new_n429_), .B2(new_n447_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n681_), .B(new_n678_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n676_), .B1(new_n680_), .B2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n673_), .B1(new_n685_), .B2(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n680_), .A2(new_n684_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n676_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(KEYINPUT104), .A3(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n692_));
  AND4_X1   g491(.A1(new_n692_), .A2(new_n687_), .A3(KEYINPUT44), .A4(new_n688_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n685_), .B2(KEYINPUT44), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n686_), .B(new_n691_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(KEYINPUT106), .B1(new_n695_), .B2(new_n434_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT104), .B1(new_n689_), .B2(new_n690_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n685_), .A2(new_n673_), .A3(KEYINPUT44), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n687_), .A2(KEYINPUT44), .A3(new_n688_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT105), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n685_), .A2(new_n692_), .A3(KEYINPUT44), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n699_), .A2(new_n700_), .A3(new_n648_), .A4(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n696_), .A2(G29gat), .A3(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n641_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n600_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n708_), .A2(new_n644_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n500_), .A2(new_n709_), .ZN(new_n710_));
  OR3_X1    g509(.A1(new_n710_), .A2(G29gat), .A3(new_n434_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n706_), .A2(new_n711_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT107), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n706_), .A2(new_n714_), .A3(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1328gat));
  INV_X1    g515(.A(KEYINPUT108), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n717_), .B1(new_n695_), .B2(new_n446_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n699_), .A2(KEYINPUT108), .A3(new_n653_), .A4(new_n704_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(G36gat), .A3(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n446_), .B(KEYINPUT109), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n710_), .A2(G36gat), .A3(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n720_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT110), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(KEYINPUT46), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(new_n729_));
  OAI211_X1 g528(.A(new_n720_), .B(new_n725_), .C1(new_n727_), .C2(KEYINPUT46), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1329gat));
  OAI21_X1  g530(.A(G43gat), .B1(new_n695_), .B2(new_n258_), .ZN(new_n732_));
  OR3_X1    g531(.A1(new_n710_), .A2(G43gat), .A3(new_n258_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g534(.A(G50gat), .B1(new_n695_), .B2(new_n353_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n353_), .A2(G50gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n710_), .B2(new_n737_), .ZN(G1331gat));
  NOR3_X1   g537(.A1(new_n585_), .A2(new_n497_), .A3(new_n600_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n643_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(G57gat), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n434_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n455_), .A2(new_n497_), .A3(new_n585_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n630_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n434_), .B1(new_n744_), .B2(KEYINPUT111), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n745_), .B1(KEYINPUT111), .B2(new_n744_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n742_), .B1(new_n741_), .B2(new_n746_), .ZN(G1332gat));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748_));
  INV_X1    g547(.A(new_n740_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n721_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n748_), .B1(new_n750_), .B2(G64gat), .ZN(new_n751_));
  INV_X1    g550(.A(G64gat), .ZN(new_n752_));
  AOI211_X1 g551(.A(KEYINPUT48), .B(new_n752_), .C1(new_n749_), .C2(new_n721_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n721_), .A2(new_n752_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT112), .ZN(new_n755_));
  OAI22_X1  g554(.A1(new_n751_), .A2(new_n753_), .B1(new_n744_), .B2(new_n755_), .ZN(G1333gat));
  INV_X1    g555(.A(KEYINPUT49), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n749_), .A2(new_n449_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n758_), .B2(G71gat), .ZN(new_n759_));
  INV_X1    g558(.A(G71gat), .ZN(new_n760_));
  AOI211_X1 g559(.A(KEYINPUT49), .B(new_n760_), .C1(new_n749_), .C2(new_n449_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n449_), .A2(new_n760_), .ZN(new_n762_));
  OAI22_X1  g561(.A1(new_n759_), .A2(new_n761_), .B1(new_n744_), .B2(new_n762_), .ZN(G1334gat));
  OR3_X1    g562(.A1(new_n744_), .A2(G78gat), .A3(new_n353_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n749_), .A2(new_n433_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(G78gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(G78gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(G1335gat));
  NAND3_X1  g568(.A1(new_n743_), .A2(new_n707_), .A3(new_n600_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(G85gat), .B1(new_n771_), .B2(new_n648_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n687_), .A2(KEYINPUT113), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n585_), .A2(new_n497_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n600_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n687_), .A2(KEYINPUT113), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n773_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n648_), .A2(new_n537_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n772_), .B1(new_n779_), .B2(new_n780_), .ZN(G1336gat));
  AOI21_X1  g580(.A(G92gat), .B1(new_n771_), .B2(new_n653_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n722_), .A2(new_n377_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n779_), .B2(new_n783_), .ZN(G1337gat));
  OAI21_X1  g583(.A(G99gat), .B1(new_n778_), .B2(new_n258_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n771_), .A2(new_n449_), .A3(new_n530_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI211_X1 g587(.A(new_n353_), .B(new_n775_), .C1(new_n680_), .C2(new_n684_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(new_n515_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT52), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n790_), .B(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n771_), .A2(new_n515_), .A3(new_n433_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g594(.A1(new_n631_), .A2(new_n498_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT54), .Z(new_n797_));
  NAND2_X1  g596(.A1(new_n497_), .A2(new_n569_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n566_), .B2(KEYINPUT114), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT55), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n561_), .A2(new_n555_), .A3(new_n564_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n566_), .B2(new_n799_), .ZN(new_n804_));
  OAI221_X1 g603(.A(new_n801_), .B1(new_n565_), .B2(new_n802_), .C1(new_n800_), .C2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n504_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT56), .B1(new_n805_), .B2(new_n806_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n798_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n810_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(new_n808_), .A3(new_n807_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n577_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n478_), .A2(new_n479_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n485_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n480_), .B1(new_n485_), .B2(new_n817_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n816_), .B(new_n489_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n820_), .A2(KEYINPUT118), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(KEYINPUT118), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n492_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n815_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n814_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n641_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OR2_X1    g627(.A1(new_n807_), .A2(KEYINPUT119), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n829_), .A2(new_n569_), .A3(new_n823_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n812_), .A2(KEYINPUT119), .A3(new_n807_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT58), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(new_n677_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(KEYINPUT58), .A3(new_n831_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n825_), .A2(KEYINPUT57), .A3(new_n641_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n828_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n797_), .B1(new_n837_), .B2(new_n600_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n453_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n653_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n648_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n838_), .A2(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(G113gat), .B1(new_n842_), .B2(new_n497_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n837_), .A2(new_n600_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n797_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847_));
  INV_X1    g646(.A(new_n841_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n846_), .A2(new_n847_), .A3(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT59), .B1(new_n838_), .B2(new_n841_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n497_), .A2(G113gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n843_), .B1(new_n851_), .B2(new_n852_), .ZN(G1340gat));
  NAND3_X1  g652(.A1(new_n849_), .A2(new_n850_), .A3(new_n644_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G120gat), .ZN(new_n855_));
  INV_X1    g654(.A(new_n842_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT60), .ZN(new_n857_));
  AOI21_X1  g656(.A(G120gat), .B1(new_n644_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n859_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n857_), .A2(G120gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n855_), .B1(new_n856_), .B2(new_n863_), .ZN(G1341gat));
  AOI21_X1  g663(.A(G127gat), .B1(new_n842_), .B2(new_n599_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n599_), .A2(G127gat), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n851_), .B2(new_n866_), .ZN(G1342gat));
  INV_X1    g666(.A(G134gat), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n677_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n849_), .A2(new_n850_), .A3(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n846_), .A2(new_n707_), .A3(new_n848_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n868_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n870_), .A2(KEYINPUT121), .A3(new_n872_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1343gat));
  NOR2_X1   g676(.A1(new_n353_), .A2(new_n449_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n722_), .A2(new_n648_), .A3(new_n878_), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n879_), .B(KEYINPUT122), .Z(new_n880_));
  NAND3_X1  g679(.A1(new_n846_), .A2(KEYINPUT123), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n882_));
  INV_X1    g681(.A(new_n880_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n838_), .B2(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n498_), .B1(new_n881_), .B2(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(new_n283_), .ZN(G1344gat));
  AOI21_X1  g685(.A(new_n585_), .B1(new_n881_), .B2(new_n884_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT124), .B(G148gat), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n887_), .B(new_n889_), .ZN(G1345gat));
  NAND2_X1  g689(.A1(new_n881_), .A2(new_n884_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT61), .B(G155gat), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n891_), .A2(new_n599_), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n891_), .B2(new_n599_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1346gat));
  AOI21_X1  g694(.A(G162gat), .B1(new_n891_), .B2(new_n707_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n681_), .A2(G162gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n891_), .B2(new_n897_), .ZN(G1347gat));
  NOR2_X1   g697(.A1(new_n838_), .A2(new_n722_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n839_), .A2(new_n648_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(G169gat), .B1(new_n901_), .B2(new_n498_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT62), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  OAI211_X1 g703(.A(KEYINPUT62), .B(G169gat), .C1(new_n901_), .C2(new_n498_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n899_), .A2(new_n391_), .A3(new_n497_), .A4(new_n900_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n904_), .A2(new_n905_), .A3(new_n906_), .ZN(G1348gat));
  NOR2_X1   g706(.A1(new_n901_), .A2(new_n585_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(new_n392_), .ZN(G1349gat));
  NOR2_X1   g708(.A1(new_n901_), .A2(new_n600_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n225_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n911_), .B1(new_n237_), .B2(new_n910_), .ZN(G1350gat));
  NOR2_X1   g711(.A1(new_n387_), .A2(new_n388_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n641_), .A2(new_n913_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n899_), .A2(new_n900_), .A3(new_n914_), .ZN(new_n915_));
  AND4_X1   g714(.A1(new_n681_), .A2(new_n846_), .A3(new_n721_), .A4(new_n900_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n916_), .B2(new_n229_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(KEYINPUT125), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n919_), .B(new_n915_), .C1(new_n916_), .C2(new_n229_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n920_), .ZN(G1351gat));
  NAND2_X1  g720(.A1(new_n878_), .A2(new_n434_), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n838_), .A2(new_n722_), .A3(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n497_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n644_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g726(.A1(new_n923_), .A2(new_n599_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT63), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n928_), .A2(new_n929_), .A3(new_n311_), .ZN(new_n930_));
  XOR2_X1   g729(.A(KEYINPUT63), .B(G211gat), .Z(new_n931_));
  NAND3_X1  g730(.A1(new_n923_), .A2(new_n599_), .A3(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n923_), .A2(KEYINPUT126), .A3(new_n599_), .A4(new_n931_), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n930_), .A2(new_n934_), .A3(new_n935_), .ZN(G1354gat));
  NOR2_X1   g735(.A1(new_n641_), .A2(G218gat), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n923_), .A2(new_n937_), .ZN(new_n938_));
  NOR4_X1   g737(.A1(new_n838_), .A2(new_n677_), .A3(new_n722_), .A4(new_n922_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n939_), .B2(new_n312_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(KEYINPUT127), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n938_), .B(new_n942_), .C1(new_n312_), .C2(new_n939_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1355gat));
endmodule


