//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n902_, new_n903_, new_n905_, new_n906_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT70), .ZN(new_n203_));
  INV_X1    g002(.A(G29gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(G36gat), .ZN(new_n205_));
  INV_X1    g004(.A(G36gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(G29gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n203_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(G29gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n204_), .A2(G36gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT70), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G43gat), .B(G50gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n212_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n202_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n208_), .A2(new_n211_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n212_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(new_n213_), .A3(KEYINPUT15), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G106gat), .ZN(new_n222_));
  OR2_X1    g021(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n224_));
  AND3_X1   g023(.A1(new_n223_), .A2(KEYINPUT64), .A3(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(KEYINPUT64), .B1(new_n223_), .B2(new_n224_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n222_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT6), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(G85gat), .A2(G92gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT9), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT65), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT9), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n233_), .A2(new_n235_), .A3(new_n237_), .A4(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT66), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n234_), .A2(KEYINPUT65), .A3(G85gat), .A4(G92gat), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n240_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n227_), .B(new_n232_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT7), .ZN(new_n245_));
  INV_X1    g044(.A(G99gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(new_n222_), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n247_), .A2(new_n230_), .A3(new_n231_), .A4(new_n248_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n233_), .A2(new_n238_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT8), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT8), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(new_n253_), .A3(new_n250_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n244_), .A2(new_n255_), .ZN(new_n256_));
  AND3_X1   g055(.A1(new_n221_), .A2(new_n256_), .A3(KEYINPUT71), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT71), .B1(new_n221_), .B2(new_n256_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n219_), .A2(new_n213_), .ZN(new_n259_));
  OAI22_X1  g058(.A1(new_n257_), .A2(new_n258_), .B1(new_n259_), .B2(new_n256_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n221_), .A2(new_n256_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n221_), .A2(new_n256_), .A3(KEYINPUT71), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT72), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G232gat), .A2(G233gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT35), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n260_), .B1(new_n265_), .B2(new_n269_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n268_), .A2(KEYINPUT35), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n272_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n269_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n271_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n270_), .B1(new_n275_), .B2(new_n260_), .ZN(new_n276_));
  XOR2_X1   g075(.A(G134gat), .B(G162gat), .Z(new_n277_));
  XNOR2_X1  g076(.A(G190gat), .B(G218gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT36), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT73), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT74), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n276_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT75), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n279_), .B(KEYINPUT36), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n270_), .B(new_n287_), .C1(new_n275_), .C2(new_n260_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n276_), .A2(KEYINPUT75), .A3(new_n283_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n286_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT37), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n284_), .A2(new_n291_), .A3(new_n288_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT76), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT76), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n284_), .A2(new_n294_), .A3(new_n291_), .A4(new_n288_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(KEYINPUT37), .A2(new_n290_), .B1(new_n293_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G57gat), .B(G64gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G71gat), .B(G78gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n298_), .A2(new_n299_), .A3(KEYINPUT11), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(KEYINPUT11), .ZN(new_n301_));
  INV_X1    g100(.A(new_n299_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n298_), .A2(KEYINPUT11), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n300_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G231gat), .A2(G233gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT77), .ZN(new_n308_));
  XOR2_X1   g107(.A(G1gat), .B(G8gat), .Z(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G15gat), .B(G22gat), .ZN(new_n311_));
  INV_X1    g110(.A(G1gat), .ZN(new_n312_));
  INV_X1    g111(.A(G8gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT14), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n309_), .A2(new_n314_), .A3(new_n311_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n308_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n308_), .A2(new_n318_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  XOR2_X1   g120(.A(G127gat), .B(G155gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT16), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G183gat), .B(G211gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT17), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n325_), .A2(new_n326_), .ZN(new_n328_));
  OR4_X1    g127(.A1(new_n319_), .A2(new_n321_), .A3(new_n327_), .A4(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n327_), .B1(new_n321_), .B2(new_n319_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n297_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n333_), .B(KEYINPUT78), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G190gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT80), .B(G183gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT25), .ZN(new_n338_));
  OR2_X1    g137(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n336_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT24), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT81), .ZN(new_n343_));
  NOR3_X1   g142(.A1(new_n343_), .A2(G169gat), .A3(G176gat), .ZN(new_n344_));
  INV_X1    g143(.A(G169gat), .ZN(new_n345_));
  INV_X1    g144(.A(G176gat), .ZN(new_n346_));
  AOI21_X1  g145(.A(KEYINPUT81), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n342_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT23), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n345_), .A2(new_n346_), .A3(KEYINPUT81), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n343_), .B1(G169gat), .B2(G176gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(KEYINPUT24), .A4(new_n353_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n348_), .A2(new_n350_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n341_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n350_), .B1(G190gat), .B2(new_n337_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n353_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT22), .B(G169gat), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(new_n346_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n356_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT30), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n363_), .A2(KEYINPUT83), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(KEYINPUT83), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G227gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT82), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G71gat), .B(G99gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G15gat), .B(G43gat), .Z(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n364_), .A2(new_n365_), .A3(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n365_), .A2(new_n371_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT85), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT85), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n372_), .A2(new_n376_), .A3(new_n373_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G127gat), .B(G134gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G113gat), .B(G120gat), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT84), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n378_), .B(new_n379_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n380_), .B1(new_n381_), .B2(KEYINPUT84), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT31), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n375_), .A2(new_n377_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n383_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n374_), .A2(KEYINPUT85), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT18), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G64gat), .B(G92gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(KEYINPUT32), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT20), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT92), .B(G204gat), .ZN(new_n395_));
  INV_X1    g194(.A(G197gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT94), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT21), .ZN(new_n398_));
  NOR2_X1   g197(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT94), .ZN(new_n401_));
  NAND2_X1  g200(.A1(KEYINPUT92), .A2(G204gat), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(G197gat), .A4(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT91), .B(G197gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(G204gat), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n397_), .A2(new_n398_), .A3(new_n403_), .A4(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G211gat), .B(G218gat), .ZN(new_n407_));
  AND2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n395_), .A2(new_n396_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT93), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n395_), .A2(KEYINPUT93), .A3(new_n396_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n404_), .ZN(new_n413_));
  INV_X1    g212(.A(G204gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n411_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT21), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n397_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n407_), .A2(new_n398_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n408_), .A2(new_n417_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  XOR2_X1   g219(.A(KEYINPUT25), .B(G183gat), .Z(new_n421_));
  OAI21_X1  g220(.A(new_n355_), .B1(new_n336_), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n350_), .B1(G183gat), .B2(G190gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n360_), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n394_), .B1(new_n420_), .B2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n418_), .A2(new_n419_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n409_), .A2(new_n410_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n398_), .B1(new_n428_), .B2(new_n412_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n406_), .A2(new_n407_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n427_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT96), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n431_), .A2(new_n432_), .A3(new_n362_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n432_), .B1(new_n431_), .B2(new_n362_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n426_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G226gat), .A2(G233gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n436_), .B(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT100), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n422_), .A2(new_n424_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n431_), .A2(new_n440_), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n341_), .A2(new_n355_), .B1(new_n360_), .B2(new_n357_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n442_), .B(new_n427_), .C1(new_n429_), .C2(new_n430_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n438_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n441_), .A2(new_n443_), .A3(KEYINPUT20), .A4(new_n444_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n435_), .A2(new_n438_), .B1(new_n439_), .B2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n394_), .B1(new_n431_), .B2(new_n440_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n447_), .A2(KEYINPUT100), .A3(new_n444_), .A4(new_n443_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n393_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n449_));
  OAI211_X1 g248(.A(new_n426_), .B(new_n444_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n443_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n438_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(new_n452_), .A3(new_n393_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G1gat), .B(G29gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(G85gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(KEYINPUT0), .B(G57gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(G155gat), .A2(G162gat), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G155gat), .A2(G162gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT87), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n461_), .A2(new_n462_), .A3(KEYINPUT1), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(new_n461_), .B2(KEYINPUT1), .ZN(new_n464_));
  OAI221_X1 g263(.A(new_n460_), .B1(KEYINPUT1), .B2(new_n461_), .C1(new_n463_), .C2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G141gat), .A2(G148gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT86), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(G141gat), .A3(G148gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(G141gat), .ZN(new_n471_));
  INV_X1    g270(.A(G148gat), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n465_), .A2(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n460_), .A2(new_n461_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n470_), .A2(KEYINPUT2), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT3), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n477_), .A2(new_n471_), .A3(new_n472_), .A4(KEYINPUT88), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT88), .ZN(new_n479_));
  OAI22_X1  g278(.A1(new_n479_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n475_), .B1(new_n476_), .B2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n474_), .A2(new_n381_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n381_), .A2(KEYINPUT84), .ZN(new_n485_));
  INV_X1    g284(.A(new_n380_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n480_), .A2(new_n481_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n488_), .B(new_n478_), .C1(KEYINPUT2), .C2(new_n470_), .ZN(new_n489_));
  AOI22_X1  g288(.A1(new_n489_), .A2(new_n475_), .B1(new_n465_), .B2(new_n473_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n484_), .B(KEYINPUT4), .C1(new_n487_), .C2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G225gat), .A2(G233gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n492_), .B(KEYINPUT97), .Z(new_n493_));
  AND2_X1   g292(.A1(new_n491_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n474_), .A2(new_n483_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT4), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n382_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT98), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n495_), .A2(new_n382_), .A3(KEYINPUT98), .A4(new_n496_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n494_), .A2(new_n501_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n484_), .B(new_n492_), .C1(new_n487_), .C2(new_n490_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n458_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n503_), .ZN(new_n505_));
  AOI211_X1 g304(.A(new_n457_), .B(new_n505_), .C1(new_n494_), .C2(new_n501_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n453_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(KEYINPUT101), .B1(new_n449_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n445_), .A2(new_n439_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT20), .B1(new_n431_), .B2(new_n440_), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT96), .B1(new_n420_), .B2(new_n442_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n431_), .A2(new_n432_), .A3(new_n362_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n510_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n509_), .B(new_n448_), .C1(new_n513_), .C2(new_n444_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(KEYINPUT32), .A3(new_n392_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n502_), .A2(new_n503_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n457_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n502_), .A2(new_n458_), .A3(new_n503_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT101), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n515_), .A2(new_n519_), .A3(new_n520_), .A4(new_n453_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT99), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(KEYINPUT33), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n484_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n458_), .B1(new_n526_), .B2(new_n493_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n501_), .A2(new_n492_), .A3(new_n491_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n506_), .A2(new_n524_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n450_), .A2(new_n452_), .A3(new_n392_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n392_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n518_), .A2(new_n523_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n529_), .A2(new_n530_), .A3(new_n532_), .A4(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n508_), .A2(new_n521_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(G78gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n495_), .A2(KEYINPUT29), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n431_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n536_), .B1(new_n431_), .B2(new_n537_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n222_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n540_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n542_), .A2(G106gat), .A3(new_n538_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G22gat), .B(G50gat), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n495_), .A2(KEYINPUT29), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n549_), .A2(KEYINPUT28), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(KEYINPUT28), .ZN(new_n551_));
  INV_X1    g350(.A(G233gat), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT89), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n553_), .A2(G228gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(G228gat), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n552_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n556_), .B(KEYINPUT90), .Z(new_n557_));
  AND3_X1   g356(.A1(new_n550_), .A2(new_n551_), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n557_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n559_));
  OAI22_X1  g358(.A1(new_n547_), .A2(new_n548_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n548_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n558_), .A2(new_n559_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(new_n546_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n535_), .A2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n392_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n530_), .A2(KEYINPUT27), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT102), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n530_), .A2(KEYINPUT27), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT102), .ZN(new_n571_));
  INV_X1    g370(.A(new_n392_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n514_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n569_), .A2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n519_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT27), .B1(new_n532_), .B2(new_n530_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n575_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n388_), .B1(new_n566_), .B2(new_n579_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n567_), .A2(KEYINPUT102), .A3(new_n568_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n571_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n578_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT103), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n575_), .A2(KEYINPUT103), .A3(new_n578_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n564_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n387_), .A2(new_n519_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n580_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G113gat), .B(G141gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G169gat), .B(G197gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n318_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n594_), .A2(KEYINPUT79), .A3(new_n213_), .A4(new_n219_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT79), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n596_), .B1(new_n259_), .B2(new_n318_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n221_), .A2(new_n318_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G229gat), .A2(G233gat), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n259_), .A2(new_n318_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n600_), .B1(new_n598_), .B2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n593_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n598_), .A2(new_n603_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n592_), .B(new_n601_), .C1(new_n606_), .C2(new_n600_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n589_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n244_), .A2(new_n255_), .A3(new_n305_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G230gat), .A2(G233gat), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n611_), .A2(KEYINPUT68), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT68), .B1(new_n611_), .B2(new_n612_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT12), .ZN(new_n615_));
  INV_X1    g414(.A(new_n305_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n256_), .B2(new_n616_), .ZN(new_n617_));
  AOI211_X1 g416(.A(KEYINPUT12), .B(new_n305_), .C1(new_n244_), .C2(new_n255_), .ZN(new_n618_));
  OAI22_X1  g417(.A1(new_n613_), .A2(new_n614_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n256_), .A2(new_n616_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT67), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n621_), .A3(new_n611_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n612_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n256_), .A2(KEYINPUT67), .A3(new_n616_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n622_), .A2(new_n623_), .A3(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n619_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G120gat), .B(G148gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT5), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n628_), .B(new_n629_), .Z(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n626_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n619_), .A2(new_n625_), .A3(new_n631_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT13), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n334_), .A2(new_n610_), .A3(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n636_), .A2(new_n312_), .A3(new_n519_), .ZN(new_n637_));
  XOR2_X1   g436(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n284_), .A2(new_n288_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n589_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n635_), .A2(new_n608_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(new_n331_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT105), .ZN(new_n645_));
  INV_X1    g444(.A(new_n519_), .ZN(new_n646_));
  OAI21_X1  g445(.A(G1gat), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n639_), .A2(new_n647_), .ZN(G1324gat));
  AOI21_X1  g447(.A(KEYINPUT103), .B1(new_n575_), .B2(new_n578_), .ZN(new_n649_));
  AOI211_X1 g448(.A(new_n584_), .B(new_n577_), .C1(new_n569_), .C2(new_n574_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n636_), .A2(new_n313_), .A3(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n641_), .A2(new_n651_), .A3(new_n643_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G8gat), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(KEYINPUT106), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n653_), .A2(new_n657_), .A3(G8gat), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n655_), .A2(new_n656_), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n656_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n652_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT40), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  OAI211_X1 g462(.A(KEYINPUT40), .B(new_n652_), .C1(new_n659_), .C2(new_n660_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1325gat));
  OAI21_X1  g464(.A(G15gat), .B1(new_n645_), .B2(new_n387_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT41), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(G15gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n636_), .A2(new_n669_), .A3(new_n388_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n668_), .A2(new_n670_), .ZN(G1326gat));
  OAI21_X1  g470(.A(G22gat), .B1(new_n645_), .B2(new_n565_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT42), .ZN(new_n673_));
  INV_X1    g472(.A(G22gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n636_), .A2(new_n674_), .A3(new_n564_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1327gat));
  INV_X1    g475(.A(new_n635_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n331_), .A2(new_n640_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n610_), .A2(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(G29gat), .B1(new_n680_), .B2(new_n519_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n642_), .A2(new_n332_), .ZN(new_n682_));
  OR2_X1    g481(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n589_), .B2(new_n297_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n566_), .A2(new_n579_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(new_n387_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n588_), .B(new_n565_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT107), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .A4(new_n296_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n684_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n297_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n689_), .B1(new_n693_), .B2(new_n690_), .ZN(new_n694_));
  OAI211_X1 g493(.A(new_n682_), .B(new_n683_), .C1(new_n692_), .C2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n688_), .A2(new_n690_), .A3(new_n296_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT107), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n698_), .A2(new_n684_), .A3(new_n691_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n683_), .B1(new_n699_), .B2(new_n682_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n696_), .A2(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n646_), .A2(new_n204_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n681_), .B1(new_n701_), .B2(new_n702_), .ZN(G1328gat));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n206_), .B1(new_n701_), .B2(new_n651_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT45), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n651_), .B(KEYINPUT109), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n610_), .A2(new_n206_), .A3(new_n679_), .A4(new_n707_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(KEYINPUT110), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(KEYINPUT110), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  OR2_X1    g510(.A1(new_n708_), .A2(KEYINPUT110), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n708_), .A2(KEYINPUT110), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n712_), .A2(KEYINPUT45), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n704_), .B1(new_n705_), .B2(new_n715_), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n711_), .A2(new_n714_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n651_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n696_), .A2(new_n700_), .A3(new_n718_), .ZN(new_n719_));
  OAI211_X1 g518(.A(new_n717_), .B(KEYINPUT46), .C1(new_n206_), .C2(new_n719_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n716_), .A2(new_n720_), .ZN(G1329gat));
  INV_X1    g520(.A(G43gat), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n387_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n701_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n680_), .A2(new_n388_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n724_), .A2(new_n726_), .A3(new_n728_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1330gat));
  AOI21_X1  g531(.A(G50gat), .B1(new_n680_), .B2(new_n564_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n564_), .A2(G50gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n701_), .B2(new_n734_), .ZN(G1331gat));
  NOR2_X1   g534(.A1(new_n589_), .A2(new_n608_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n334_), .A2(new_n736_), .A3(new_n677_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT112), .Z(new_n738_));
  AOI21_X1  g537(.A(G57gat), .B1(new_n738_), .B2(new_n519_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n331_), .A2(new_n608_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n641_), .A2(new_n677_), .A3(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n741_), .A2(G57gat), .A3(new_n519_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT113), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n739_), .A2(new_n743_), .ZN(G1332gat));
  NAND2_X1  g543(.A1(new_n741_), .A2(new_n707_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(G64gat), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT48), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n737_), .B(KEYINPUT112), .ZN(new_n748_));
  INV_X1    g547(.A(new_n707_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n749_), .A2(G64gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n747_), .B1(new_n748_), .B2(new_n750_), .ZN(G1333gat));
  INV_X1    g550(.A(G71gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n741_), .B2(new_n388_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT49), .Z(new_n754_));
  NAND2_X1  g553(.A1(new_n388_), .A2(new_n752_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT114), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n748_), .B2(new_n756_), .ZN(G1334gat));
  NAND2_X1  g556(.A1(new_n741_), .A2(new_n564_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(G78gat), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT50), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n759_), .B(new_n760_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n748_), .A2(G78gat), .A3(new_n565_), .ZN(new_n762_));
  OAI21_X1  g561(.A(KEYINPUT115), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n759_), .B(KEYINPUT50), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n738_), .A2(new_n536_), .A3(new_n564_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n763_), .A2(new_n767_), .ZN(G1335gat));
  NOR3_X1   g567(.A1(new_n635_), .A2(new_n332_), .A3(new_n608_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n699_), .A2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(G85gat), .B1(new_n770_), .B2(new_n646_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n635_), .A2(new_n678_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n736_), .A2(new_n772_), .ZN(new_n773_));
  OR2_X1    g572(.A1(new_n646_), .A2(G85gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n771_), .B1(new_n773_), .B2(new_n774_), .ZN(G1336gat));
  OAI21_X1  g574(.A(G92gat), .B1(new_n770_), .B2(new_n749_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n718_), .A2(G92gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n773_), .B2(new_n777_), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n770_), .B2(new_n387_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n388_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n779_), .B1(new_n773_), .B2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g581(.A1(new_n736_), .A2(new_n222_), .A3(new_n564_), .A4(new_n772_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n699_), .A2(new_n564_), .A3(new_n769_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(G106gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G106gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT53), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n790_), .B(new_n783_), .C1(new_n786_), .C2(new_n787_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1339gat));
  INV_X1    g591(.A(KEYINPUT59), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794_));
  AND3_X1   g593(.A1(new_n608_), .A2(new_n794_), .A3(new_n633_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n608_), .B2(new_n633_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n619_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n611_), .A2(new_n612_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT68), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n611_), .A2(KEYINPUT68), .A3(new_n612_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n620_), .A2(KEYINPUT12), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n256_), .A2(new_n615_), .A3(new_n616_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n805_), .A2(new_n808_), .A3(KEYINPUT117), .A4(KEYINPUT55), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n800_), .A2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n611_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n619_), .A2(new_n799_), .B1(new_n811_), .B2(new_n623_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT56), .B1(new_n813_), .B2(new_n630_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  AOI211_X1 g614(.A(new_n815_), .B(new_n631_), .C1(new_n810_), .C2(new_n812_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n797_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n600_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n598_), .A2(new_n599_), .A3(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n593_), .B(new_n819_), .C1(new_n606_), .C2(new_n818_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n607_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n821_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n640_), .B1(new_n817_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT57), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n811_), .A2(new_n623_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n803_), .A2(new_n804_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(KEYINPUT55), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n800_), .B2(new_n809_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n815_), .B1(new_n831_), .B2(new_n631_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n813_), .A2(KEYINPUT56), .A3(new_n630_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n822_), .B1(new_n834_), .B2(new_n797_), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT118), .B(new_n827_), .C1(new_n835_), .C2(new_n640_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n821_), .B1(new_n626_), .B2(new_n631_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(KEYINPUT58), .A3(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT58), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n296_), .A2(new_n838_), .A3(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n826_), .A2(new_n836_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n635_), .A2(new_n740_), .ZN(new_n844_));
  OR3_X1    g643(.A1(new_n296_), .A2(new_n844_), .A3(KEYINPUT54), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT54), .B1(new_n296_), .B2(new_n844_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n843_), .A2(new_n331_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT120), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n793_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n387_), .A2(new_n646_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n850_), .B(new_n565_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT119), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n847_), .A2(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n849_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n843_), .A2(new_n331_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n845_), .A2(new_n846_), .ZN(new_n857_));
  AOI221_X4 g656(.A(new_n853_), .B1(new_n848_), .B2(new_n793_), .C1(new_n856_), .C2(new_n857_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n855_), .A2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G113gat), .B1(new_n859_), .B2(new_n609_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n856_), .A2(new_n857_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n853_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  OR3_X1    g662(.A1(new_n863_), .A2(G113gat), .A3(new_n609_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n860_), .A2(new_n864_), .ZN(G1340gat));
  INV_X1    g664(.A(G120gat), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n635_), .B2(KEYINPUT60), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(KEYINPUT121), .Z(new_n868_));
  OAI211_X1 g667(.A(new_n854_), .B(new_n868_), .C1(KEYINPUT60), .C2(new_n866_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT122), .ZN(new_n870_));
  OAI21_X1  g669(.A(G120gat), .B1(new_n859_), .B2(new_n635_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1341gat));
  INV_X1    g671(.A(G127gat), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n331_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(KEYINPUT123), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n861_), .A2(KEYINPUT120), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n863_), .A3(new_n793_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n849_), .A2(new_n854_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n875_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n873_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n863_), .A2(new_n331_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n879_), .A2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT124), .B1(new_n881_), .B2(new_n884_), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n880_), .B(new_n874_), .C1(new_n855_), .C2(new_n858_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(G127gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n882_), .B1(new_n859_), .B2(new_n875_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT124), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n885_), .A2(new_n890_), .ZN(G1342gat));
  OAI21_X1  g690(.A(G134gat), .B1(new_n859_), .B2(new_n297_), .ZN(new_n892_));
  INV_X1    g691(.A(G134gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n854_), .A2(new_n893_), .A3(new_n640_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(G1343gat));
  NOR2_X1   g694(.A1(new_n847_), .A2(new_n388_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n896_), .A2(new_n519_), .A3(new_n564_), .A4(new_n749_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n609_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n471_), .ZN(G1344gat));
  NOR2_X1   g698(.A1(new_n897_), .A2(new_n635_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(new_n472_), .ZN(G1345gat));
  NOR2_X1   g700(.A1(new_n897_), .A2(new_n331_), .ZN(new_n902_));
  XOR2_X1   g701(.A(KEYINPUT61), .B(G155gat), .Z(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1346gat));
  OAI21_X1  g703(.A(G162gat), .B1(new_n897_), .B2(new_n297_), .ZN(new_n905_));
  INV_X1    g704(.A(G162gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n640_), .A2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n905_), .B1(new_n897_), .B2(new_n907_), .ZN(G1347gat));
  NAND2_X1  g707(.A1(new_n707_), .A2(new_n588_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(KEYINPUT125), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n847_), .A2(new_n564_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n608_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G169gat), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n913_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n912_), .A2(new_n359_), .A3(new_n608_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n916_), .A2(new_n917_), .A3(new_n918_), .ZN(G1348gat));
  AOI21_X1  g718(.A(G176gat), .B1(new_n912_), .B2(new_n677_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n911_), .B(KEYINPUT126), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n910_), .A2(G176gat), .A3(new_n677_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n921_), .B2(new_n922_), .ZN(G1349gat));
  NAND3_X1  g722(.A1(new_n921_), .A2(new_n332_), .A3(new_n910_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n337_), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n332_), .A2(new_n421_), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n924_), .A2(new_n925_), .B1(new_n912_), .B2(new_n926_), .ZN(G1350gat));
  INV_X1    g726(.A(new_n912_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G190gat), .B1(new_n928_), .B2(new_n297_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n640_), .A2(new_n335_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT127), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n929_), .B1(new_n928_), .B2(new_n931_), .ZN(G1351gat));
  NAND3_X1  g731(.A1(new_n896_), .A2(new_n576_), .A3(new_n707_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n609_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(new_n396_), .ZN(G1352gat));
  NOR2_X1   g734(.A1(new_n933_), .A2(new_n635_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(G204gat), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n937_), .B1(new_n395_), .B2(new_n936_), .ZN(G1353gat));
  NOR2_X1   g737(.A1(new_n933_), .A2(new_n331_), .ZN(new_n939_));
  NOR3_X1   g738(.A1(new_n939_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940_));
  XOR2_X1   g739(.A(KEYINPUT63), .B(G211gat), .Z(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n939_), .B2(new_n941_), .ZN(G1354gat));
  OAI21_X1  g741(.A(G218gat), .B1(new_n933_), .B2(new_n297_), .ZN(new_n943_));
  INV_X1    g742(.A(G218gat), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n640_), .A2(new_n944_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n943_), .B1(new_n933_), .B2(new_n945_), .ZN(G1355gat));
endmodule


