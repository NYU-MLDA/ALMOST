//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n807_, new_n808_,
    new_n809_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n962_, new_n963_, new_n964_, new_n965_,
    new_n966_, new_n967_, new_n968_, new_n969_, new_n970_, new_n972_,
    new_n973_, new_n975_, new_n976_, new_n977_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n992_, new_n993_;
  INV_X1    g000(.A(KEYINPUT101), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT29), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT88), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT88), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(new_n208_), .A3(KEYINPUT1), .ZN(new_n209_));
  OR2_X1    g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n206_), .A2(new_n207_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n211_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT89), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT2), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n214_), .A2(new_n217_), .A3(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n212_), .A2(new_n223_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n219_), .A2(new_n221_), .A3(new_n222_), .A4(new_n224_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n210_), .A2(new_n204_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n203_), .B1(new_n216_), .B2(new_n227_), .ZN(new_n228_));
  AND2_X1   g027(.A1(G228gat), .A2(G233gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT21), .ZN(new_n230_));
  INV_X1    g029(.A(G204gat), .ZN(new_n231_));
  INV_X1    g030(.A(G197gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT91), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT91), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G197gat), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n231_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(G197gat), .A2(G204gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n230_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(G218gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(G211gat), .ZN(new_n240_));
  INV_X1    g039(.A(G211gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(G218gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n233_), .A2(new_n235_), .A3(new_n231_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n230_), .B1(G197gat), .B2(G204gat), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n236_), .A2(new_n237_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n230_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n248_));
  AOI22_X1  g047(.A1(new_n238_), .A2(new_n246_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n228_), .A2(new_n229_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n216_), .A2(new_n227_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT92), .B(KEYINPUT29), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n238_), .A2(new_n246_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n247_), .A2(new_n248_), .ZN(new_n255_));
  AND3_X1   g054(.A1(new_n254_), .A2(KEYINPUT93), .A3(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(KEYINPUT93), .B1(new_n254_), .B2(new_n255_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n253_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n250_), .B1(new_n258_), .B2(new_n229_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G78gat), .B(G106gat), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT94), .B1(new_n259_), .B2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n261_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n259_), .A2(KEYINPUT94), .A3(new_n261_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G22gat), .B(G50gat), .Z(new_n267_));
  OAI21_X1  g066(.A(new_n267_), .B1(new_n251_), .B2(KEYINPUT29), .ZN(new_n268_));
  AOI22_X1  g067(.A1(new_n225_), .A2(new_n226_), .B1(new_n211_), .B2(new_n215_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n267_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(new_n203_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n272_), .B(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n266_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT95), .ZN(new_n277_));
  INV_X1    g076(.A(new_n275_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n278_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT95), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AOI211_X1 g080(.A(new_n260_), .B(new_n250_), .C1(new_n229_), .C2(new_n258_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n282_), .A2(new_n275_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT96), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n284_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n285_));
  OR3_X1    g084(.A1(new_n259_), .A2(new_n284_), .A3(new_n261_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n283_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n277_), .A2(new_n281_), .A3(new_n287_), .ZN(new_n288_));
  XOR2_X1   g087(.A(G8gat), .B(G36gat), .Z(new_n289_));
  XNOR2_X1  g088(.A(new_n289_), .B(KEYINPUT18), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G64gat), .B(G92gat), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G226gat), .A2(G233gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT19), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G183gat), .A2(G190gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT26), .B(G190gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT25), .B(G183gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n300_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(G169gat), .ZN(new_n304_));
  INV_X1    g103(.A(G176gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(KEYINPUT24), .A3(new_n307_), .ZN(new_n308_));
  OR3_X1    g107(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n298_), .B(new_n299_), .C1(G183gat), .C2(G190gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n307_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(KEYINPUT22), .B(G169gat), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n312_), .B1(new_n313_), .B2(new_n305_), .ZN(new_n314_));
  AOI22_X1  g113(.A1(new_n303_), .A2(new_n310_), .B1(new_n311_), .B2(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n295_), .B1(new_n249_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT85), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT22), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G169gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n304_), .A2(KEYINPUT22), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n317_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n317_), .B1(new_n304_), .B2(KEYINPUT22), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n305_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT86), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(G176gat), .B1(new_n319_), .B2(new_n317_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT86), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n325_), .B(new_n326_), .C1(new_n317_), .C2(new_n313_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n300_), .ZN(new_n329_));
  OR2_X1    g128(.A1(KEYINPUT83), .A2(G183gat), .ZN(new_n330_));
  INV_X1    g129(.A(G190gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(KEYINPUT83), .A2(G183gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n312_), .B1(new_n329_), .B2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n330_), .A2(KEYINPUT25), .A3(new_n332_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT26), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(KEYINPUT84), .A3(G190gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(G190gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT84), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT25), .ZN(new_n341_));
  AOI22_X1  g140(.A1(new_n341_), .A2(G183gat), .B1(new_n331_), .B2(KEYINPUT26), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n335_), .A2(new_n337_), .A3(new_n340_), .A4(new_n342_), .ZN(new_n343_));
  AND4_X1   g142(.A1(new_n298_), .A2(new_n308_), .A3(new_n299_), .A4(new_n309_), .ZN(new_n344_));
  AOI22_X1  g143(.A1(new_n328_), .A2(new_n334_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n316_), .B(KEYINPUT20), .C1(new_n345_), .C2(new_n249_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n295_), .B(KEYINPUT97), .Z(new_n348_));
  INV_X1    g147(.A(KEYINPUT20), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n254_), .A2(new_n255_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n303_), .A2(new_n310_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n314_), .A2(new_n311_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n349_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n328_), .A2(new_n334_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n344_), .A2(new_n343_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(new_n249_), .A3(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n348_), .B1(new_n354_), .B2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n293_), .B1(new_n347_), .B2(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n354_), .A2(new_n357_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n292_), .B(new_n346_), .C1(new_n360_), .C2(new_n348_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G1gat), .B(G29gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G57gat), .B(G85gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G127gat), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n369_), .A2(G134gat), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(G134gat), .ZN(new_n371_));
  INV_X1    g170(.A(G113gat), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n372_), .A2(G120gat), .ZN(new_n373_));
  INV_X1    g172(.A(G120gat), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n374_), .A2(G113gat), .ZN(new_n375_));
  OAI22_X1  g174(.A1(new_n370_), .A2(new_n371_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G127gat), .B(G134gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G113gat), .B(G120gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n376_), .A2(new_n379_), .A3(KEYINPUT87), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT87), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n377_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n251_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n376_), .A2(new_n379_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n216_), .A2(new_n227_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n368_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n380_), .A2(new_n382_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n386_), .B(KEYINPUT4), .C1(new_n390_), .C2(new_n269_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT98), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n384_), .A2(KEYINPUT98), .A3(KEYINPUT4), .A4(new_n386_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n384_), .A2(KEYINPUT4), .ZN(new_n396_));
  INV_X1    g195(.A(new_n388_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n389_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n362_), .A2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n387_), .A2(new_n397_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n393_), .A2(new_n394_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n397_), .B1(new_n384_), .B2(KEYINPUT4), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n402_), .B(new_n367_), .C1(new_n403_), .C2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT33), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n408_), .A2(new_n401_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n409_), .A2(KEYINPUT33), .A3(new_n367_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n400_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n256_), .A2(new_n257_), .A3(new_n353_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT20), .B1(new_n345_), .B2(new_n249_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n295_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT100), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT100), .ZN(new_n416_));
  OAI211_X1 g215(.A(new_n416_), .B(new_n295_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n360_), .A2(new_n348_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n292_), .A2(KEYINPUT32), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n368_), .B1(new_n408_), .B2(new_n401_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n405_), .A2(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n420_), .B(new_n346_), .C1(new_n360_), .C2(new_n348_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n422_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n411_), .A2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n202_), .B1(new_n288_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n361_), .A2(KEYINPUT27), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n419_), .B2(new_n293_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT27), .B1(new_n359_), .B2(new_n361_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n405_), .A2(KEYINPUT102), .A3(new_n423_), .ZN(new_n433_));
  AOI21_X1  g232(.A(KEYINPUT102), .B1(new_n405_), .B2(new_n423_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n287_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n436_));
  AOI211_X1 g235(.A(KEYINPUT95), .B(new_n278_), .C1(new_n264_), .C2(new_n265_), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n432_), .B(new_n435_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n283_), .A2(new_n285_), .A3(new_n286_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n276_), .B2(KEYINPUT95), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n411_), .A2(new_n426_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(KEYINPUT101), .A4(new_n281_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n428_), .A2(new_n438_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G227gat), .A2(G233gat), .ZN(new_n444_));
  INV_X1    g243(.A(G15gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n444_), .B(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT30), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT31), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G71gat), .B(G99gat), .ZN(new_n449_));
  INV_X1    g248(.A(G43gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OR2_X1    g251(.A1(new_n345_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n345_), .A2(new_n452_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n383_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n453_), .A2(new_n383_), .A3(new_n454_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n448_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n457_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n448_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n459_), .A2(new_n455_), .A3(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT103), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n463_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n431_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n414_), .A2(KEYINPUT100), .B1(new_n348_), .B2(new_n360_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n292_), .B1(new_n466_), .B2(new_n417_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n465_), .B(KEYINPUT103), .C1(new_n467_), .C2(new_n429_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n464_), .A2(new_n468_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n433_), .A2(new_n462_), .A3(new_n434_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n469_), .A2(new_n281_), .A3(new_n440_), .A4(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT104), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n436_), .A2(new_n437_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT104), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n473_), .A2(new_n469_), .A3(new_n474_), .A4(new_n470_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n443_), .A2(new_n462_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G1gat), .B(G8gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G1gat), .ZN(new_n479_));
  INV_X1    g278(.A(G8gat), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT14), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n478_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n481_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(new_n477_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G29gat), .B(G36gat), .Z(new_n487_));
  XOR2_X1   g286(.A(G43gat), .B(G50gat), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G29gat), .B(G36gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT75), .B(KEYINPUT15), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n489_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n489_), .B2(new_n492_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n486_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G229gat), .A2(G233gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n489_), .A2(new_n492_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n498_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT79), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n486_), .A2(new_n492_), .A3(new_n489_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n499_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n497_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT79), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n496_), .A2(new_n506_), .A3(new_n497_), .A4(new_n499_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G113gat), .B(G141gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G169gat), .B(G197gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n508_), .B(new_n509_), .Z(new_n510_));
  NAND4_X1  g309(.A1(new_n501_), .A2(new_n505_), .A3(new_n507_), .A4(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT80), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n507_), .A2(new_n505_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n514_), .A2(KEYINPUT80), .A3(new_n501_), .A4(new_n510_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n501_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n510_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT81), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT82), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n476_), .A2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n524_), .B(KEYINPUT105), .Z(new_n525_));
  INV_X1    g324(.A(G106gat), .ZN(new_n526_));
  OR2_X1    g325(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n527_), .A2(KEYINPUT65), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT65), .B1(new_n527_), .B2(new_n528_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n526_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT66), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT10), .B(G99gat), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT65), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n529_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT66), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n537_), .A2(new_n538_), .A3(new_n526_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n533_), .A2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT68), .B1(G85gat), .B2(G92gat), .ZN(new_n541_));
  NAND3_X1  g340(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n542_), .ZN(new_n544_));
  XOR2_X1   g343(.A(KEYINPUT67), .B(G92gat), .Z(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(G85gat), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT9), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n544_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT68), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n543_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G99gat), .A2(G106gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT6), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n540_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G57gat), .B(G64gat), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n554_), .A2(KEYINPUT11), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(KEYINPUT11), .ZN(new_n556_));
  XOR2_X1   g355(.A(G71gat), .B(G78gat), .Z(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  OR2_X1    g357(.A1(new_n556_), .A2(new_n557_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G85gat), .B(G92gat), .ZN(new_n561_));
  NOR2_X1   g360(.A1(G99gat), .A2(G106gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT7), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n561_), .B1(new_n563_), .B2(new_n552_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT8), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT70), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT7), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n562_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT6), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n551_), .B(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT69), .B1(new_n568_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT69), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n563_), .A2(new_n572_), .A3(new_n552_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n561_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n571_), .A2(new_n573_), .A3(new_n565_), .A4(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n574_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT70), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n576_), .A2(new_n577_), .A3(KEYINPUT8), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n566_), .A2(new_n575_), .A3(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n553_), .A2(new_n560_), .A3(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT71), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n560_), .B1(new_n553_), .B2(new_n579_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n553_), .A2(KEYINPUT71), .A3(new_n579_), .A4(new_n560_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n582_), .A2(new_n584_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G230gat), .A2(G233gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n587_), .B(KEYINPUT64), .Z(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(KEYINPUT72), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n583_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n553_), .A2(new_n579_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n560_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n594_), .A2(new_n595_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n580_), .A2(new_n588_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n593_), .A2(new_n598_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n590_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G120gat), .B(G148gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT5), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G176gat), .B(G204gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n604_), .B(new_n605_), .Z(new_n606_));
  NAND2_X1  g405(.A1(new_n602_), .A2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n583_), .A2(new_n592_), .ZN(new_n608_));
  AOI211_X1 g407(.A(new_n560_), .B(new_n596_), .C1(new_n553_), .C2(new_n579_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  AOI22_X1  g409(.A1(new_n610_), .A2(new_n600_), .B1(new_n586_), .B2(new_n589_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n606_), .ZN(new_n612_));
  AOI21_X1  g411(.A(KEYINPUT73), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  AND4_X1   g412(.A1(KEYINPUT73), .A2(new_n590_), .A3(new_n601_), .A4(new_n612_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n607_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT13), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT74), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n615_), .B(KEYINPUT13), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(KEYINPUT74), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G190gat), .B(G218gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT36), .Z(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n494_), .A2(new_n495_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n594_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G232gat), .A2(G233gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT34), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT35), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n553_), .A2(new_n498_), .A3(new_n579_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n629_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n632_), .A2(new_n633_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n637_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n629_), .A2(new_n639_), .A3(new_n634_), .A4(new_n635_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n627_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n625_), .A2(KEYINPUT36), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n638_), .A2(new_n642_), .A3(new_n640_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT76), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT76), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n638_), .A2(new_n640_), .A3(new_n645_), .A4(new_n642_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n641_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT37), .ZN(new_n648_));
  NAND2_X1  g447(.A1(G231gat), .A2(G233gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n486_), .B(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(new_n560_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G127gat), .B(G155gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT16), .ZN(new_n653_));
  XOR2_X1   g452(.A(G183gat), .B(G211gat), .Z(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT17), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n655_), .A2(new_n656_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n651_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(KEYINPUT77), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT77), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n662_), .B1(new_n651_), .B2(new_n658_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n661_), .B1(new_n660_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n648_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n622_), .A2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT78), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n525_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n435_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n670_), .A2(new_n479_), .A3(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT38), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n622_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n522_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n675_), .A2(new_n676_), .A3(new_n665_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n476_), .A2(new_n647_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI21_X1  g478(.A(G1gat), .B1(new_n679_), .B2(new_n435_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n672_), .A2(new_n673_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n674_), .A2(new_n680_), .A3(new_n681_), .ZN(G1324gat));
  OAI21_X1  g481(.A(G8gat), .B1(new_n679_), .B2(new_n469_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n683_), .A2(KEYINPUT39), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(KEYINPUT39), .ZN(new_n685_));
  INV_X1    g484(.A(new_n469_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(new_n480_), .ZN(new_n687_));
  OAI22_X1  g486(.A1(new_n684_), .A2(new_n685_), .B1(new_n669_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT40), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(G1325gat));
  OAI21_X1  g489(.A(G15gat), .B1(new_n679_), .B2(new_n462_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT41), .Z(new_n692_));
  INV_X1    g491(.A(new_n462_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n670_), .A2(new_n445_), .A3(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1326gat));
  XNOR2_X1  g494(.A(new_n473_), .B(KEYINPUT106), .ZN(new_n696_));
  OAI21_X1  g495(.A(G22gat), .B1(new_n679_), .B2(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n697_), .A2(KEYINPUT42), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n697_), .A2(KEYINPUT42), .ZN(new_n699_));
  OR2_X1    g498(.A1(new_n696_), .A2(G22gat), .ZN(new_n700_));
  OAI22_X1  g499(.A1(new_n698_), .A2(new_n699_), .B1(new_n669_), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT107), .ZN(G1327gat));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n442_), .A2(new_n438_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT101), .B1(new_n473_), .B2(new_n441_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n462_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n472_), .A2(new_n475_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n648_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT109), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT37), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n647_), .B(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT109), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n715_), .A3(new_n709_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT108), .B1(new_n714_), .B2(new_n709_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n718_), .B(KEYINPUT43), .C1(new_n476_), .C2(new_n713_), .ZN(new_n719_));
  AOI22_X1  g518(.A1(new_n711_), .A2(new_n716_), .B1(new_n717_), .B2(new_n719_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n675_), .A2(new_n676_), .A3(new_n664_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n703_), .B1(new_n720_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n708_), .A2(new_n648_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n718_), .B1(new_n724_), .B2(KEYINPUT43), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n714_), .A2(KEYINPUT108), .A3(new_n709_), .ZN(new_n726_));
  NOR4_X1   g525(.A1(new_n476_), .A2(KEYINPUT109), .A3(KEYINPUT43), .A4(new_n713_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n715_), .B1(new_n714_), .B2(new_n709_), .ZN(new_n728_));
  OAI22_X1  g527(.A1(new_n725_), .A2(new_n726_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(KEYINPUT44), .A3(new_n721_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n723_), .A2(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n671_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G29gat), .ZN(new_n733_));
  INV_X1    g532(.A(new_n647_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n734_), .A2(new_n664_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n622_), .A2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n525_), .A2(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n435_), .A2(G29gat), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT110), .Z(new_n739_));
  OAI21_X1  g538(.A(new_n733_), .B1(new_n737_), .B2(new_n739_), .ZN(G1328gat));
  NAND3_X1  g539(.A1(new_n723_), .A2(new_n730_), .A3(new_n686_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G36gat), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n469_), .A2(G36gat), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n525_), .A2(new_n736_), .A3(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT45), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n525_), .A2(new_n746_), .A3(new_n736_), .A4(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n742_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT46), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n742_), .A2(new_n748_), .A3(KEYINPUT46), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1329gat));
  NOR2_X1   g552(.A1(new_n462_), .A2(new_n450_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n723_), .A2(new_n730_), .A3(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT111), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n723_), .A2(new_n730_), .A3(KEYINPUT111), .A4(new_n754_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n450_), .B1(new_n737_), .B2(new_n462_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT47), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n757_), .A2(new_n762_), .A3(new_n758_), .A4(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1330gat));
  INV_X1    g563(.A(G50gat), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n473_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n696_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n525_), .A2(new_n767_), .A3(new_n736_), .ZN(new_n768_));
  AOI22_X1  g567(.A1(new_n731_), .A2(new_n766_), .B1(new_n765_), .B2(new_n768_), .ZN(G1331gat));
  NOR3_X1   g568(.A1(new_n622_), .A2(new_n476_), .A3(new_n522_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n666_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT112), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n772_), .A2(G57gat), .A3(new_n435_), .ZN(new_n773_));
  INV_X1    g572(.A(G57gat), .ZN(new_n774_));
  AND4_X1   g573(.A1(new_n523_), .A2(new_n678_), .A3(new_n675_), .A4(new_n664_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n775_), .B2(new_n671_), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n773_), .A2(new_n776_), .ZN(G1332gat));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n686_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(G64gat), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(KEYINPUT48), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n779_), .A2(KEYINPUT48), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n469_), .A2(G64gat), .ZN(new_n782_));
  OAI22_X1  g581(.A1(new_n780_), .A2(new_n781_), .B1(new_n772_), .B2(new_n782_), .ZN(G1333gat));
  NAND2_X1  g582(.A1(new_n775_), .A2(new_n693_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(G71gat), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n785_), .A2(KEYINPUT49), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(KEYINPUT49), .ZN(new_n787_));
  OR2_X1    g586(.A1(new_n462_), .A2(G71gat), .ZN(new_n788_));
  OAI22_X1  g587(.A1(new_n786_), .A2(new_n787_), .B1(new_n772_), .B2(new_n788_), .ZN(G1334gat));
  NAND2_X1  g588(.A1(new_n775_), .A2(new_n767_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(G78gat), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n791_), .A2(KEYINPUT50), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(KEYINPUT50), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n696_), .A2(G78gat), .ZN(new_n794_));
  OAI22_X1  g593(.A1(new_n792_), .A2(new_n793_), .B1(new_n772_), .B2(new_n794_), .ZN(G1335gat));
  NAND2_X1  g594(.A1(new_n770_), .A2(new_n735_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(G85gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(new_n671_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT113), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n622_), .A2(new_n522_), .A3(new_n664_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n720_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n729_), .A2(KEYINPUT113), .A3(new_n801_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n435_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n799_), .B1(new_n805_), .B2(new_n798_), .ZN(G1336gat));
  AOI21_X1  g605(.A(G92gat), .B1(new_n797_), .B2(new_n686_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n803_), .A2(new_n804_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n686_), .A2(new_n545_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n808_), .B2(new_n809_), .ZN(G1337gat));
  NAND3_X1  g609(.A1(new_n797_), .A2(new_n693_), .A3(new_n537_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n811_), .B(KEYINPUT114), .ZN(new_n812_));
  INV_X1    g611(.A(G99gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n462_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT51), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n812_), .B(new_n817_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1338gat));
  XNOR2_X1  g618(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n720_), .A2(new_n473_), .A3(new_n802_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT52), .B1(new_n821_), .B2(new_n526_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n729_), .A2(new_n288_), .A3(new_n801_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(G106gat), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n796_), .A2(G106gat), .A3(new_n473_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n820_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n820_), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n830_), .B(new_n827_), .C1(new_n822_), .C2(new_n825_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n829_), .A2(new_n831_), .ZN(G1339gat));
  INV_X1    g631(.A(KEYINPUT57), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n611_), .A2(KEYINPUT73), .A3(new_n612_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n590_), .A2(new_n601_), .A3(new_n612_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT73), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n598_), .B1(new_n583_), .B2(new_n592_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n582_), .A2(new_n585_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n589_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n839_), .B2(new_n599_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n593_), .A2(new_n600_), .A3(KEYINPUT55), .A4(new_n598_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n841_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  AND3_X1   g644(.A1(new_n845_), .A2(KEYINPUT56), .A3(new_n606_), .ZN(new_n846_));
  AOI21_X1  g645(.A(KEYINPUT56), .B1(new_n845_), .B2(new_n606_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n522_), .B(new_n838_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n503_), .A2(new_n497_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n496_), .A2(new_n504_), .A3(new_n499_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n851_), .A3(new_n518_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n849_), .B1(new_n516_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n516_), .A2(new_n849_), .A3(new_n852_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n615_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n848_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n833_), .B1(new_n858_), .B2(new_n734_), .ZN(new_n859_));
  AOI211_X1 g658(.A(KEYINPUT57), .B(new_n647_), .C1(new_n848_), .C2(new_n857_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n855_), .ZN(new_n861_));
  OAI22_X1  g660(.A1(new_n613_), .A2(new_n614_), .B1(new_n861_), .B2(new_n853_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT117), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n845_), .A2(new_n606_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT56), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n845_), .A2(KEYINPUT56), .A3(new_n606_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n838_), .A2(new_n856_), .A3(new_n869_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n863_), .A2(new_n868_), .A3(KEYINPUT58), .A4(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n648_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n837_), .A2(new_n834_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n873_), .A2(new_n869_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT58), .B1(new_n874_), .B2(new_n863_), .ZN(new_n875_));
  OAI22_X1  g674(.A1(new_n859_), .A2(new_n860_), .B1(new_n872_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT118), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n868_), .A2(new_n870_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n873_), .A2(new_n869_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(new_n648_), .A3(new_n871_), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n883_), .B(KEYINPUT118), .C1(new_n859_), .C2(new_n860_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n878_), .A2(new_n665_), .A3(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n620_), .A2(new_n523_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n713_), .A2(new_n664_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT54), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n666_), .A2(new_n620_), .A3(new_n889_), .A4(new_n523_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n885_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n885_), .A2(KEYINPUT119), .A3(new_n891_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n686_), .A2(new_n288_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n693_), .A3(new_n671_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n894_), .A2(new_n895_), .A3(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n900_), .A2(new_n372_), .A3(new_n522_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n876_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n891_), .B1(new_n902_), .B2(new_n664_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n903_), .A2(new_n898_), .A3(new_n904_), .ZN(new_n905_));
  AOI211_X1 g704(.A(new_n523_), .B(new_n905_), .C1(new_n899_), .C2(KEYINPUT59), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n901_), .B1(new_n906_), .B2(new_n372_), .ZN(G1340gat));
  AOI211_X1 g706(.A(new_n622_), .B(new_n905_), .C1(new_n899_), .C2(KEYINPUT59), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n374_), .B1(new_n622_), .B2(KEYINPUT60), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n909_), .B1(KEYINPUT60), .B2(new_n374_), .ZN(new_n910_));
  OAI22_X1  g709(.A1(new_n908_), .A2(new_n374_), .B1(new_n899_), .B2(new_n910_), .ZN(G1341gat));
  NAND3_X1  g710(.A1(new_n900_), .A2(new_n369_), .A3(new_n664_), .ZN(new_n912_));
  AOI211_X1 g711(.A(new_n665_), .B(new_n905_), .C1(new_n899_), .C2(KEYINPUT59), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n369_), .ZN(G1342gat));
  AOI21_X1  g713(.A(G134gat), .B1(new_n900_), .B2(new_n647_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n905_), .B1(new_n899_), .B2(KEYINPUT59), .ZN(new_n916_));
  XOR2_X1   g715(.A(KEYINPUT121), .B(G134gat), .Z(new_n917_));
  NOR2_X1   g716(.A1(new_n713_), .A2(new_n917_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n915_), .B1(new_n916_), .B2(new_n918_), .ZN(G1343gat));
  AND2_X1   g718(.A1(new_n888_), .A2(new_n890_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n664_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n921_));
  AOI211_X1 g720(.A(new_n893_), .B(new_n920_), .C1(new_n921_), .C2(new_n884_), .ZN(new_n922_));
  AOI21_X1  g721(.A(KEYINPUT119), .B1(new_n885_), .B2(new_n891_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND4_X1  g723(.A1(new_n288_), .A2(new_n469_), .A3(new_n462_), .A4(new_n671_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT122), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n924_), .A2(new_n522_), .A3(new_n926_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(new_n927_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g727(.A1(new_n924_), .A2(new_n675_), .A3(new_n926_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g729(.A1(new_n894_), .A2(new_n664_), .A3(new_n895_), .A4(new_n926_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(KEYINPUT123), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n933_));
  NAND4_X1  g732(.A1(new_n924_), .A2(new_n933_), .A3(new_n664_), .A4(new_n926_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(KEYINPUT61), .B(G155gat), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n932_), .A2(new_n934_), .A3(new_n935_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n932_), .B2(new_n934_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1346gat));
  NAND2_X1  g737(.A1(new_n924_), .A2(new_n926_), .ZN(new_n939_));
  OAI21_X1  g738(.A(G162gat), .B1(new_n939_), .B2(new_n713_), .ZN(new_n940_));
  OR2_X1    g739(.A1(new_n734_), .A2(G162gat), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n939_), .B2(new_n941_), .ZN(G1347gat));
  NAND2_X1  g741(.A1(new_n686_), .A2(new_n470_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n943_), .ZN(new_n944_));
  NAND3_X1  g743(.A1(new_n903_), .A2(new_n696_), .A3(new_n944_), .ZN(new_n945_));
  INV_X1    g744(.A(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n304_), .B1(new_n946_), .B2(new_n522_), .ZN(new_n947_));
  OR2_X1    g746(.A1(new_n947_), .A2(KEYINPUT124), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(KEYINPUT124), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n948_), .A2(KEYINPUT62), .A3(new_n949_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n947_), .A2(KEYINPUT124), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT62), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n945_), .A2(new_n676_), .ZN(new_n953_));
  AOI22_X1  g752(.A1(new_n951_), .A2(new_n952_), .B1(new_n313_), .B2(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n950_), .A2(new_n954_), .ZN(G1348gat));
  AOI21_X1  g754(.A(G176gat), .B1(new_n946_), .B2(new_n675_), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n894_), .A2(new_n473_), .A3(new_n895_), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n957_), .B(new_n958_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n622_), .A2(new_n305_), .A3(new_n943_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n956_), .B1(new_n959_), .B2(new_n960_), .ZN(G1349gat));
  NOR3_X1   g760(.A1(new_n943_), .A2(new_n302_), .A3(new_n665_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n903_), .A2(new_n696_), .A3(new_n962_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(KEYINPUT126), .ZN(new_n964_));
  NOR2_X1   g763(.A1(new_n943_), .A2(new_n665_), .ZN(new_n965_));
  AOI21_X1  g764(.A(KEYINPUT125), .B1(new_n924_), .B2(new_n473_), .ZN(new_n966_));
  NOR4_X1   g765(.A1(new_n922_), .A2(new_n923_), .A3(new_n958_), .A4(new_n288_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n965_), .B1(new_n966_), .B2(new_n967_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n330_), .A2(new_n332_), .ZN(new_n969_));
  INV_X1    g768(.A(new_n969_), .ZN(new_n970_));
  AOI21_X1  g769(.A(new_n964_), .B1(new_n968_), .B2(new_n970_), .ZN(G1350gat));
  OAI21_X1  g770(.A(G190gat), .B1(new_n945_), .B2(new_n713_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n647_), .A2(new_n301_), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n972_), .B1(new_n945_), .B2(new_n973_), .ZN(G1351gat));
  NAND2_X1  g773(.A1(new_n288_), .A2(new_n435_), .ZN(new_n975_));
  NOR3_X1   g774(.A1(new_n975_), .A2(new_n693_), .A3(new_n469_), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n924_), .A2(new_n522_), .A3(new_n976_), .ZN(new_n977_));
  XNOR2_X1  g776(.A(new_n977_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g777(.A1(new_n894_), .A2(new_n895_), .ZN(new_n979_));
  INV_X1    g778(.A(new_n976_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(new_n979_), .A2(new_n980_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n981_), .A2(new_n675_), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n982_), .B1(KEYINPUT127), .B2(G204gat), .ZN(new_n983_));
  XNOR2_X1  g782(.A(KEYINPUT127), .B(G204gat), .ZN(new_n984_));
  NAND3_X1  g783(.A1(new_n981_), .A2(new_n675_), .A3(new_n984_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n983_), .A2(new_n985_), .ZN(G1353gat));
  NAND2_X1  g785(.A1(new_n981_), .A2(new_n664_), .ZN(new_n987_));
  OAI21_X1  g786(.A(new_n987_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n988_));
  XNOR2_X1  g787(.A(KEYINPUT63), .B(G211gat), .ZN(new_n989_));
  NAND3_X1  g788(.A1(new_n981_), .A2(new_n664_), .A3(new_n989_), .ZN(new_n990_));
  NAND2_X1  g789(.A1(new_n988_), .A2(new_n990_), .ZN(G1354gat));
  NAND3_X1  g790(.A1(new_n981_), .A2(new_n239_), .A3(new_n647_), .ZN(new_n992_));
  NOR3_X1   g791(.A1(new_n979_), .A2(new_n713_), .A3(new_n980_), .ZN(new_n993_));
  OAI21_X1  g792(.A(new_n992_), .B1(new_n239_), .B2(new_n993_), .ZN(G1355gat));
endmodule


