//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 1 1 1 1 1 0 0 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_;
  XNOR2_X1  g000(.A(G71gat), .B(G99gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT93), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G15gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G227gat), .A2(G233gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(KEYINPUT31), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(G169gat), .ZN(new_n210_));
  INV_X1    g009(.A(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(G190gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT23), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT90), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n213_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  OAI211_X1 g016(.A(KEYINPUT90), .B(KEYINPUT23), .C1(new_n211_), .C2(new_n212_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n210_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(G190gat), .B1(KEYINPUT87), .B2(KEYINPUT26), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT87), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT26), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n223_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT86), .B1(new_n225_), .B2(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT86), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n228_), .A2(new_n212_), .A3(KEYINPUT26), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n227_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT85), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT25), .B1(new_n231_), .B2(new_n211_), .ZN(new_n232_));
  OR3_X1    g031(.A1(new_n231_), .A2(new_n211_), .A3(KEYINPUT25), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n226_), .A2(new_n230_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT88), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G169gat), .ZN(new_n238_));
  INV_X1    g037(.A(G176gat), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n237_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n234_), .A2(new_n235_), .A3(new_n240_), .ZN(new_n241_));
  OR4_X1    g040(.A1(KEYINPUT89), .A2(new_n211_), .A3(new_n212_), .A4(KEYINPUT23), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n213_), .A2(new_n215_), .A3(KEYINPUT89), .ZN(new_n243_));
  OR3_X1    g042(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n241_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n235_), .B1(new_n234_), .B2(new_n240_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n221_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT91), .B(KEYINPUT30), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT92), .B(G43gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(KEYINPUT94), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n234_), .A2(new_n240_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT88), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(new_n241_), .A3(new_n245_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(new_n221_), .A3(new_n249_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n251_), .A2(new_n254_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n254_), .B1(new_n251_), .B2(new_n258_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G127gat), .B(G134gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT95), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G113gat), .B(G120gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT95), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n262_), .B(new_n267_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n268_), .A2(new_n264_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n266_), .A2(new_n269_), .ZN(new_n270_));
  NOR3_X1   g069(.A1(new_n260_), .A2(new_n261_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n251_), .A2(new_n258_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n253_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n272_), .B1(new_n274_), .B2(new_n259_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n208_), .B1(new_n271_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n270_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n274_), .A2(new_n272_), .A3(new_n259_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n207_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n268_), .A2(new_n264_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n263_), .A2(new_n265_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G141gat), .A2(G148gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT96), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT96), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n285_), .A2(G141gat), .A3(G148gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT2), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT3), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT3), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n288_), .A2(new_n291_), .A3(new_n293_), .A4(new_n294_), .ZN(new_n295_));
  OR2_X1    g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G155gat), .A2(G162gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT97), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n296_), .A2(KEYINPUT97), .A3(new_n297_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n295_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n298_), .A2(KEYINPUT1), .ZN(new_n303_));
  NAND3_X1  g102(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n304_));
  AND4_X1   g103(.A1(new_n284_), .A2(new_n290_), .A3(new_n286_), .A4(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n281_), .B(new_n282_), .C1(new_n302_), .C2(new_n307_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n300_), .A2(new_n301_), .ZN(new_n309_));
  AOI22_X1  g108(.A1(new_n309_), .A2(new_n295_), .B1(new_n303_), .B2(new_n305_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n310_), .B1(new_n266_), .B2(new_n269_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n308_), .A2(new_n311_), .A3(KEYINPUT4), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT4), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n270_), .B(new_n313_), .C1(new_n307_), .C2(new_n302_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n308_), .A2(new_n311_), .A3(new_n315_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT102), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT102), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n308_), .A2(new_n311_), .A3(new_n320_), .A4(new_n315_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n317_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G1gat), .B(G29gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G85gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT0), .B(G57gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n326_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n317_), .A2(new_n319_), .A3(new_n328_), .A4(new_n321_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G228gat), .A2(G233gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n309_), .A2(new_n295_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n335_), .B2(new_n306_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G211gat), .B(G218gat), .ZN(new_n337_));
  INV_X1    g136(.A(G204gat), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n338_), .A2(G197gat), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n337_), .B(KEYINPUT21), .C1(KEYINPUT99), .C2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G197gat), .B(G204gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n337_), .A2(KEYINPUT21), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n344_), .A2(new_n341_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n343_), .B1(new_n340_), .B2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n333_), .B1(new_n336_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n340_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n348_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n349_), .B(new_n332_), .C1(new_n334_), .C2(new_n310_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G78gat), .B(G106gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n352_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n347_), .A2(new_n350_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n310_), .A2(new_n334_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT98), .B(KEYINPUT28), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n357_), .B(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n354_), .B1(new_n347_), .B2(new_n350_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n361_), .B1(new_n362_), .B2(KEYINPUT100), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n356_), .A2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n353_), .A2(KEYINPUT100), .A3(new_n361_), .A4(new_n355_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n280_), .A2(new_n331_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT20), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n242_), .B(new_n243_), .C1(G183gat), .C2(G190gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n210_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT25), .B(G183gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT26), .B(G190gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  AND3_X1   g172(.A1(new_n373_), .A2(new_n240_), .A3(new_n244_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n219_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT101), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n373_), .A2(new_n240_), .A3(new_n244_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT101), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n219_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n370_), .B1(new_n376_), .B2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n368_), .B1(new_n380_), .B2(new_n349_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT19), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n257_), .A2(new_n221_), .A3(new_n346_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n381_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT104), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n381_), .A2(KEYINPUT104), .A3(new_n384_), .A4(new_n385_), .ZN(new_n389_));
  OAI211_X1 g188(.A(new_n346_), .B(new_n370_), .C1(new_n219_), .C2(new_n377_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT103), .B(KEYINPUT20), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n346_), .B1(new_n257_), .B2(new_n221_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n383_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n388_), .A2(new_n389_), .A3(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G8gat), .B(G36gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT18), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G64gat), .B(G92gat), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n397_), .B(new_n398_), .Z(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n395_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT27), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n384_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n384_), .A2(KEYINPUT20), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n374_), .A2(KEYINPUT101), .A3(new_n375_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n378_), .B1(new_n377_), .B2(new_n219_), .ZN(new_n406_));
  AOI22_X1  g205(.A1(new_n405_), .A2(new_n406_), .B1(new_n210_), .B2(new_n369_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n407_), .B2(new_n346_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n248_), .A2(new_n349_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n403_), .A2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n402_), .B1(new_n411_), .B2(new_n399_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n401_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n403_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n408_), .A2(new_n409_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n399_), .A3(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n400_), .B1(new_n403_), .B2(new_n410_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT105), .B(KEYINPUT27), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n413_), .A2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n367_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n399_), .A2(KEYINPUT32), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n395_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n411_), .A2(new_n423_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n330_), .A3(new_n426_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n312_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n308_), .A2(new_n311_), .A3(new_n316_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n326_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT33), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n329_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n319_), .A2(new_n321_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n433_), .A2(KEYINPUT33), .A3(new_n328_), .A4(new_n317_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n432_), .A2(new_n434_), .A3(new_n416_), .A4(new_n417_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n427_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n366_), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n401_), .A2(new_n412_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n366_), .A2(new_n330_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n280_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n422_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  XOR2_X1   g242(.A(KEYINPUT10), .B(G99gat), .Z(new_n444_));
  INV_X1    g243(.A(G106gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G99gat), .A2(G106gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT6), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT6), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(G99gat), .A3(G106gat), .ZN(new_n450_));
  AND2_X1   g249(.A1(G85gat), .A2(G92gat), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT9), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n448_), .A2(new_n450_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(G85gat), .A2(G92gat), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT9), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n446_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(new_n451_), .A2(new_n454_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n448_), .A2(new_n450_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n459_), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT8), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT65), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n448_), .A2(new_n450_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT7), .ZN(new_n469_));
  INV_X1    g268(.A(G99gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n445_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(new_n460_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n455_), .B1(new_n468_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT65), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(KEYINPUT8), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n467_), .A2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n466_), .B(new_n455_), .C1(new_n468_), .C2(new_n472_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT64), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n463_), .A2(new_n464_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT64), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n479_), .A2(new_n480_), .A3(new_n466_), .A4(new_n455_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n478_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n458_), .B1(new_n476_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G29gat), .B(G36gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G43gat), .B(G50gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(KEYINPUT15), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n467_), .A2(new_n475_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n457_), .B(KEYINPUT68), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n488_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G232gat), .A2(G233gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT74), .ZN(new_n493_));
  XNOR2_X1  g292(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT35), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n487_), .A2(new_n491_), .A3(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n495_), .A2(new_n496_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n498_), .A2(new_n499_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G190gat), .B(G218gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT75), .ZN(new_n505_));
  XOR2_X1   g304(.A(G134gat), .B(G162gat), .Z(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT36), .ZN(new_n508_));
  AND2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n503_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT37), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n507_), .B(new_n508_), .ZN(new_n512_));
  OAI211_X1 g311(.A(new_n510_), .B(new_n511_), .C1(new_n503_), .C2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n502_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n514_), .A2(new_n509_), .A3(new_n500_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n512_), .B1(new_n514_), .B2(new_n500_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT37), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(KEYINPUT76), .B(G8gat), .Z(new_n520_));
  INV_X1    g319(.A(G1gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT14), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G15gat), .B(G22gat), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G1gat), .B(G8gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n522_), .A2(new_n523_), .A3(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G231gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT77), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n529_), .B(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(G64gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(G57gat), .ZN(new_n534_));
  INV_X1    g333(.A(G57gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(G64gat), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT66), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n534_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n537_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT11), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n534_), .A2(new_n536_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT66), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT11), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(new_n538_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G71gat), .B(G78gat), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n541_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  OAI211_X1 g347(.A(KEYINPUT11), .B(new_n546_), .C1(new_n539_), .C2(new_n540_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n532_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n532_), .A2(new_n550_), .ZN(new_n552_));
  XOR2_X1   g351(.A(G127gat), .B(G155gat), .Z(new_n553_));
  XNOR2_X1  g352(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G183gat), .B(G211gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  AOI22_X1  g356(.A1(new_n551_), .A2(new_n552_), .B1(KEYINPUT17), .B2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(KEYINPUT17), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n551_), .A2(new_n552_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n558_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n519_), .A2(KEYINPUT79), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT79), .ZN(new_n563_));
  INV_X1    g362(.A(new_n561_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n563_), .B1(new_n518_), .B2(new_n564_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n443_), .A2(new_n562_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n529_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n486_), .B(KEYINPUT80), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT80), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n486_), .B(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n529_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(G229gat), .A3(G233gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n567_), .A2(new_n488_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G229gat), .A2(G233gat), .ZN(new_n576_));
  XOR2_X1   g375(.A(new_n576_), .B(KEYINPUT81), .Z(new_n577_));
  NAND3_X1  g376(.A1(new_n575_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n574_), .A2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G113gat), .B(G141gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(new_n580_), .B(KEYINPUT82), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n581_), .B(KEYINPUT83), .Z(new_n582_));
  XNOR2_X1  g381(.A(G169gat), .B(G197gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n579_), .A2(KEYINPUT84), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n585_), .B1(new_n579_), .B2(KEYINPUT84), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT72), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G230gat), .A2(G233gat), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT67), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n483_), .B2(new_n550_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n476_), .A2(new_n482_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n550_), .A3(new_n457_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n483_), .A2(new_n592_), .A3(new_n550_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n591_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n599_));
  OAI21_X1  g398(.A(new_n599_), .B1(new_n483_), .B2(new_n550_), .ZN(new_n600_));
  AND3_X1   g399(.A1(new_n548_), .A2(KEYINPUT12), .A3(new_n549_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n601_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n600_), .A2(new_n590_), .A3(new_n602_), .A4(new_n595_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G120gat), .B(G148gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT5), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G176gat), .B(G204gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n598_), .A2(new_n603_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT71), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n598_), .A2(KEYINPUT71), .A3(new_n603_), .A4(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n598_), .A2(new_n603_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n607_), .B(KEYINPUT70), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n612_), .A2(KEYINPUT13), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT13), .B1(new_n612_), .B2(new_n615_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n589_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n612_), .A2(new_n615_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT13), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(KEYINPUT72), .A3(new_n616_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n619_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n566_), .A2(new_n588_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(new_n521_), .A3(new_n330_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT38), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT107), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n622_), .A2(new_n616_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n588_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n443_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n515_), .A2(new_n516_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(new_n561_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT106), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n330_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n630_), .B1(new_n638_), .B2(G1gat), .ZN(new_n639_));
  AOI211_X1 g438(.A(KEYINPUT107), .B(new_n521_), .C1(new_n637_), .C2(new_n330_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n629_), .B1(new_n639_), .B2(new_n640_), .ZN(G1324gat));
  OAI21_X1  g440(.A(G8gat), .B1(new_n636_), .B2(new_n438_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT39), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n421_), .A2(new_n520_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT108), .B1(new_n627_), .B2(new_n645_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n627_), .A2(KEYINPUT108), .A3(new_n645_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n643_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT40), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n643_), .B(KEYINPUT40), .C1(new_n646_), .C2(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1325gat));
  OR3_X1    g451(.A1(new_n626_), .A2(G15gat), .A3(new_n442_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n637_), .A2(new_n280_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n654_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(KEYINPUT41), .B1(new_n654_), .B2(G15gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(G1326gat));
  OR3_X1    g456(.A1(new_n626_), .A2(G22gat), .A3(new_n366_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n366_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n637_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n660_), .A2(new_n661_), .A3(G22gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n660_), .B2(G22gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n658_), .B1(new_n662_), .B2(new_n663_), .ZN(G1327gat));
  INV_X1    g463(.A(new_n634_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(new_n564_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n633_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G29gat), .B1(new_n668_), .B2(new_n330_), .ZN(new_n669_));
  NOR3_X1   g468(.A1(new_n631_), .A2(new_n632_), .A3(new_n564_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n439_), .A2(new_n413_), .A3(new_n420_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n659_), .B1(new_n427_), .B2(new_n435_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n442_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n438_), .A2(new_n331_), .A3(new_n280_), .A4(new_n366_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n671_), .B1(new_n676_), .B2(new_n519_), .ZN(new_n677_));
  AOI211_X1 g476(.A(KEYINPUT43), .B(new_n518_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n670_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI211_X1 g480(.A(KEYINPUT44), .B(new_n670_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n330_), .A2(G29gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n669_), .B1(new_n684_), .B2(new_n685_), .ZN(G1328gat));
  NOR2_X1   g485(.A1(new_n631_), .A2(new_n632_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n438_), .A2(G36gat), .ZN(new_n688_));
  NAND4_X1  g487(.A1(new_n687_), .A2(new_n676_), .A3(new_n666_), .A4(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT110), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT45), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n681_), .A2(new_n421_), .A3(new_n682_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT109), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(G36gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n692_), .B2(G36gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n691_), .B(KEYINPUT46), .C1(new_n694_), .C2(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1329gat));
  XNOR2_X1  g499(.A(KEYINPUT111), .B(G43gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n701_), .B1(new_n667_), .B2(new_n442_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n280_), .A2(G43gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n683_), .B2(new_n703_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g504(.A(G50gat), .B1(new_n683_), .B2(new_n366_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n366_), .A2(G50gat), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT112), .Z(new_n708_));
  OAI21_X1  g507(.A(new_n706_), .B1(new_n667_), .B2(new_n708_), .ZN(G1331gat));
  AND3_X1   g508(.A1(new_n566_), .A2(new_n631_), .A3(new_n632_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n710_), .A2(new_n535_), .A3(new_n330_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n588_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n624_), .A2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n635_), .ZN(new_n714_));
  OAI21_X1  g513(.A(G57gat), .B1(new_n714_), .B2(new_n331_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n711_), .A2(new_n715_), .ZN(G1332gat));
  OAI21_X1  g515(.A(G64gat), .B1(new_n714_), .B2(new_n438_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n710_), .A2(new_n533_), .A3(new_n421_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(G1333gat));
  OAI21_X1  g520(.A(G71gat), .B1(new_n714_), .B2(new_n442_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT49), .ZN(new_n723_));
  INV_X1    g522(.A(G71gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n710_), .A2(new_n724_), .A3(new_n280_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1334gat));
  INV_X1    g525(.A(G78gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n710_), .A2(new_n727_), .A3(new_n659_), .ZN(new_n728_));
  OAI21_X1  g527(.A(G78gat), .B1(new_n714_), .B2(new_n366_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(KEYINPUT50), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(KEYINPUT50), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n728_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT114), .ZN(G1335gat));
  NAND3_X1  g532(.A1(new_n631_), .A2(new_n632_), .A3(new_n561_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT43), .B1(new_n443_), .B2(new_n518_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n676_), .A2(new_n671_), .A3(new_n519_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n331_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n624_), .A2(new_n666_), .A3(new_n712_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT115), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n624_), .A2(new_n712_), .A3(KEYINPUT115), .A4(new_n666_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n331_), .A2(G85gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n739_), .B1(new_n745_), .B2(new_n746_), .ZN(G1336gat));
  OAI21_X1  g546(.A(G92gat), .B1(new_n738_), .B2(new_n438_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n438_), .A2(G92gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n748_), .B1(new_n745_), .B2(new_n749_), .ZN(G1337gat));
  OAI21_X1  g549(.A(G99gat), .B1(new_n738_), .B2(new_n442_), .ZN(new_n751_));
  XOR2_X1   g550(.A(KEYINPUT117), .B(KEYINPUT51), .Z(new_n752_));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n280_), .A2(new_n444_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n753_), .B1(new_n744_), .B2(new_n755_), .ZN(new_n756_));
  AOI211_X1 g555(.A(KEYINPUT116), .B(new_n754_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n751_), .B(new_n752_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n758_), .A2(KEYINPUT118), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n758_), .A2(KEYINPUT118), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n751_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT51), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n759_), .B1(new_n760_), .B2(new_n762_), .ZN(G1338gat));
  NAND3_X1  g562(.A1(new_n744_), .A2(new_n445_), .A3(new_n659_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT52), .ZN(new_n765_));
  INV_X1    g564(.A(new_n734_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n766_), .B(new_n659_), .C1(new_n677_), .C2(new_n678_), .ZN(new_n767_));
  OAI21_X1  g566(.A(G106gat), .B1(new_n767_), .B2(KEYINPUT119), .ZN(new_n768_));
  INV_X1    g567(.A(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(KEYINPUT119), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n765_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT119), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n737_), .B2(new_n659_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n768_), .A2(new_n773_), .A3(KEYINPUT52), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n764_), .B1(new_n771_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT53), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n777_), .B(new_n764_), .C1(new_n771_), .C2(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1339gat));
  INV_X1    g578(.A(new_n599_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n594_), .A2(new_n457_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n550_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n602_), .A2(new_n595_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n591_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT121), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT121), .B(new_n591_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n603_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n784_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n791_), .A2(KEYINPUT55), .A3(new_n590_), .A4(new_n600_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n787_), .A2(new_n788_), .A3(new_n790_), .A4(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n614_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT56), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n793_), .A2(new_n796_), .A3(new_n614_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n795_), .A2(new_n612_), .A3(new_n588_), .A4(new_n797_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n575_), .A2(new_n572_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n799_), .A2(new_n577_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n569_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n585_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n579_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(new_n585_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n620_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n798_), .A2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n665_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n794_), .A2(KEYINPUT56), .B1(new_n610_), .B2(new_n611_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(new_n804_), .A3(new_n797_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n810_), .A2(KEYINPUT58), .A3(new_n804_), .A4(new_n797_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n519_), .A3(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n806_), .A2(KEYINPUT57), .A3(new_n665_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n809_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n561_), .ZN(new_n818_));
  AOI211_X1 g617(.A(new_n588_), .B(new_n561_), .C1(new_n513_), .C2(new_n517_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(new_n622_), .A3(new_n616_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n631_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n821_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n819_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n818_), .A2(new_n827_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n442_), .A2(new_n421_), .A3(new_n659_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(new_n330_), .A3(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(G113gat), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n588_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n830_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n826_), .B1(new_n817_), .B2(new_n561_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n836_), .A2(new_n331_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(KEYINPUT59), .A3(new_n829_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n632_), .B1(new_n835_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n833_), .B1(new_n839_), .B2(new_n832_), .ZN(G1340gat));
  INV_X1    g639(.A(G120gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n823_), .B2(KEYINPUT60), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n831_), .B(new_n842_), .C1(KEYINPUT60), .C2(new_n841_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n625_), .B1(new_n835_), .B2(new_n838_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n841_), .ZN(G1341gat));
  INV_X1    g644(.A(G127gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n831_), .A2(new_n846_), .A3(new_n564_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n561_), .B1(new_n835_), .B2(new_n838_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n848_), .B2(new_n846_), .ZN(G1342gat));
  NAND3_X1  g648(.A1(new_n837_), .A2(new_n634_), .A3(new_n829_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n851_));
  INV_X1    g650(.A(G134gat), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(KEYINPUT123), .B(G134gat), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n519_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n855_), .B1(new_n835_), .B2(new_n838_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n851_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n853_), .A2(new_n856_), .A3(new_n857_), .ZN(G1343gat));
  NAND2_X1  g657(.A1(new_n442_), .A2(new_n659_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n421_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n837_), .A2(new_n588_), .A3(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g661(.A1(new_n837_), .A2(new_n624_), .A3(new_n860_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g663(.A1(new_n837_), .A2(new_n860_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n561_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT61), .B(G155gat), .Z(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1346gat));
  OAI21_X1  g667(.A(G162gat), .B1(new_n865_), .B2(new_n518_), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n665_), .A2(G162gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n865_), .B2(new_n870_), .ZN(G1347gat));
  INV_X1    g670(.A(new_n367_), .ZN(new_n872_));
  AOI21_X1  g671(.A(KEYINPUT57), .B1(new_n806_), .B2(new_n665_), .ZN(new_n873_));
  AOI211_X1 g672(.A(new_n808_), .B(new_n634_), .C1(new_n798_), .C2(new_n805_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n564_), .B1(new_n875_), .B2(new_n815_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n421_), .B(new_n872_), .C1(new_n876_), .C2(new_n826_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NAND4_X1  g678(.A1(new_n828_), .A2(KEYINPUT124), .A3(new_n421_), .A4(new_n872_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(KEYINPUT22), .B(G169gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n588_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  INV_X1    g683(.A(new_n877_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n588_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n886_), .B2(G169gat), .ZN(new_n887_));
  AOI211_X1 g686(.A(KEYINPUT62), .B(new_n238_), .C1(new_n885_), .C2(new_n588_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n883_), .B1(new_n887_), .B2(new_n888_), .ZN(G1348gat));
  INV_X1    g688(.A(KEYINPUT125), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n823_), .A2(G176gat), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n893_));
  OAI21_X1  g692(.A(G176gat), .B1(new_n877_), .B2(new_n625_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n890_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n438_), .B1(new_n818_), .B2(new_n827_), .ZN(new_n897_));
  AOI21_X1  g696(.A(KEYINPUT124), .B1(new_n897_), .B2(new_n872_), .ZN(new_n898_));
  NOR4_X1   g697(.A1(new_n836_), .A2(new_n878_), .A3(new_n438_), .A4(new_n367_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n891_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n900_), .A2(KEYINPUT125), .A3(new_n894_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n896_), .A2(new_n901_), .ZN(G1349gat));
  NOR2_X1   g701(.A1(new_n877_), .A2(new_n561_), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n903_), .A2(KEYINPUT126), .ZN(new_n904_));
  AOI21_X1  g703(.A(G183gat), .B1(new_n903_), .B2(KEYINPUT126), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n561_), .A2(new_n371_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n904_), .A2(new_n905_), .B1(new_n881_), .B2(new_n906_), .ZN(G1350gat));
  NAND3_X1  g706(.A1(new_n881_), .A2(new_n372_), .A3(new_n634_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n518_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n212_), .B2(new_n909_), .ZN(G1351gat));
  NOR2_X1   g709(.A1(new_n859_), .A2(new_n330_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  NOR3_X1   g711(.A1(new_n836_), .A2(new_n438_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n588_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g714(.A1(new_n913_), .A2(new_n624_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g716(.A1(new_n913_), .A2(new_n564_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n919_));
  AND2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n918_), .A2(new_n919_), .A3(new_n920_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n918_), .B2(new_n919_), .ZN(G1354gat));
  INV_X1    g721(.A(G218gat), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n913_), .A2(new_n923_), .A3(new_n634_), .ZN(new_n924_));
  NOR4_X1   g723(.A1(new_n836_), .A2(new_n438_), .A3(new_n518_), .A4(new_n912_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(new_n923_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n924_), .B(KEYINPUT127), .C1(new_n923_), .C2(new_n925_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1355gat));
endmodule


