//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n884_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n938_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT82), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT31), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT81), .ZN(new_n207_));
  INV_X1    g006(.A(G169gat), .ZN(new_n208_));
  OR3_X1    g007(.A1(new_n208_), .A2(KEYINPUT22), .A3(G176gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G183gat), .A2(G190gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n211_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n214_), .A2(new_n215_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT24), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n208_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(G183gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT25), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT25), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G183gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(KEYINPUT26), .B(G190gat), .Z(new_n228_));
  OAI211_X1 g027(.A(new_n219_), .B(new_n222_), .C1(new_n227_), .C2(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n230_));
  AND2_X1   g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT78), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT78), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n234_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n218_), .B1(new_n229_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT30), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n237_), .A2(new_n238_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n207_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n217_), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n219_), .A2(new_n242_), .B1(new_n210_), .B2(new_n209_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n236_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n222_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n227_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT26), .B(G190gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n245_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n243_), .B1(new_n244_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT30), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n237_), .A2(new_n238_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(KEYINPUT81), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(G227gat), .A2(G233gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT79), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G15gat), .B(G43gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G71gat), .B(G99gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT80), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n256_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n241_), .A2(new_n252_), .A3(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n259_), .A2(KEYINPUT81), .A3(new_n251_), .A4(new_n250_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n206_), .A2(new_n261_), .A3(KEYINPUT83), .A4(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(KEYINPUT83), .ZN(new_n264_));
  INV_X1    g063(.A(new_n206_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(KEYINPUT83), .B1(new_n261_), .B2(new_n262_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n263_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n204_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G155gat), .B(G162gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G141gat), .A2(G148gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT2), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT85), .A3(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n272_), .B1(new_n271_), .B2(KEYINPUT85), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NOR3_X1   g076(.A1(new_n274_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT84), .ZN(new_n279_));
  NOR2_X1   g078(.A1(G141gat), .A2(G148gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT3), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n279_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n280_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n270_), .B1(new_n278_), .B2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n270_), .A2(KEYINPUT1), .ZN(new_n287_));
  INV_X1    g086(.A(new_n280_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n288_), .A2(new_n271_), .A3(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n269_), .B1(new_n286_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n270_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n271_), .A2(KEYINPUT85), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT2), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(new_n273_), .A3(new_n276_), .ZN(new_n296_));
  NOR4_X1   g095(.A1(KEYINPUT84), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n297_), .A2(new_n282_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n293_), .B1(new_n296_), .B2(new_n298_), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n287_), .A2(new_n290_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n299_), .A2(new_n300_), .A3(new_n204_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n292_), .A2(KEYINPUT4), .A3(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G225gat), .A2(G233gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n204_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT4), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n292_), .A2(new_n301_), .A3(new_n303_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G1gat), .B(G29gat), .ZN(new_n309_));
  INV_X1    g108(.A(G85gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT0), .B(G57gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n307_), .A2(new_n308_), .A3(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n313_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n268_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT21), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT88), .ZN(new_n320_));
  INV_X1    g119(.A(G204gat), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n320_), .B1(new_n321_), .B2(G197gat), .ZN(new_n322_));
  AND2_X1   g121(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n323_));
  NOR2_X1   g122(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n322_), .B1(new_n325_), .B2(G197gat), .ZN(new_n326_));
  OR2_X1    g125(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n327_), .A2(KEYINPUT88), .A3(G197gat), .A4(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n319_), .B1(new_n326_), .B2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G211gat), .B(G218gat), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G197gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n325_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n319_), .B1(G197gat), .B2(G204gat), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n333_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n326_), .A2(new_n330_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n332_), .A2(new_n319_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n331_), .A2(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n342_));
  OAI21_X1  g141(.A(G106gat), .B1(new_n340_), .B2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G228gat), .A2(G233gat), .ZN(new_n344_));
  INV_X1    g143(.A(G78gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT29), .B1(new_n286_), .B2(new_n291_), .ZN(new_n347_));
  INV_X1    g146(.A(G106gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n327_), .A2(G197gat), .A3(new_n328_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n322_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n339_), .A3(new_n329_), .ZN(new_n352_));
  AOI21_X1  g151(.A(KEYINPUT21), .B1(new_n351_), .B2(new_n329_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT87), .B(G204gat), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n354_), .A2(G197gat), .ZN(new_n355_));
  INV_X1    g154(.A(new_n336_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n332_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n352_), .B1(new_n353_), .B2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n347_), .A2(new_n348_), .A3(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n343_), .A2(new_n346_), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n346_), .B1(new_n343_), .B2(new_n359_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT89), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n346_), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n340_), .A2(new_n342_), .A3(G106gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n348_), .B1(new_n347_), .B2(new_n358_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n343_), .A2(new_n359_), .A3(new_n346_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(KEYINPUT86), .A3(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n299_), .A2(new_n341_), .A3(new_n300_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT28), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n299_), .A2(new_n371_), .A3(new_n300_), .A4(new_n341_), .ZN(new_n372_));
  XOR2_X1   g171(.A(G22gat), .B(G50gat), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT89), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n370_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n362_), .A2(new_n368_), .A3(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n377_), .A2(new_n366_), .A3(KEYINPUT86), .A4(new_n367_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  XOR2_X1   g180(.A(G8gat), .B(G36gat), .Z(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT18), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT90), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n225_), .A2(G183gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n223_), .A2(KEYINPUT25), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n387_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n224_), .A2(new_n226_), .A3(KEYINPUT90), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(new_n247_), .A3(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n245_), .A2(new_n232_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT91), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n243_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n392_), .A2(new_n393_), .A3(KEYINPUT91), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n331_), .A2(new_n337_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n396_), .A2(new_n397_), .B1(new_n398_), .B2(new_n352_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT20), .B1(new_n358_), .B2(new_n237_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G226gat), .A2(G233gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT19), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n399_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n402_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n340_), .A2(new_n218_), .A3(new_n394_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT20), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n406_), .B1(new_n358_), .B2(new_n237_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n386_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n402_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n340_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n411_), .A2(new_n407_), .A3(new_n404_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n410_), .A2(new_n412_), .A3(new_n385_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n409_), .A2(KEYINPUT27), .A3(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(KEYINPUT93), .B(KEYINPUT27), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n396_), .A2(new_n397_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n358_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n406_), .B1(new_n340_), .B2(new_n249_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n404_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n411_), .A2(new_n407_), .A3(new_n404_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n386_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n415_), .B1(new_n421_), .B2(new_n413_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n414_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n318_), .A2(new_n381_), .A3(new_n423_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n379_), .A2(new_n380_), .A3(new_n316_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n385_), .A2(KEYINPUT32), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n410_), .A2(new_n412_), .A3(new_n426_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n428_), .B(new_n429_), .C1(new_n314_), .C2(new_n315_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n303_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n313_), .B1(new_n302_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n292_), .A2(new_n301_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT92), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n431_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n434_), .A2(KEYINPUT92), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n433_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n421_), .A2(new_n438_), .A3(new_n413_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n307_), .A2(new_n308_), .A3(new_n313_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT33), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n307_), .A2(KEYINPUT33), .A3(new_n308_), .A4(new_n313_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n430_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n445_));
  AOI22_X1  g244(.A1(new_n425_), .A2(new_n423_), .B1(new_n445_), .B2(new_n381_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n268_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n424_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G190gat), .B(G218gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G134gat), .B(G162gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT36), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G99gat), .A2(G106gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT6), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT6), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(G99gat), .A3(G106gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n457_), .B1(new_n460_), .B2(G106gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(G85gat), .B(G92gat), .C1(KEYINPUT64), .C2(KEYINPUT9), .ZN(new_n463_));
  OAI211_X1 g262(.A(KEYINPUT64), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(KEYINPUT64), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n462_), .A2(KEYINPUT65), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT65), .ZN(new_n469_));
  INV_X1    g268(.A(new_n467_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n469_), .B1(new_n470_), .B2(new_n461_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT66), .ZN(new_n472_));
  INV_X1    g271(.A(G99gat), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(new_n348_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT7), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT7), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n472_), .A2(new_n476_), .A3(new_n473_), .A4(new_n348_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n457_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT8), .ZN(new_n479_));
  XOR2_X1   g278(.A(G85gat), .B(G92gat), .Z(new_n480_));
  AND3_X1   g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n479_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n482_));
  OAI211_X1 g281(.A(new_n468_), .B(new_n471_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n483_));
  XOR2_X1   g282(.A(G29gat), .B(G36gat), .Z(new_n484_));
  XOR2_X1   g283(.A(G43gat), .B(G50gat), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G232gat), .A2(G233gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT34), .ZN(new_n489_));
  OAI22_X1  g288(.A1(new_n483_), .A2(new_n487_), .B1(KEYINPUT35), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n468_), .A2(new_n471_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n481_), .A2(new_n482_), .A3(KEYINPUT68), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT68), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n478_), .A2(new_n480_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT8), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n495_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n493_), .B1(new_n494_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT15), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n486_), .B(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT71), .B1(new_n500_), .B2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT68), .B1(new_n481_), .B2(new_n482_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n497_), .A2(new_n495_), .A3(new_n498_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n492_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT71), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n507_), .A2(new_n508_), .A3(new_n502_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n491_), .B1(new_n504_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n489_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT35), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n500_), .A2(KEYINPUT71), .A3(new_n503_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n508_), .B1(new_n507_), .B2(new_n502_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n513_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n491_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n452_), .B1(new_n514_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT72), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n514_), .A2(new_n521_), .A3(new_n519_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n451_), .A2(KEYINPUT36), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n514_), .A2(new_n521_), .A3(new_n519_), .A4(new_n523_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n520_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  AND2_X1   g326(.A1(new_n448_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT77), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT73), .B(G8gat), .ZN(new_n530_));
  INV_X1    g329(.A(G1gat), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT14), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G15gat), .B(G22gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G1gat), .B(G8gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n532_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n486_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n539_), .A2(new_n486_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n529_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  AND2_X1   g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n537_), .A2(new_n538_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n487_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n546_), .A2(KEYINPUT77), .A3(new_n540_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n543_), .A2(new_n544_), .A3(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n540_), .B1(new_n502_), .B2(new_n539_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n548_), .B1(new_n544_), .B2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G169gat), .B(G197gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n550_), .A2(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n548_), .B(new_n553_), .C1(new_n544_), .C2(new_n549_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT5), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G176gat), .B(G204gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G57gat), .B(G64gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT11), .ZN(new_n564_));
  XOR2_X1   g363(.A(G71gat), .B(G78gat), .Z(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n563_), .A2(KEYINPUT11), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n564_), .A2(new_n565_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n483_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(KEYINPUT12), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n571_), .B1(new_n500_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G230gat), .A2(G233gat), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n483_), .A2(new_n570_), .ZN(new_n576_));
  XOR2_X1   g375(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n577_));
  AND3_X1   g376(.A1(new_n576_), .A2(KEYINPUT70), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT70), .B1(new_n576_), .B2(new_n577_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n574_), .B(new_n575_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n575_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n571_), .A2(KEYINPUT67), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(new_n576_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n571_), .A2(KEYINPUT67), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n581_), .B1(new_n583_), .B2(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n562_), .B1(new_n580_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n580_), .A2(new_n585_), .A3(new_n562_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n587_), .A2(KEYINPUT13), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT13), .ZN(new_n590_));
  INV_X1    g389(.A(new_n588_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n590_), .B1(new_n591_), .B2(new_n586_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(G231gat), .ZN(new_n595_));
  INV_X1    g394(.A(G233gat), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n597_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n569_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n597_), .ZN(new_n600_));
  OAI211_X1 g399(.A(new_n599_), .B(new_n600_), .C1(new_n567_), .C2(new_n566_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(new_n539_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n545_), .A2(new_n598_), .A3(new_n601_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(G183gat), .B(G211gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT17), .B1(new_n605_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT75), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n603_), .A2(new_n612_), .A3(new_n604_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n610_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(KEYINPUT17), .A3(new_n610_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n528_), .A2(new_n557_), .A3(new_n594_), .A4(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(G1gat), .B1(new_n618_), .B2(new_n316_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n520_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n518_), .B1(new_n517_), .B2(new_n491_), .ZN(new_n621_));
  AOI211_X1 g420(.A(new_n513_), .B(new_n490_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n523_), .B1(new_n623_), .B2(new_n521_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n526_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n620_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT37), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT37), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n527_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n615_), .A2(KEYINPUT76), .A3(new_n616_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT76), .B1(new_n615_), .B2(new_n616_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n630_), .A2(new_n593_), .A3(new_n633_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n448_), .A2(new_n557_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NOR3_X1   g435(.A1(new_n636_), .A2(G1gat), .A3(new_n316_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n619_), .B1(new_n637_), .B2(KEYINPUT38), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n638_), .B1(KEYINPUT38), .B2(new_n637_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT94), .ZN(G1324gat));
  OAI21_X1  g439(.A(G8gat), .B1(new_n618_), .B2(new_n423_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT39), .ZN(new_n642_));
  INV_X1    g441(.A(new_n423_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n530_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n642_), .B1(new_n636_), .B2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(KEYINPUT95), .B(KEYINPUT40), .Z(new_n646_));
  XNOR2_X1  g445(.A(new_n645_), .B(new_n646_), .ZN(G1325gat));
  OAI21_X1  g446(.A(G15gat), .B1(new_n618_), .B2(new_n268_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT41), .Z(new_n649_));
  OR2_X1    g448(.A1(new_n268_), .A2(G15gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n649_), .B1(new_n636_), .B2(new_n650_), .ZN(G1326gat));
  OAI21_X1  g450(.A(G22gat), .B1(new_n618_), .B2(new_n381_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT42), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n381_), .A2(G22gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT96), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n653_), .B1(new_n636_), .B2(new_n655_), .ZN(G1327gat));
  NAND4_X1  g455(.A1(new_n635_), .A2(new_n594_), .A3(new_n626_), .A4(new_n633_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT101), .ZN(new_n658_));
  INV_X1    g457(.A(G29gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n658_), .A2(new_n659_), .A3(new_n317_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT99), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n589_), .A2(new_n592_), .A3(new_n557_), .A4(new_n633_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT97), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n525_), .A2(new_n526_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n628_), .B1(new_n664_), .B2(new_n620_), .ZN(new_n665_));
  AOI211_X1 g464(.A(KEYINPUT37), .B(new_n520_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n448_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT43), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT43), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n448_), .B(new_n669_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n663_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n316_), .B1(new_n671_), .B2(KEYINPUT44), .ZN(new_n672_));
  INV_X1    g471(.A(new_n663_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n669_), .B1(new_n630_), .B2(new_n448_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n670_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT98), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT98), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n671_), .A2(new_n679_), .A3(KEYINPUT44), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n661_), .B(new_n672_), .C1(new_n678_), .C2(new_n680_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(G29gat), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT100), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n676_), .A2(KEYINPUT98), .A3(new_n677_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n679_), .B1(new_n671_), .B2(KEYINPUT44), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n661_), .B1(new_n686_), .B2(new_n672_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n682_), .A2(new_n683_), .A3(new_n687_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT44), .B(new_n673_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n317_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n685_), .B2(new_n684_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n659_), .B1(new_n691_), .B2(new_n661_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n686_), .A2(new_n672_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT99), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT100), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n660_), .B1(new_n688_), .B2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT102), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n698_), .B(new_n660_), .C1(new_n688_), .C2(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1328gat));
  INV_X1    g499(.A(G36gat), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n643_), .A2(KEYINPUT103), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n643_), .A2(KEYINPUT103), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n658_), .A2(new_n701_), .A3(new_n704_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT45), .Z(new_n706_));
  AND2_X1   g505(.A1(new_n686_), .A2(new_n689_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n701_), .B1(new_n707_), .B2(new_n643_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  OR2_X1    g508(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n709_), .B(new_n710_), .ZN(G1329gat));
  AOI21_X1  g510(.A(G43gat), .B1(new_n658_), .B2(new_n447_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n447_), .A2(G43gat), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n707_), .B2(new_n714_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g515(.A(new_n381_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G50gat), .B1(new_n658_), .B2(new_n717_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n717_), .A2(G50gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n707_), .B2(new_n719_), .ZN(G1331gat));
  INV_X1    g519(.A(new_n557_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n633_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n528_), .A2(new_n721_), .A3(new_n593_), .A4(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(G57gat), .B1(new_n723_), .B2(new_n316_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n630_), .A2(new_n594_), .A3(new_n633_), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n725_), .A2(KEYINPUT105), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n448_), .A2(new_n721_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n725_), .A2(KEYINPUT105), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n726_), .A2(new_n727_), .A3(new_n728_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n316_), .A2(G57gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n724_), .B1(new_n729_), .B2(new_n730_), .ZN(G1332gat));
  INV_X1    g530(.A(new_n704_), .ZN(new_n732_));
  OAI21_X1  g531(.A(G64gat), .B1(new_n723_), .B2(new_n732_), .ZN(new_n733_));
  XOR2_X1   g532(.A(KEYINPUT106), .B(KEYINPUT48), .Z(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n732_), .A2(G64gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n729_), .B2(new_n736_), .ZN(G1333gat));
  OAI21_X1  g536(.A(G71gat), .B1(new_n723_), .B2(new_n268_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT49), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n268_), .A2(G71gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n729_), .B2(new_n740_), .ZN(G1334gat));
  OAI21_X1  g540(.A(G78gat), .B1(new_n723_), .B2(new_n381_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT50), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n717_), .A2(new_n345_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n729_), .B2(new_n744_), .ZN(G1335gat));
  NAND2_X1  g544(.A1(new_n668_), .A2(new_n670_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n594_), .A2(new_n557_), .A3(new_n722_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n748_), .A2(KEYINPUT107), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(KEYINPUT107), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n310_), .B1(new_n751_), .B2(new_n317_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n594_), .A2(new_n527_), .A3(new_n722_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n727_), .A2(new_n753_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n754_), .A2(G85gat), .A3(new_n316_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n752_), .A2(new_n755_), .ZN(G1336gat));
  INV_X1    g555(.A(new_n754_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G92gat), .B1(new_n757_), .B2(new_n643_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n704_), .A2(G92gat), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT108), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n758_), .B1(new_n751_), .B2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT109), .ZN(G1337gat));
  NOR3_X1   g561(.A1(new_n754_), .A2(new_n268_), .A3(new_n460_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n751_), .A2(new_n447_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(G99gat), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT110), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n765_), .A2(KEYINPUT110), .A3(new_n766_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n765_), .A2(KEYINPUT111), .A3(new_n766_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT111), .B1(new_n765_), .B2(new_n766_), .ZN(new_n772_));
  OAI22_X1  g571(.A1(new_n769_), .A2(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(G1338gat));
  NAND3_X1  g572(.A1(new_n746_), .A2(new_n717_), .A3(new_n747_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT112), .B1(new_n774_), .B2(G106gat), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(KEYINPUT112), .A3(G106gat), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n754_), .A2(G106gat), .A3(new_n381_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g582(.A1(new_n447_), .A2(new_n381_), .A3(new_n423_), .A4(new_n317_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT117), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n617_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n543_), .A2(new_n547_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n549_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n544_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n549_), .A2(new_n789_), .ZN(new_n792_));
  OAI221_X1 g591(.A(new_n554_), .B1(new_n788_), .B2(new_n544_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n793_), .A2(new_n556_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n794_), .A2(new_n588_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796_));
  OR3_X1    g595(.A1(new_n580_), .A2(KEYINPUT115), .A3(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(KEYINPUT115), .B1(new_n580_), .B2(new_n796_), .ZN(new_n798_));
  XOR2_X1   g597(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n799_));
  OAI21_X1  g598(.A(new_n574_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n581_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n580_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n797_), .B(new_n798_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n803_), .A2(KEYINPUT56), .A3(new_n561_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT56), .B1(new_n803_), .B2(new_n561_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n795_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n795_), .B(KEYINPUT58), .C1(new_n805_), .C2(new_n806_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n630_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n557_), .A2(new_n588_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT113), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n587_), .A2(new_n588_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n794_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n626_), .B1(new_n815_), .B2(new_n817_), .ZN(new_n818_));
  OAI22_X1  g617(.A1(new_n810_), .A2(new_n812_), .B1(new_n818_), .B2(KEYINPUT57), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n813_), .B(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n806_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n804_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n817_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n527_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n787_), .B1(new_n819_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n634_), .A2(new_n721_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT54), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n634_), .A2(new_n831_), .A3(new_n721_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n786_), .B1(new_n828_), .B2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(G113gat), .B1(new_n834_), .B2(new_n557_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n811_), .A2(new_n630_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n809_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n825_), .A2(new_n826_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n818_), .A2(KEYINPUT57), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n840_), .A2(new_n787_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT59), .B1(new_n841_), .B2(new_n786_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n786_), .A2(KEYINPUT59), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n809_), .A2(new_n836_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n722_), .B1(new_n844_), .B2(new_n839_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n833_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n843_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n842_), .A2(new_n847_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT118), .B(G113gat), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n557_), .A2(new_n849_), .ZN(new_n850_));
  XNOR2_X1  g649(.A(new_n850_), .B(KEYINPUT119), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n835_), .B1(new_n848_), .B2(new_n851_), .ZN(G1340gat));
  INV_X1    g651(.A(G120gat), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n842_), .A2(new_n593_), .A3(new_n847_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n855_), .B2(new_n854_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n853_), .B1(new_n594_), .B2(KEYINPUT60), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n834_), .B(new_n858_), .C1(KEYINPUT60), .C2(new_n853_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(G1341gat));
  NAND2_X1  g659(.A1(new_n848_), .A2(new_n617_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(G127gat), .ZN(new_n862_));
  INV_X1    g661(.A(new_n834_), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n633_), .A2(G127gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n862_), .B1(new_n863_), .B2(new_n864_), .ZN(G1342gat));
  NAND4_X1  g664(.A1(new_n842_), .A2(new_n847_), .A3(G134gat), .A4(new_n630_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867_));
  AOI211_X1 g666(.A(new_n867_), .B(G134gat), .C1(new_n834_), .C2(new_n626_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n828_), .A2(new_n833_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n869_), .A2(new_n626_), .A3(new_n785_), .ZN(new_n870_));
  INV_X1    g669(.A(G134gat), .ZN(new_n871_));
  AOI21_X1  g670(.A(KEYINPUT121), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n866_), .B1(new_n868_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  OAI211_X1 g674(.A(KEYINPUT122), .B(new_n866_), .C1(new_n868_), .C2(new_n872_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1343gat));
  NOR2_X1   g676(.A1(new_n841_), .A2(new_n447_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n704_), .A2(new_n381_), .A3(new_n316_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n557_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n593_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g684(.A1(new_n880_), .A2(new_n633_), .ZN(new_n886_));
  XOR2_X1   g685(.A(KEYINPUT61), .B(G155gat), .Z(new_n887_));
  XNOR2_X1  g686(.A(new_n886_), .B(new_n887_), .ZN(G1346gat));
  AOI21_X1  g687(.A(G162gat), .B1(new_n881_), .B2(new_n626_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n630_), .A2(G162gat), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(KEYINPUT123), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n889_), .B1(new_n881_), .B2(new_n891_), .ZN(G1347gat));
  OR2_X1    g691(.A1(new_n845_), .A2(new_n846_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n704_), .A2(new_n381_), .A3(new_n318_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n893_), .A2(new_n557_), .A3(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n896_), .A2(new_n897_), .A3(G169gat), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n897_), .B1(new_n896_), .B2(G169gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n893_), .A2(new_n895_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(KEYINPUT22), .B(G169gat), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n557_), .A2(new_n901_), .ZN(new_n902_));
  XOR2_X1   g701(.A(new_n902_), .B(KEYINPUT124), .Z(new_n903_));
  OAI22_X1  g702(.A1(new_n898_), .A2(new_n899_), .B1(new_n900_), .B2(new_n903_), .ZN(G1348gat));
  INV_X1    g703(.A(new_n900_), .ZN(new_n905_));
  AOI21_X1  g704(.A(G176gat), .B1(new_n905_), .B2(new_n593_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n841_), .A2(new_n894_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n907_), .A2(G176gat), .A3(new_n593_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT125), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n908_), .A2(new_n909_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n906_), .A2(new_n910_), .A3(new_n911_), .ZN(G1349gat));
  AOI21_X1  g711(.A(G183gat), .B1(new_n907_), .B2(new_n722_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n787_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n913_), .B1(new_n905_), .B2(new_n914_), .ZN(G1350gat));
  INV_X1    g714(.A(new_n630_), .ZN(new_n916_));
  OAI21_X1  g715(.A(G190gat), .B1(new_n900_), .B2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n626_), .A2(new_n247_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n900_), .B2(new_n918_), .ZN(G1351gat));
  AND2_X1   g718(.A1(new_n704_), .A2(new_n425_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n878_), .A2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n721_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(new_n334_), .ZN(G1352gat));
  INV_X1    g722(.A(KEYINPUT126), .ZN(new_n924_));
  NOR4_X1   g723(.A1(new_n921_), .A2(new_n924_), .A3(new_n354_), .A4(new_n594_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n921_), .A2(new_n594_), .ZN(new_n926_));
  AOI21_X1  g725(.A(KEYINPUT126), .B1(new_n926_), .B2(new_n325_), .ZN(new_n927_));
  OAI21_X1  g726(.A(G204gat), .B1(new_n921_), .B2(new_n594_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n925_), .B1(new_n927_), .B2(new_n928_), .ZN(G1353gat));
  XOR2_X1   g728(.A(KEYINPUT63), .B(G211gat), .Z(new_n930_));
  NAND4_X1  g729(.A1(new_n878_), .A2(new_n617_), .A3(new_n920_), .A4(new_n930_), .ZN(new_n931_));
  OR2_X1    g730(.A1(new_n931_), .A2(KEYINPUT127), .ZN(new_n932_));
  NOR2_X1   g731(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n933_), .B1(new_n921_), .B2(new_n787_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n931_), .A2(KEYINPUT127), .ZN(new_n935_));
  AND3_X1   g734(.A1(new_n932_), .A2(new_n934_), .A3(new_n935_), .ZN(G1354gat));
  OAI21_X1  g735(.A(G218gat), .B1(new_n921_), .B2(new_n916_), .ZN(new_n937_));
  OR2_X1    g736(.A1(new_n527_), .A2(G218gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n921_), .B2(new_n938_), .ZN(G1355gat));
endmodule


