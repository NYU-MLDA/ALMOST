//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT86), .ZN(new_n207_));
  INV_X1    g006(.A(G204gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n207_), .B1(new_n208_), .B2(G197gat), .ZN(new_n209_));
  INV_X1    g008(.A(G197gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(KEYINPUT86), .A3(G204gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT21), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n208_), .A2(G197gat), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n209_), .A2(new_n211_), .A3(new_n212_), .A4(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n213_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n208_), .A2(G197gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT21), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(G211gat), .B(G218gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT87), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G211gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(G218gat), .ZN(new_n222_));
  INV_X1    g021(.A(G218gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n223_), .A2(G211gat), .ZN(new_n224_));
  NOR3_X1   g023(.A1(new_n222_), .A2(new_n224_), .A3(KEYINPUT87), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n214_), .B(new_n217_), .C1(new_n220_), .C2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n218_), .A2(new_n219_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT87), .B1(new_n222_), .B2(new_n224_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n209_), .A2(new_n211_), .A3(new_n213_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(KEYINPUT21), .A4(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n226_), .A2(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT25), .B(G183gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT26), .B(G190gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G183gat), .ZN(new_n235_));
  INV_X1    g034(.A(G190gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT23), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n238_), .A2(G183gat), .A3(G190gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G169gat), .A2(G176gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G169gat), .A2(G176gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(KEYINPUT24), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT24), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n241_), .A2(new_n245_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n234_), .A2(new_n240_), .A3(new_n244_), .A4(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT79), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n237_), .A2(new_n248_), .A3(new_n239_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n238_), .A2(KEYINPUT79), .A3(G183gat), .A4(G190gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n235_), .A2(new_n236_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n249_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT78), .B(G176gat), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT77), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT22), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(new_n255_), .A3(G169gat), .ZN(new_n256_));
  INV_X1    g055(.A(G169gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT22), .B1(new_n257_), .B2(KEYINPUT77), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n253_), .A2(new_n256_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(new_n243_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n247_), .B1(new_n252_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT80), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT80), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n263_), .B(new_n247_), .C1(new_n252_), .C2(new_n260_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n231_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n232_), .A2(new_n233_), .B1(new_n245_), .B2(new_n241_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n266_), .A2(new_n244_), .A3(new_n250_), .A4(new_n249_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT22), .B(G169gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n253_), .A2(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(KEYINPUT93), .A3(new_n243_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n240_), .A2(new_n251_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n253_), .A2(new_n268_), .B1(G169gat), .B2(G176gat), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(KEYINPUT93), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n267_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n226_), .A2(new_n230_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT20), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G226gat), .A2(G233gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n265_), .A2(new_n277_), .A3(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n262_), .A2(new_n231_), .A3(new_n264_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT20), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n280_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n206_), .B1(new_n282_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n285_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n281_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n264_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n249_), .A2(new_n250_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n251_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n243_), .B(new_n259_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n263_), .B1(new_n293_), .B2(new_n247_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n276_), .B1(new_n290_), .B2(new_n294_), .ZN(new_n295_));
  AOI22_X1  g094(.A1(new_n273_), .A2(KEYINPUT93), .B1(new_n240_), .B2(new_n251_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n273_), .A2(KEYINPUT93), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n266_), .A2(new_n244_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n291_), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n296_), .A2(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n284_), .B1(new_n300_), .B2(new_n231_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n295_), .A2(new_n301_), .A3(new_n280_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n289_), .A2(new_n205_), .A3(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n287_), .A2(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n304_), .A2(KEYINPUT27), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n283_), .A2(new_n285_), .A3(new_n280_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n281_), .B1(new_n265_), .B2(new_n277_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(KEYINPUT96), .B2(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n280_), .B1(new_n295_), .B2(new_n301_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT96), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n205_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n303_), .A2(KEYINPUT27), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT97), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  OAI22_X1  g113(.A1(new_n309_), .A2(new_n310_), .B1(new_n281_), .B2(new_n288_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n307_), .A2(KEYINPUT96), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n206_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n303_), .A2(KEYINPUT27), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT97), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n305_), .B1(new_n314_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT82), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT82), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n325_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT2), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(G141gat), .ZN(new_n331_));
  INV_X1    g130(.A(G148gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(KEYINPUT3), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT3), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(G141gat), .B2(G148gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n327_), .A2(new_n330_), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT83), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G155gat), .B(G162gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT83), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n327_), .A2(new_n336_), .A3(new_n341_), .A4(new_n330_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n338_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n339_), .A2(KEYINPUT1), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n331_), .A2(new_n332_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(new_n328_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n344_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n343_), .A2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G127gat), .B(G134gat), .Z(new_n351_));
  XOR2_X1   g150(.A(G113gat), .B(G120gat), .Z(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  NAND2_X1  g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n339_), .B1(new_n337_), .B2(KEYINPUT83), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n348_), .B1(new_n355_), .B2(new_n342_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n353_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n354_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n354_), .A2(KEYINPUT4), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT94), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n354_), .A2(KEYINPUT4), .A3(new_n358_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n359_), .A2(KEYINPUT94), .A3(KEYINPUT4), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n362_), .B1(new_n368_), .B2(new_n361_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G1gat), .B(G29gat), .Z(new_n370_));
  XNOR2_X1  g169(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G57gat), .B(G85gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n372_), .B(new_n373_), .Z(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n369_), .A2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n360_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n377_), .A2(new_n374_), .A3(new_n362_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G228gat), .A2(G233gat), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT29), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n276_), .B1(new_n356_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT85), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n381_), .B(new_n382_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n231_), .B1(new_n350_), .B2(KEYINPUT29), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT88), .B1(new_n387_), .B2(KEYINPUT85), .ZN(new_n388_));
  INV_X1    g187(.A(new_n382_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(new_n384_), .B2(new_n381_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n386_), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G78gat), .B(G106gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT89), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n391_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT91), .ZN(new_n395_));
  INV_X1    g194(.A(new_n392_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT91), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n391_), .A2(new_n398_), .A3(new_n393_), .ZN(new_n399_));
  XOR2_X1   g198(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n350_), .B2(KEYINPUT29), .ZN(new_n401_));
  XOR2_X1   g200(.A(G22gat), .B(G50gat), .Z(new_n402_));
  INV_X1    g201(.A(new_n400_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n356_), .A2(new_n383_), .A3(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n401_), .A2(new_n402_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n402_), .B1(new_n401_), .B2(new_n404_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n395_), .A2(new_n397_), .A3(new_n399_), .A4(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT90), .ZN(new_n409_));
  INV_X1    g208(.A(new_n393_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n386_), .B(new_n410_), .C1(new_n388_), .C2(new_n390_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n394_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n407_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n409_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  AOI211_X1 g213(.A(KEYINPUT90), .B(new_n407_), .C1(new_n394_), .C2(new_n411_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n408_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n290_), .A2(new_n294_), .ZN(new_n417_));
  XOR2_X1   g216(.A(G71gat), .B(G99gat), .Z(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT81), .B(G43gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n417_), .B(new_n420_), .ZN(new_n421_));
  AND2_X1   g220(.A1(new_n421_), .A2(new_n357_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n357_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G227gat), .A2(G233gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n424_), .B(G15gat), .Z(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT30), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT31), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  OR3_X1    g227(.A1(new_n422_), .A2(new_n423_), .A3(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n428_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NOR4_X1   g231(.A1(new_n322_), .A2(new_n380_), .A3(new_n416_), .A4(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n416_), .A2(new_n321_), .A3(new_n379_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT98), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT98), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n416_), .A2(new_n321_), .A3(new_n436_), .A4(new_n379_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT33), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n369_), .B2(new_n375_), .ZN(new_n439_));
  OAI211_X1 g238(.A(KEYINPUT33), .B(new_n374_), .C1(new_n377_), .C2(new_n362_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n374_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n441_), .B1(new_n368_), .B2(new_n361_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n439_), .A2(new_n304_), .A3(new_n440_), .A4(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n282_), .A2(new_n286_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n308_), .A2(new_n311_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n446_), .B1(new_n447_), .B2(new_n445_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n416_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n435_), .A2(new_n437_), .A3(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n433_), .B1(new_n453_), .B2(new_n432_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT74), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G29gat), .B(G36gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT69), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G43gat), .B(G50gat), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n456_), .A2(KEYINPUT69), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n456_), .A2(KEYINPUT69), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n462_), .A3(new_n458_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G15gat), .B(G22gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(KEYINPUT72), .B(G8gat), .ZN(new_n466_));
  INV_X1    g265(.A(G1gat), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT14), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n465_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G1gat), .B(G8gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n465_), .B(new_n471_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n455_), .B1(new_n464_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n460_), .A2(new_n463_), .ZN(new_n477_));
  NAND4_X1  g276(.A1(new_n477_), .A2(KEYINPUT74), .A3(new_n474_), .A4(new_n473_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n464_), .A2(KEYINPUT73), .A3(new_n475_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(KEYINPUT73), .B1(new_n464_), .B2(new_n475_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n479_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT75), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G229gat), .A2(G233gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n482_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n480_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(KEYINPUT75), .A3(new_n479_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n485_), .A2(new_n487_), .A3(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n481_), .A2(new_n482_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n477_), .B(KEYINPUT15), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n493_), .A2(new_n475_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n486_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(G113gat), .B(G141gat), .Z(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT76), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G169gat), .B(G197gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n498_), .B(new_n499_), .Z(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n500_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n491_), .A2(new_n495_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n501_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n454_), .A2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(KEYINPUT10), .B(G99gat), .Z(new_n507_));
  INV_X1    g306(.A(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G85gat), .B(G92gat), .Z(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT9), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT6), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(G99gat), .A3(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(G85gat), .ZN(new_n517_));
  INV_X1    g316(.A(G92gat), .ZN(new_n518_));
  OR3_X1    g317(.A1(new_n517_), .A2(new_n518_), .A3(KEYINPUT9), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n509_), .A2(new_n511_), .A3(new_n516_), .A4(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT8), .ZN(new_n521_));
  NOR2_X1   g320(.A1(G99gat), .A2(G106gat), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT7), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT64), .B1(new_n513_), .B2(new_n515_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n513_), .A2(new_n515_), .A3(KEYINPUT64), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n521_), .B1(new_n529_), .B2(new_n510_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n516_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n521_), .B(new_n510_), .C1(new_n524_), .C2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n520_), .B1(new_n530_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n493_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n520_), .ZN(new_n536_));
  NOR3_X1   g335(.A1(new_n524_), .A2(new_n527_), .A3(new_n525_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n510_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT8), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n536_), .B1(new_n539_), .B2(new_n532_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(new_n477_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n535_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G232gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n542_), .A2(KEYINPUT70), .A3(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT35), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n535_), .A2(new_n548_), .A3(new_n541_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n546_), .B1(new_n542_), .B2(KEYINPUT70), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n547_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G190gat), .B(G218gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G134gat), .B(G162gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n554_), .B(KEYINPUT36), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n551_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n542_), .A2(KEYINPUT70), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(new_n549_), .A3(new_n545_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n554_), .A2(KEYINPUT36), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n542_), .A2(KEYINPUT70), .A3(new_n546_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT37), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n557_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT71), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n555_), .B1(new_n551_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n559_), .A2(new_n561_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n567_), .A2(KEYINPUT71), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n562_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT37), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n564_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572_));
  XOR2_X1   g371(.A(G127gat), .B(G155gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT16), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n475_), .B(new_n577_), .Z(new_n578_));
  XNOR2_X1  g377(.A(G57gat), .B(G64gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT11), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT65), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n579_), .A2(KEYINPUT11), .ZN(new_n582_));
  XOR2_X1   g381(.A(G71gat), .B(G78gat), .Z(new_n583_));
  INV_X1    g382(.A(KEYINPUT65), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n579_), .A2(new_n584_), .A3(KEYINPUT11), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n581_), .A2(new_n582_), .A3(new_n583_), .A4(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n583_), .B1(KEYINPUT11), .B2(new_n579_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n579_), .A2(new_n584_), .A3(KEYINPUT11), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n584_), .B1(new_n579_), .B2(KEYINPUT11), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n587_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n586_), .A2(new_n590_), .ZN(new_n591_));
  AOI211_X1 g390(.A(new_n572_), .B(new_n576_), .C1(new_n578_), .C2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n591_), .B2(new_n578_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT66), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n586_), .A2(new_n590_), .A3(KEYINPUT66), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n578_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n578_), .A2(new_n597_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n576_), .B(KEYINPUT17), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n593_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n571_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n595_), .A2(new_n596_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(new_n540_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n586_), .A2(new_n590_), .A3(KEYINPUT12), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n534_), .A2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT68), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G230gat), .A2(G233gat), .ZN(new_n611_));
  XOR2_X1   g410(.A(KEYINPUT67), .B(KEYINPUT12), .Z(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n613_), .B1(new_n605_), .B2(new_n540_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n609_), .A2(new_n610_), .A3(new_n611_), .A4(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n614_), .A2(new_n611_), .A3(new_n606_), .A4(new_n608_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT68), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n597_), .A2(new_n534_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(new_n606_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n619_), .A2(G230gat), .A3(G233gat), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n615_), .A2(new_n617_), .A3(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G120gat), .B(G148gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT5), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G176gat), .B(G204gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n623_), .B(new_n624_), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n621_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n625_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n615_), .A2(new_n617_), .A3(new_n620_), .A4(new_n627_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n626_), .A2(KEYINPUT13), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT13), .B1(new_n626_), .B2(new_n628_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n604_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n506_), .A2(new_n633_), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n634_), .A2(G1gat), .A3(new_n379_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n635_), .A2(KEYINPUT38), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(KEYINPUT38), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n556_), .B1(new_n567_), .B2(KEYINPUT71), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n551_), .A2(new_n565_), .ZN(new_n639_));
  AOI22_X1  g438(.A1(new_n638_), .A2(new_n639_), .B1(new_n560_), .B2(new_n551_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n454_), .A2(new_n602_), .A3(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n632_), .A2(new_n505_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n379_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n636_), .A2(new_n637_), .A3(new_n644_), .ZN(G1324gat));
  OAI21_X1  g444(.A(G8gat), .B1(new_n643_), .B2(new_n321_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT39), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n322_), .A2(new_n466_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n647_), .B1(new_n634_), .B2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n649_), .B(new_n651_), .ZN(G1325gat));
  OAI21_X1  g451(.A(G15gat), .B1(new_n643_), .B2(new_n432_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT41), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n634_), .A2(G15gat), .A3(new_n432_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1326gat));
  OAI21_X1  g455(.A(G22gat), .B1(new_n643_), .B2(new_n451_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT42), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n451_), .A2(G22gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n658_), .B1(new_n634_), .B2(new_n659_), .ZN(G1327gat));
  NAND2_X1  g459(.A1(new_n640_), .A2(new_n602_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n632_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n506_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT103), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n506_), .A2(new_n665_), .A3(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  OR3_X1    g466(.A1(new_n667_), .A2(G29gat), .A3(new_n379_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n642_), .A2(new_n602_), .ZN(new_n670_));
  OAI21_X1  g469(.A(KEYINPUT43), .B1(new_n454_), .B2(new_n571_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT43), .ZN(new_n672_));
  OAI22_X1  g471(.A1(new_n640_), .A2(KEYINPUT37), .B1(new_n557_), .B2(new_n563_), .ZN(new_n673_));
  AOI22_X1  g472(.A1(new_n434_), .A2(KEYINPUT98), .B1(new_n450_), .B2(new_n451_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n431_), .B1(new_n674_), .B2(new_n437_), .ZN(new_n675_));
  OAI211_X1 g474(.A(new_n672_), .B(new_n673_), .C1(new_n675_), .C2(new_n433_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n670_), .B1(new_n671_), .B2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n669_), .B1(new_n677_), .B2(KEYINPUT44), .ZN(new_n678_));
  INV_X1    g477(.A(new_n670_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n453_), .A2(new_n432_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n433_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n672_), .B1(new_n682_), .B2(new_n673_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n454_), .A2(KEYINPUT43), .A3(new_n571_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n679_), .B1(new_n683_), .B2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n685_), .A2(KEYINPUT100), .A3(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(KEYINPUT44), .B(new_n679_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT101), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT101), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n677_), .A2(new_n690_), .A3(KEYINPUT44), .ZN(new_n691_));
  AOI22_X1  g490(.A1(new_n678_), .A2(new_n687_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(KEYINPUT102), .A3(new_n380_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(G29gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT102), .B1(new_n692_), .B2(new_n380_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n668_), .B1(new_n694_), .B2(new_n695_), .ZN(G1328gat));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n692_), .B2(new_n322_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n664_), .A2(new_n698_), .A3(new_n322_), .A4(new_n666_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT45), .Z(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n699_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n687_), .A2(new_n678_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n689_), .A2(new_n691_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G36gat), .B1(new_n705_), .B2(new_n321_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n700_), .B(KEYINPUT45), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(KEYINPUT46), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n702_), .A2(new_n708_), .ZN(G1329gat));
  INV_X1    g508(.A(G43gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n710_), .B1(new_n667_), .B2(new_n432_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n431_), .A2(G43gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n711_), .B1(new_n705_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT47), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n711_), .B(new_n715_), .C1(new_n705_), .C2(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1330gat));
  INV_X1    g516(.A(new_n667_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G50gat), .B1(new_n718_), .B2(new_n416_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n416_), .A2(G50gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n692_), .B2(new_n720_), .ZN(G1331gat));
  INV_X1    g520(.A(G57gat), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n454_), .A2(new_n504_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n723_), .A2(new_n632_), .A3(new_n603_), .A4(new_n571_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n722_), .B1(new_n724_), .B2(new_n379_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT104), .Z(new_n726_));
  NOR2_X1   g525(.A1(new_n631_), .A2(new_n504_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n641_), .A2(new_n727_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n728_), .A2(new_n722_), .A3(new_n379_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n726_), .A2(new_n729_), .ZN(G1332gat));
  OAI21_X1  g529(.A(G64gat), .B1(new_n728_), .B2(new_n321_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(KEYINPUT105), .B(KEYINPUT48), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n731_), .B(new_n732_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n321_), .A2(G64gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n724_), .B2(new_n734_), .ZN(G1333gat));
  OAI21_X1  g534(.A(G71gat), .B1(new_n728_), .B2(new_n432_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(KEYINPUT106), .B(KEYINPUT49), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n432_), .A2(G71gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n738_), .B1(new_n724_), .B2(new_n739_), .ZN(G1334gat));
  OAI21_X1  g539(.A(G78gat), .B1(new_n728_), .B2(new_n451_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n741_), .B(new_n742_), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n451_), .A2(G78gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n743_), .B1(new_n724_), .B2(new_n744_), .ZN(G1335gat));
  NAND2_X1  g544(.A1(new_n727_), .A2(new_n602_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n746_), .B1(new_n671_), .B2(new_n676_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(G85gat), .B1(new_n748_), .B2(new_n379_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n723_), .A2(new_n632_), .A3(new_n602_), .A4(new_n640_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n751_), .A2(new_n517_), .A3(new_n380_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n749_), .A2(new_n752_), .ZN(G1336gat));
  OAI21_X1  g552(.A(G92gat), .B1(new_n748_), .B2(new_n321_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n518_), .A3(new_n322_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1337gat));
  OAI21_X1  g555(.A(G99gat), .B1(new_n748_), .B2(new_n432_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n751_), .A2(new_n431_), .A3(new_n507_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g559(.A1(new_n751_), .A2(new_n508_), .A3(new_n416_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n508_), .B1(new_n747_), .B2(new_n416_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n762_), .A2(new_n763_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g566(.A1(new_n571_), .A2(new_n505_), .A3(new_n631_), .A4(new_n603_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT54), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n485_), .A2(new_n490_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n486_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n494_), .B1(new_n488_), .B2(new_n480_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n500_), .B1(new_n773_), .B2(new_n487_), .ZN(new_n774_));
  AOI22_X1  g573(.A1(new_n496_), .A2(new_n500_), .B1(new_n772_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n606_), .A2(new_n608_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n612_), .B1(new_n597_), .B2(new_n534_), .ZN(new_n777_));
  OAI211_X1 g576(.A(G230gat), .B(G233gat), .C1(new_n776_), .C2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT55), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(new_n616_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n615_), .A2(new_n617_), .A3(new_n779_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n627_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  OAI211_X1 g583(.A(new_n628_), .B(new_n775_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n615_), .A2(new_n617_), .A3(new_n779_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n625_), .B1(new_n786_), .B2(new_n780_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n787_), .A2(KEYINPUT56), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n770_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n775_), .A2(new_n628_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n783_), .A2(new_n784_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n787_), .A2(KEYINPUT56), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n790_), .A2(KEYINPUT58), .A3(new_n791_), .A4(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n673_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n626_), .A2(new_n628_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n775_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(KEYINPUT108), .A2(KEYINPUT56), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n625_), .B(new_n799_), .C1(new_n786_), .C2(new_n780_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n628_), .A2(new_n799_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n504_), .B(new_n800_), .C1(new_n783_), .C2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n775_), .A2(new_n795_), .A3(KEYINPUT109), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n798_), .A2(new_n802_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT110), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(KEYINPUT57), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(new_n569_), .A3(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n794_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n804_), .B2(new_n569_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n602_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n769_), .A2(new_n811_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n322_), .A2(new_n416_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(new_n380_), .A3(new_n431_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT111), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(KEYINPUT59), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n814_), .B1(new_n769_), .B2(new_n811_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  OAI21_X1  g619(.A(KEYINPUT111), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT112), .B(new_n602_), .C1(new_n809_), .C2(new_n810_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n804_), .A2(new_n569_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n806_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n826_), .A2(new_n794_), .A3(new_n808_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT112), .B1(new_n827_), .B2(new_n602_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n769_), .B1(new_n824_), .B2(new_n828_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(new_n820_), .A3(new_n815_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n504_), .A2(G113gat), .ZN(new_n831_));
  XOR2_X1   g630(.A(new_n831_), .B(KEYINPUT113), .Z(new_n832_));
  NAND3_X1  g631(.A1(new_n822_), .A2(new_n830_), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(G113gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n816_), .B2(new_n505_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT114), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1340gat));
  INV_X1    g637(.A(G120gat), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n631_), .B2(KEYINPUT60), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n819_), .B(new_n840_), .C1(KEYINPUT60), .C2(new_n839_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n822_), .A2(new_n830_), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n842_), .A2(new_n632_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n843_), .B2(new_n839_), .ZN(G1341gat));
  AOI21_X1  g643(.A(G127gat), .B1(new_n819_), .B2(new_n603_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT115), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n603_), .A2(G127gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n842_), .B2(new_n847_), .ZN(G1342gat));
  AOI21_X1  g647(.A(G134gat), .B1(new_n819_), .B2(new_n640_), .ZN(new_n849_));
  XOR2_X1   g648(.A(new_n849_), .B(KEYINPUT116), .Z(new_n850_));
  XNOR2_X1  g649(.A(KEYINPUT117), .B(G134gat), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n673_), .A2(new_n851_), .ZN(new_n852_));
  XOR2_X1   g651(.A(new_n852_), .B(KEYINPUT118), .Z(new_n853_));
  AOI21_X1  g652(.A(new_n850_), .B1(new_n842_), .B2(new_n853_), .ZN(G1343gat));
  NOR3_X1   g653(.A1(new_n451_), .A2(new_n322_), .A3(new_n379_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n812_), .A2(new_n432_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT119), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT119), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n812_), .A2(new_n858_), .A3(new_n432_), .A4(new_n855_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n857_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n504_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n632_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n860_), .B2(new_n603_), .ZN(new_n866_));
  AOI211_X1 g665(.A(KEYINPUT120), .B(new_n602_), .C1(new_n857_), .C2(new_n859_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT61), .B(G155gat), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OR3_X1    g668(.A1(new_n866_), .A2(new_n867_), .A3(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1346gat));
  INV_X1    g671(.A(G162gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n860_), .A2(new_n873_), .A3(new_n640_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n571_), .B1(new_n857_), .B2(new_n859_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n873_), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(KEYINPUT121), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT121), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n874_), .B(new_n878_), .C1(new_n873_), .C2(new_n875_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1347gat));
  XOR2_X1   g679(.A(new_n768_), .B(KEYINPUT54), .Z(new_n881_));
  INV_X1    g680(.A(KEYINPUT112), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n811_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n883_), .B2(new_n823_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n322_), .A2(new_n379_), .A3(new_n431_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n416_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT123), .B1(new_n884_), .B2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT123), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n829_), .A2(new_n889_), .A3(new_n886_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n888_), .A2(new_n890_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(new_n504_), .A3(new_n268_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n885_), .A2(new_n505_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT122), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n451_), .ZN(new_n895_));
  OAI21_X1  g694(.A(G169gat), .B1(new_n884_), .B2(new_n895_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT62), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n892_), .A2(new_n897_), .ZN(G1348gat));
  NAND3_X1  g697(.A1(new_n888_), .A2(new_n890_), .A3(new_n632_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n900_));
  AND3_X1   g699(.A1(new_n899_), .A2(new_n900_), .A3(new_n253_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n899_), .B2(new_n253_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n887_), .B1(new_n769_), .B2(new_n811_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n903_), .A2(G176gat), .A3(new_n632_), .ZN(new_n904_));
  XOR2_X1   g703(.A(new_n904_), .B(KEYINPUT125), .Z(new_n905_));
  NOR3_X1   g704(.A1(new_n901_), .A2(new_n902_), .A3(new_n905_), .ZN(G1349gat));
  AOI21_X1  g705(.A(G183gat), .B1(new_n903_), .B2(new_n603_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n602_), .A2(new_n232_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n891_), .B2(new_n908_), .ZN(G1350gat));
  NAND3_X1  g708(.A1(new_n888_), .A2(new_n890_), .A3(new_n673_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(G190gat), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n888_), .A2(new_n890_), .A3(new_n233_), .A4(new_n640_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT126), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n911_), .A2(new_n915_), .A3(new_n912_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1351gat));
  NOR3_X1   g716(.A1(new_n451_), .A2(new_n380_), .A3(new_n321_), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n812_), .A2(new_n432_), .A3(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n919_), .A2(new_n504_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g720(.A1(new_n919_), .A2(new_n632_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g722(.A1(new_n919_), .A2(new_n603_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n926_), .B(KEYINPUT127), .Z(new_n927_));
  AND2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n924_), .A2(new_n925_), .A3(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1354gat));
  INV_X1    g729(.A(new_n919_), .ZN(new_n931_));
  OAI21_X1  g730(.A(G218gat), .B1(new_n931_), .B2(new_n571_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n919_), .A2(new_n223_), .A3(new_n640_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1355gat));
endmodule


