//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n756_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_;
  INV_X1    g000(.A(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  AOI211_X1 g002(.A(KEYINPUT68), .B(KEYINPUT7), .C1(new_n202_), .C2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n208_));
  NAND4_X1  g007(.A1(new_n207_), .A2(new_n202_), .A3(new_n203_), .A4(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n205_), .A2(KEYINPUT69), .A3(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT6), .B1(new_n202_), .B2(new_n203_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT69), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n208_), .A2(new_n202_), .A3(new_n203_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(new_n206_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n217_), .B2(new_n204_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n210_), .A2(new_n214_), .A3(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G85gat), .B(G92gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(KEYINPUT8), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT67), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n214_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT67), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XOR2_X1   g025(.A(KEYINPUT10), .B(G99gat), .Z(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(new_n203_), .ZN(new_n228_));
  INV_X1    g027(.A(G92gat), .ZN(new_n229_));
  OR2_X1    g028(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT65), .B1(new_n232_), .B2(KEYINPUT9), .ZN(new_n233_));
  NAND3_X1  g032(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(KEYINPUT66), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n236_), .B1(G85gat), .B2(G92gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n235_), .B1(new_n234_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  NOR3_X1   g038(.A1(new_n232_), .A2(KEYINPUT65), .A3(KEYINPUT9), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n226_), .B(new_n228_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT8), .ZN(new_n242_));
  AOI22_X1  g041(.A1(new_n224_), .A2(new_n225_), .B1(new_n205_), .B2(new_n209_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n242_), .B1(new_n243_), .B2(new_n220_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n222_), .A2(new_n241_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT71), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n222_), .A2(new_n241_), .A3(new_n244_), .A4(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G57gat), .B(G64gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G71gat), .B(G78gat), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n251_), .A3(KEYINPUT11), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n253_));
  INV_X1    g052(.A(new_n251_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n252_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT12), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n249_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n257_), .B(KEYINPUT70), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n245_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT12), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n245_), .A2(new_n261_), .ZN(new_n265_));
  AND2_X1   g064(.A1(G230gat), .A2(G233gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n260_), .A2(KEYINPUT72), .A3(new_n264_), .A4(new_n267_), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n267_), .B(new_n264_), .C1(new_n249_), .C2(new_n259_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n262_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n266_), .B1(new_n273_), .B2(new_n265_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G120gat), .B(G148gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT5), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G176gat), .B(G204gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n279_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n272_), .A2(new_n274_), .A3(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT13), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n280_), .A2(KEYINPUT13), .A3(new_n282_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT77), .B(G15gat), .ZN(new_n288_));
  INV_X1    g087(.A(G22gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n288_), .B(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G1gat), .ZN(new_n291_));
  INV_X1    g090(.A(G8gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT14), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G1gat), .B(G8gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G29gat), .B(G36gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT73), .ZN(new_n298_));
  AND2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n297_), .A2(new_n298_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G43gat), .B(G50gat), .Z(new_n301_));
  OR3_X1    g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n301_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n296_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G229gat), .A2(G233gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT15), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n304_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n296_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n296_), .A2(new_n304_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n306_), .A3(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n308_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G113gat), .B(G141gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G169gat), .B(G197gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n315_), .B(new_n316_), .Z(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT82), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n314_), .A2(KEYINPUT82), .A3(new_n317_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n314_), .A2(new_n317_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT83), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n287_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT2), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT93), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT93), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n328_), .A2(new_n332_), .A3(new_n329_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT94), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n334_), .A2(new_n337_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT92), .ZN(new_n343_));
  INV_X1    g142(.A(G155gat), .ZN(new_n344_));
  INV_X1    g143(.A(G162gat), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(KEYINPUT92), .B1(G155gat), .B2(G162gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT95), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT95), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n348_), .A2(new_n352_), .A3(new_n349_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n342_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT1), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n349_), .B(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n348_), .ZN(new_n357_));
  OR3_X1    g156(.A1(KEYINPUT91), .A2(G141gat), .A3(G148gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT91), .B1(G141gat), .B2(G148gat), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n358_), .A2(new_n359_), .A3(new_n328_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n354_), .A2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT28), .B1(new_n362_), .B2(KEYINPUT29), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n348_), .A2(new_n352_), .A3(new_n349_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n352_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n366_), .A2(new_n342_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT28), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT29), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n372_), .B(KEYINPUT96), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n371_), .B(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n369_), .B1(new_n354_), .B2(new_n361_), .ZN(new_n375_));
  XOR2_X1   g174(.A(G211gat), .B(G218gat), .Z(new_n376_));
  INV_X1    g175(.A(KEYINPUT21), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G197gat), .B(G204gat), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n378_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT21), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n380_), .A2(new_n376_), .A3(KEYINPUT21), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(G78gat), .B1(new_n375_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(G78gat), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n387_), .B(new_n384_), .C1(new_n367_), .C2(new_n369_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n388_), .A3(G106gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(G106gat), .B1(new_n386_), .B2(new_n388_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G22gat), .B(G50gat), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n392_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n386_), .A2(new_n388_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n203_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n394_), .B1(new_n396_), .B2(new_n389_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n374_), .B1(new_n393_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n374_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n392_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(new_n389_), .A3(new_n394_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G85gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT0), .B(G57gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G127gat), .B(G134gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G113gat), .B(G120gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n354_), .A2(new_n361_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT99), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n409_), .A2(new_n410_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n414_), .A2(KEYINPUT89), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n415_), .B1(new_n411_), .B2(KEYINPUT89), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n362_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G225gat), .A2(G233gat), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT99), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n354_), .A2(new_n419_), .A3(new_n361_), .A4(new_n411_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n413_), .A2(new_n417_), .A3(new_n418_), .A4(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT4), .B1(new_n362_), .B2(new_n416_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n413_), .A2(new_n417_), .A3(new_n420_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n422_), .B1(new_n423_), .B2(KEYINPUT4), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n408_), .B(new_n421_), .C1(new_n424_), .C2(new_n418_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT100), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT33), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(KEYINPUT100), .A3(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(G8gat), .B(G36gat), .Z(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G64gat), .B(G92gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G226gat), .A2(G233gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT19), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n438_));
  NOR2_X1   g237(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(G169gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G183gat), .A2(G190gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT23), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(KEYINPUT87), .A2(KEYINPUT23), .ZN(new_n444_));
  NOR2_X1   g243(.A1(KEYINPUT87), .A2(KEYINPUT23), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n443_), .B1(new_n446_), .B2(new_n441_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(G183gat), .A2(G190gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n440_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT86), .ZN(new_n450_));
  INV_X1    g249(.A(G183gat), .ZN(new_n451_));
  AOI21_X1  g250(.A(KEYINPUT84), .B1(new_n451_), .B2(KEYINPUT25), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(KEYINPUT25), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT26), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n456_), .A3(G190gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n451_), .A2(KEYINPUT84), .A3(KEYINPUT25), .ZN(new_n458_));
  INV_X1    g257(.A(G190gat), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT26), .B1(new_n459_), .B2(KEYINPUT85), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n454_), .A2(new_n457_), .A3(new_n458_), .A4(new_n460_), .ZN(new_n461_));
  OR2_X1    g260(.A1(G169gat), .A2(G176gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G169gat), .A2(G176gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(KEYINPUT24), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n450_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n460_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT84), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT25), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n467_), .B1(new_n468_), .B2(G183gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(G183gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n450_), .B(new_n464_), .C1(new_n466_), .C2(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n462_), .A2(KEYINPUT24), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n441_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n442_), .A2(G183gat), .A3(G190gat), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n449_), .B1(new_n465_), .B2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n438_), .B1(new_n478_), .B2(new_n384_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n462_), .A2(KEYINPUT24), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n451_), .A2(KEYINPUT25), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n470_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT26), .B(G190gat), .Z(new_n483_));
  OAI211_X1 g282(.A(new_n480_), .B(new_n464_), .C1(new_n482_), .C2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT97), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n463_), .B(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(KEYINPUT22), .B(G169gat), .Z(new_n487_));
  OAI21_X1  g286(.A(new_n486_), .B1(G176gat), .B2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n448_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n489_));
  OAI22_X1  g288(.A1(new_n484_), .A2(new_n447_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n384_), .A2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n437_), .B1(new_n479_), .B2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n438_), .B1(new_n384_), .B2(new_n490_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n493_), .B(new_n437_), .C1(new_n384_), .C2(new_n478_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n435_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n478_), .A2(new_n384_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n497_), .A2(new_n491_), .A3(KEYINPUT20), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n494_), .B(new_n434_), .C1(new_n498_), .C2(new_n437_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n407_), .B1(new_n423_), .B2(new_n418_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n423_), .A2(KEYINPUT4), .ZN(new_n502_));
  INV_X1    g301(.A(new_n422_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n501_), .B1(new_n504_), .B2(new_n418_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n500_), .A2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n427_), .A2(new_n429_), .A3(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n421_), .B1(new_n424_), .B2(new_n418_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n407_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n425_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n494_), .B1(new_n498_), .B2(new_n437_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n435_), .A2(KEYINPUT32), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n437_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT101), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n384_), .B1(new_n490_), .B2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n516_), .B1(new_n515_), .B2(new_n490_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n514_), .B1(new_n517_), .B2(new_n479_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n493_), .B1(new_n384_), .B2(new_n478_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n519_), .A2(new_n437_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n521_), .A2(new_n512_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n510_), .A2(new_n513_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n403_), .B1(new_n507_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n510_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n434_), .B1(new_n518_), .B2(new_n520_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT27), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n527_), .B1(new_n511_), .B2(new_n435_), .ZN(new_n528_));
  AOI22_X1  g327(.A1(new_n526_), .A2(new_n528_), .B1(new_n500_), .B2(new_n527_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n403_), .A2(new_n525_), .A3(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT88), .B(G43gat), .Z(new_n531_));
  OAI211_X1 g330(.A(new_n449_), .B(KEYINPUT30), .C1(new_n465_), .C2(new_n477_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n464_), .B1(new_n466_), .B2(new_n471_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT86), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n535_), .A2(new_n472_), .A3(new_n476_), .ZN(new_n536_));
  AOI21_X1  g335(.A(KEYINPUT30), .B1(new_n536_), .B2(new_n449_), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n533_), .A2(new_n537_), .A3(G99gat), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT30), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n478_), .A2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n202_), .B1(new_n540_), .B2(new_n532_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n531_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G227gat), .A2(G233gat), .ZN(new_n543_));
  INV_X1    g342(.A(G15gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(G71gat), .ZN(new_n546_));
  OAI21_X1  g345(.A(G99gat), .B1(new_n533_), .B2(new_n537_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n531_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n540_), .A2(new_n202_), .A3(new_n532_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n547_), .A2(new_n548_), .A3(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n542_), .A2(new_n546_), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT90), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n546_), .B1(new_n542_), .B2(new_n550_), .ZN(new_n553_));
  OAI21_X1  g352(.A(KEYINPUT31), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n542_), .A2(new_n550_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n546_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT31), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n557_), .A2(new_n551_), .A3(KEYINPUT90), .A4(new_n558_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n554_), .A2(new_n416_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n416_), .B1(new_n554_), .B2(new_n559_), .ZN(new_n561_));
  OAI22_X1  g360(.A1(new_n524_), .A2(new_n530_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n554_), .A2(new_n559_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n416_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n554_), .A2(new_n416_), .A3(new_n559_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n528_), .A2(new_n526_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n500_), .A2(new_n527_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n403_), .A2(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n565_), .A2(new_n525_), .A3(new_n566_), .A4(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n562_), .A2(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n327_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n310_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n245_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n304_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT35), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT34), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n575_), .A2(new_n576_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n577_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n574_), .A2(new_n581_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n583_), .B1(new_n574_), .B2(new_n581_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G190gat), .B(G218gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT74), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G134gat), .B(G162gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT36), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n592_), .B(KEYINPUT75), .Z(new_n593_));
  NAND2_X1  g392(.A1(new_n586_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n590_), .B(KEYINPUT36), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n594_), .A2(new_n596_), .A3(KEYINPUT37), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT76), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n574_), .A2(new_n581_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(new_n582_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n574_), .A2(new_n581_), .A3(new_n583_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n598_), .B1(new_n602_), .B2(new_n595_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n598_), .B(new_n595_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n594_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT37), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n597_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(G127gat), .B(G155gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(KEYINPUT79), .B(KEYINPUT16), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G183gat), .B(G211gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT17), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT80), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n296_), .B(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n261_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n617_), .A2(new_n261_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n257_), .B(KEYINPUT78), .Z(new_n621_));
  NOR2_X1   g420(.A1(new_n617_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(new_n621_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT17), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n613_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  OAI22_X1  g425(.A1(new_n619_), .A2(new_n620_), .B1(new_n622_), .B2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT81), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n608_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n573_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n510_), .B(KEYINPUT102), .Z(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n291_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n633_), .B1(KEYINPUT104), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT104), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n635_), .B1(new_n636_), .B2(KEYINPUT38), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n322_), .A2(new_n323_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n287_), .A2(new_n627_), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n606_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n562_), .B2(new_n571_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT103), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n525_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n633_), .A2(KEYINPUT104), .A3(new_n634_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n637_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n646_), .B(new_n647_), .ZN(G1324gat));
  AOI21_X1  g447(.A(new_n292_), .B1(new_n642_), .B2(new_n569_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n649_), .A2(new_n650_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n631_), .A2(new_n292_), .A3(new_n569_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(G1325gat));
  NOR2_X1   g456(.A1(new_n560_), .A2(new_n561_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n631_), .A2(new_n544_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n658_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G15gat), .B1(new_n643_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT41), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n661_), .A2(new_n662_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n659_), .B1(new_n663_), .B2(new_n664_), .ZN(G1326gat));
  NAND3_X1  g464(.A1(new_n631_), .A2(new_n289_), .A3(new_n403_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n403_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G22gat), .B1(new_n643_), .B2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n668_), .A2(KEYINPUT42), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(KEYINPUT42), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(G1327gat));
  NOR3_X1   g470(.A1(new_n287_), .A2(new_n638_), .A3(new_n628_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT43), .ZN(new_n673_));
  INV_X1    g472(.A(new_n608_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n572_), .B2(new_n674_), .ZN(new_n675_));
  AOI211_X1 g474(.A(KEYINPUT43), .B(new_n608_), .C1(new_n562_), .C2(new_n571_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT44), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n672_), .B(KEYINPUT44), .C1(new_n675_), .C2(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n632_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G29gat), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n628_), .A2(new_n606_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n573_), .A2(new_n684_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n525_), .A2(G29gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n683_), .B1(new_n685_), .B2(new_n686_), .ZN(G1328gat));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n529_), .A2(G36gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n573_), .A2(new_n684_), .A3(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT45), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n679_), .A2(new_n694_), .A3(new_n569_), .A4(new_n680_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(G36gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n679_), .A2(new_n569_), .A3(new_n680_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT108), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n693_), .B1(new_n696_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT109), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n688_), .B(new_n689_), .C1(new_n699_), .C2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT46), .B1(new_n699_), .B2(new_n688_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n691_), .B(KEYINPUT45), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n697_), .A2(KEYINPUT108), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n695_), .A2(G36gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n703_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT110), .B1(new_n706_), .B2(KEYINPUT109), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n701_), .B1(new_n702_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(G1329gat));
  OAI21_X1  g508(.A(G43gat), .B1(new_n681_), .B2(new_n660_), .ZN(new_n710_));
  OR2_X1    g509(.A1(new_n660_), .A2(G43gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n710_), .B1(new_n685_), .B2(new_n711_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT47), .Z(G1330gat));
  INV_X1    g512(.A(G50gat), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n681_), .A2(new_n714_), .A3(new_n667_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n573_), .A2(new_n403_), .A3(new_n684_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n714_), .B2(new_n716_), .ZN(G1331gat));
  INV_X1    g516(.A(new_n286_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT13), .B1(new_n280_), .B2(new_n282_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(new_n629_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n721_), .A2(KEYINPUT111), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n324_), .B1(new_n562_), .B2(new_n571_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(KEYINPUT111), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n722_), .A2(new_n723_), .A3(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G57gat), .B1(new_n726_), .B2(new_n632_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n326_), .A2(new_n628_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(new_n641_), .A3(new_n287_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT112), .B(G57gat), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n730_), .A2(new_n525_), .A3(new_n731_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n727_), .A2(new_n732_), .ZN(G1332gat));
  OAI21_X1  g532(.A(G64gat), .B1(new_n730_), .B2(new_n529_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT48), .ZN(new_n735_));
  OR2_X1    g534(.A1(new_n529_), .A2(G64gat), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n725_), .B2(new_n736_), .ZN(G1333gat));
  OAI21_X1  g536(.A(G71gat), .B1(new_n730_), .B2(new_n660_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT49), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n660_), .A2(G71gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n725_), .B2(new_n740_), .ZN(G1334gat));
  OAI21_X1  g540(.A(G78gat), .B1(new_n730_), .B2(new_n667_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT50), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n726_), .A2(new_n387_), .A3(new_n403_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1335gat));
  AND3_X1   g544(.A1(new_n723_), .A2(new_n287_), .A3(new_n684_), .ZN(new_n746_));
  AOI21_X1  g545(.A(G85gat), .B1(new_n746_), .B2(new_n632_), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n675_), .A2(new_n676_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n720_), .A2(new_n324_), .A3(new_n628_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n525_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n747_), .B1(new_n751_), .B2(new_n752_), .ZN(G1336gat));
  NAND3_X1  g552(.A1(new_n746_), .A2(new_n229_), .A3(new_n569_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n751_), .A2(new_n569_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n756_), .B2(new_n229_), .ZN(G1337gat));
  NAND3_X1  g556(.A1(new_n746_), .A2(new_n658_), .A3(new_n227_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT113), .Z(new_n759_));
  OAI21_X1  g558(.A(G99gat), .B1(new_n750_), .B2(new_n660_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n759_), .A2(new_n760_), .B1(KEYINPUT114), .B2(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n761_), .A2(KEYINPUT114), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(G1338gat));
  NAND3_X1  g563(.A1(new_n746_), .A2(new_n203_), .A3(new_n403_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G106gat), .B1(new_n750_), .B2(new_n667_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n766_), .A2(KEYINPUT52), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(KEYINPUT52), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n765_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT53), .ZN(G1339gat));
  AND2_X1   g569(.A1(new_n658_), .A2(new_n570_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n632_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT57), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT56), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n281_), .A2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n268_), .A2(new_n271_), .A3(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n269_), .ZN(new_n779_));
  OAI221_X1 g578(.A(new_n264_), .B1(new_n245_), .B2(new_n261_), .C1(new_n249_), .C2(new_n259_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n779_), .A2(KEYINPUT55), .B1(new_n780_), .B2(new_n266_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n776_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n782_), .A2(KEYINPUT115), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(KEYINPUT115), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n281_), .B1(new_n778_), .B2(new_n781_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n783_), .B(new_n784_), .C1(KEYINPUT56), .C2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n324_), .A2(new_n282_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n311_), .A2(new_n312_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n306_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(new_n789_), .B2(new_n788_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n317_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT117), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n791_), .A2(KEYINPUT117), .A3(new_n792_), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n322_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  AOI22_X1  g596(.A1(new_n786_), .A2(new_n787_), .B1(new_n283_), .B2(new_n797_), .ZN(new_n798_));
  OAI211_X1 g597(.A(KEYINPUT118), .B(new_n773_), .C1(new_n798_), .C2(new_n640_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n800_));
  OAI22_X1  g599(.A1(KEYINPUT115), .A2(new_n782_), .B1(new_n785_), .B2(KEYINPUT56), .ZN(new_n801_));
  INV_X1    g600(.A(new_n784_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n787_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n283_), .A2(new_n797_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n640_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n800_), .B1(new_n805_), .B2(KEYINPUT57), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(KEYINPUT57), .ZN(new_n807_));
  AND4_X1   g606(.A1(new_n322_), .A2(new_n282_), .A3(new_n795_), .A4(new_n796_), .ZN(new_n808_));
  OAI22_X1  g607(.A1(KEYINPUT119), .A2(new_n782_), .B1(new_n785_), .B2(KEYINPUT56), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n782_), .A2(KEYINPUT119), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n808_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n608_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n813_), .B1(new_n812_), .B2(new_n811_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n799_), .A2(new_n806_), .A3(new_n807_), .A4(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n627_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n720_), .A2(new_n628_), .A3(new_n326_), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT54), .B1(new_n817_), .B2(new_n674_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT54), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n729_), .A2(new_n720_), .A3(new_n819_), .A4(new_n608_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n772_), .B1(new_n816_), .B2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(G113gat), .B1(new_n823_), .B2(new_n324_), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n824_), .A2(KEYINPUT120), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(KEYINPUT120), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n821_), .B1(new_n815_), .B2(new_n627_), .ZN(new_n827_));
  OAI21_X1  g626(.A(KEYINPUT59), .B1(new_n827_), .B2(new_n772_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n772_), .A2(KEYINPUT59), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n814_), .A2(new_n807_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n773_), .B1(new_n798_), .B2(new_n640_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n628_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n829_), .B1(new_n832_), .B2(new_n821_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n828_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(G113gat), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n326_), .A2(new_n835_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n825_), .A2(new_n826_), .B1(new_n834_), .B2(new_n836_), .ZN(G1340gat));
  NAND3_X1  g636(.A1(new_n828_), .A2(new_n287_), .A3(new_n833_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT122), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n828_), .A2(new_n840_), .A3(new_n287_), .A4(new_n833_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(G120gat), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT60), .ZN(new_n843_));
  AOI21_X1  g642(.A(G120gat), .B1(new_n287_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n843_), .B2(G120gat), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n823_), .A2(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT121), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n842_), .A2(new_n847_), .ZN(G1341gat));
  AOI21_X1  g647(.A(G127gat), .B1(new_n823_), .B2(new_n628_), .ZN(new_n849_));
  OR2_X1    g648(.A1(new_n849_), .A2(KEYINPUT123), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(KEYINPUT123), .ZN(new_n851_));
  INV_X1    g650(.A(G127gat), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n627_), .A2(new_n852_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n850_), .A2(new_n851_), .B1(new_n834_), .B2(new_n853_), .ZN(G1342gat));
  NAND3_X1  g653(.A1(new_n828_), .A2(new_n674_), .A3(new_n833_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(G134gat), .ZN(new_n856_));
  INV_X1    g655(.A(new_n823_), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n606_), .A2(G134gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n856_), .B1(new_n857_), .B2(new_n858_), .ZN(G1343gat));
  NAND2_X1  g658(.A1(new_n816_), .A2(new_n822_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT125), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n660_), .A2(new_n403_), .A3(new_n529_), .A4(new_n632_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT124), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n860_), .A2(new_n861_), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n863_), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT125), .B1(new_n827_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT126), .B(G141gat), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n867_), .A2(new_n324_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n867_), .B2(new_n324_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1344gat));
  INV_X1    g670(.A(new_n867_), .ZN(new_n872_));
  OAI21_X1  g671(.A(G148gat), .B1(new_n872_), .B2(new_n720_), .ZN(new_n873_));
  INV_X1    g672(.A(G148gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n867_), .A2(new_n874_), .A3(new_n287_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1345gat));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  INV_X1    g676(.A(new_n628_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n872_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n877_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n867_), .A2(new_n628_), .A3(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n879_), .A2(new_n881_), .ZN(G1346gat));
  OAI21_X1  g681(.A(G162gat), .B1(new_n872_), .B2(new_n608_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n867_), .A2(new_n345_), .A3(new_n640_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1347gat));
  NOR2_X1   g684(.A1(new_n832_), .A2(new_n821_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n660_), .A2(new_n529_), .A3(new_n632_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n667_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n886_), .A2(new_n638_), .A3(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n890_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n892_));
  INV_X1    g691(.A(G169gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n889_), .B2(new_n893_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n891_), .B(new_n894_), .C1(new_n487_), .C2(new_n890_), .ZN(G1348gat));
  NOR2_X1   g694(.A1(new_n886_), .A2(new_n888_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G176gat), .B1(new_n896_), .B2(new_n287_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n827_), .A2(new_n403_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n887_), .A2(G176gat), .A3(new_n287_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(G1349gat));
  NAND3_X1  g699(.A1(new_n898_), .A2(new_n628_), .A3(new_n887_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n627_), .B1(new_n470_), .B2(new_n481_), .ZN(new_n902_));
  AOI22_X1  g701(.A1(new_n901_), .A2(new_n451_), .B1(new_n896_), .B2(new_n902_), .ZN(G1350gat));
  INV_X1    g702(.A(new_n483_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n896_), .A2(new_n904_), .A3(new_n640_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n886_), .A2(new_n608_), .A3(new_n888_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n459_), .ZN(G1351gat));
  NOR4_X1   g706(.A1(new_n658_), .A2(new_n510_), .A3(new_n667_), .A4(new_n529_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n860_), .A2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n324_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g711(.A1(new_n909_), .A2(new_n720_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(KEYINPUT127), .B(G204gat), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n913_), .B(new_n914_), .ZN(G1353gat));
  NOR2_X1   g714(.A1(new_n909_), .A2(new_n627_), .ZN(new_n916_));
  OR2_X1    g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n916_), .A2(new_n917_), .ZN(new_n918_));
  XOR2_X1   g717(.A(KEYINPUT63), .B(G211gat), .Z(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n916_), .B2(new_n919_), .ZN(G1354gat));
  OR3_X1    g719(.A1(new_n909_), .A2(G218gat), .A3(new_n606_), .ZN(new_n921_));
  OAI21_X1  g720(.A(G218gat), .B1(new_n909_), .B2(new_n608_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1355gat));
endmodule


