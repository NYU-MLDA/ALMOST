//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n584_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n594_,
    new_n595_, new_n596_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n860_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_;
  INV_X1    g000(.A(KEYINPUT93), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT26), .B(G190gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT78), .B(G183gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT25), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n203_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G183gat), .ZN(new_n209_));
  INV_X1    g008(.A(G190gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT23), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(KEYINPUT24), .A3(new_n218_), .ZN(new_n219_));
  OR3_X1    g018(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n214_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n208_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n204_), .A2(new_n210_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(new_n214_), .ZN(new_n224_));
  OAI21_X1  g023(.A(KEYINPUT79), .B1(new_n215_), .B2(KEYINPUT22), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT22), .B(G169gat), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n216_), .B(new_n225_), .C1(new_n226_), .C2(KEYINPUT79), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n227_), .A3(new_n218_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n222_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G197gat), .B(G204gat), .ZN(new_n230_));
  XOR2_X1   g029(.A(G211gat), .B(G218gat), .Z(new_n231_));
  INV_X1    g030(.A(KEYINPUT21), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n233_), .B1(new_n232_), .B2(new_n231_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n231_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(new_n230_), .A3(KEYINPUT21), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n229_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT20), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G226gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT19), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n214_), .B1(G183gat), .B2(G190gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n226_), .A2(new_n216_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n218_), .A3(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT25), .B(G183gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n203_), .A2(new_n246_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n247_), .A2(new_n214_), .A3(new_n219_), .A4(new_n220_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n242_), .B1(new_n237_), .B2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n239_), .A2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT20), .B1(new_n229_), .B2(new_n237_), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n252_), .A2(KEYINPUT87), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n252_), .A2(KEYINPUT87), .B1(new_n237_), .B2(new_n249_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n251_), .B1(new_n255_), .B2(new_n241_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G8gat), .B(G36gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(G64gat), .B(G92gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n256_), .A2(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n242_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n261_), .B1(new_n264_), .B2(new_n251_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT27), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n267_), .B1(new_n256_), .B2(new_n262_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n249_), .A2(KEYINPUT91), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n249_), .A2(KEYINPUT91), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n237_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n241_), .B1(new_n272_), .B2(new_n239_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(new_n255_), .B2(new_n241_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n261_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n268_), .A2(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(G127gat), .B(G134gat), .Z(new_n278_));
  XOR2_X1   g077(.A(G113gat), .B(G120gat), .Z(new_n279_));
  OR2_X1    g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n280_), .A2(KEYINPUT81), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(KEYINPUT81), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n278_), .A2(new_n279_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G155gat), .B(G162gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT84), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT2), .ZN(new_n288_));
  OAI22_X1  g087(.A1(KEYINPUT83), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n292_), .A2(KEYINPUT83), .A3(KEYINPUT3), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n288_), .A2(new_n291_), .A3(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n286_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(G155gat), .ZN(new_n296_));
  INV_X1    g095(.A(G162gat), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT1), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n298_), .B1(G155gat), .B2(G162gat), .ZN(new_n299_));
  NOR3_X1   g098(.A1(new_n296_), .A2(new_n297_), .A3(KEYINPUT1), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n287_), .B(new_n292_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n295_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n284_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n280_), .A2(new_n283_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n295_), .A2(new_n306_), .A3(new_n301_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n308_));
  OAI211_X1 g107(.A(KEYINPUT4), .B(new_n307_), .C1(new_n308_), .C2(new_n302_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G225gat), .A2(G233gat), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n310_), .B(KEYINPUT89), .Z(new_n311_));
  NAND3_X1  g110(.A1(new_n305_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n284_), .A2(new_n303_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(new_n307_), .A3(new_n310_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G1gat), .B(G29gat), .Z(new_n315_));
  XNOR2_X1  g114(.A(G57gat), .B(G85gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT90), .B(KEYINPUT0), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n312_), .A2(new_n314_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT92), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT92), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n312_), .A2(new_n314_), .A3(new_n322_), .A4(new_n319_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n312_), .A2(new_n314_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n319_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n321_), .A2(new_n323_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT29), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n302_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT28), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n237_), .A2(KEYINPUT86), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n329_), .B1(new_n295_), .B2(new_n301_), .ZN(new_n334_));
  OAI211_X1 g133(.A(G228gat), .B(G233gat), .C1(new_n333_), .C2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G228gat), .A2(G233gat), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT86), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n337_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n336_), .B(new_n338_), .C1(new_n302_), .C2(new_n329_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G78gat), .B(G106gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n335_), .A2(new_n339_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n341_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n332_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n335_), .A2(new_n339_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n340_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n330_), .B(KEYINPUT28), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n342_), .A3(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G22gat), .B(G50gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT85), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n345_), .A2(new_n349_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n351_), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n343_), .A2(new_n332_), .A3(new_n344_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n348_), .B1(new_n347_), .B2(new_n342_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n328_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n202_), .B1(new_n277_), .B2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n274_), .A2(KEYINPUT32), .A3(new_n262_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT32), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n256_), .B1(new_n360_), .B2(new_n261_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n327_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n320_), .A2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n312_), .A2(new_n314_), .A3(KEYINPUT33), .A4(new_n319_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n305_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n313_), .A2(new_n307_), .A3(new_n311_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(new_n367_), .A3(new_n325_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n364_), .A2(new_n365_), .A3(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n362_), .B1(new_n266_), .B2(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n356_), .A2(new_n352_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n266_), .A2(new_n267_), .B1(new_n269_), .B2(new_n275_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n374_), .A2(new_n371_), .A3(KEYINPUT93), .A4(new_n328_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n358_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n229_), .B(KEYINPUT30), .ZN(new_n377_));
  XOR2_X1   g176(.A(G71gat), .B(G99gat), .Z(new_n378_));
  NAND2_X1  g177(.A1(G227gat), .A2(G233gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n378_), .B(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G15gat), .B(G43gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT80), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n380_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n377_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(new_n308_), .ZN(new_n385_));
  XOR2_X1   g184(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n269_), .A2(new_n275_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT27), .B1(new_n263_), .B2(new_n265_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT94), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT94), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n268_), .A2(new_n391_), .A3(new_n276_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n371_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n387_), .A2(new_n327_), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n376_), .A2(new_n387_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  XOR2_X1   g194(.A(G43gat), .B(G50gat), .Z(new_n396_));
  XNOR2_X1  g195(.A(G29gat), .B(G36gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT15), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT9), .ZN(new_n401_));
  INV_X1    g200(.A(G85gat), .ZN(new_n402_));
  INV_X1    g201(.A(G92gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G85gat), .A2(G92gat), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n401_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT64), .ZN(new_n407_));
  AOI21_X1  g206(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n408_));
  OR3_X1    g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n410_));
  XOR2_X1   g209(.A(KEYINPUT10), .B(G99gat), .Z(new_n411_));
  INV_X1    g210(.A(G106gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G99gat), .A2(G106gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT6), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(G99gat), .A3(G106gat), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n411_), .A2(new_n412_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n409_), .A2(new_n410_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT8), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n414_), .A2(new_n416_), .ZN(new_n420_));
  AND2_X1   g219(.A1(KEYINPUT66), .A2(KEYINPUT67), .ZN(new_n421_));
  NOR2_X1   g220(.A1(KEYINPUT66), .A2(KEYINPUT67), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(new_n414_), .B(new_n416_), .C1(new_n422_), .C2(new_n421_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT65), .ZN(new_n426_));
  INV_X1    g225(.A(G99gat), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n412_), .A4(KEYINPUT7), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT7), .ZN(new_n429_));
  OAI22_X1  g228(.A1(new_n429_), .A2(KEYINPUT65), .B1(G99gat), .B2(G106gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n426_), .A2(KEYINPUT7), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n428_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n424_), .A2(new_n425_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n404_), .A2(new_n405_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n419_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n436_));
  AOI211_X1 g235(.A(KEYINPUT8), .B(new_n434_), .C1(new_n432_), .C2(new_n420_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n418_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n400_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G232gat), .A2(G233gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT34), .ZN(new_n441_));
  OR2_X1    g240(.A1(new_n441_), .A2(KEYINPUT35), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n439_), .B(new_n442_), .C1(new_n438_), .C2(new_n398_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n441_), .A2(KEYINPUT35), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n443_), .B(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT36), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G190gat), .B(G218gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT71), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT72), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G134gat), .B(G162gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n445_), .A2(new_n446_), .A3(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n446_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n445_), .A2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n452_), .A2(new_n454_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n395_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G71gat), .B(G78gat), .Z(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G57gat), .B(G64gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT68), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G57gat), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n462_), .A2(G64gat), .ZN(new_n463_));
  INV_X1    g262(.A(G64gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n464_), .A2(G57gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT68), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n461_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n458_), .B1(new_n467_), .B2(KEYINPUT11), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT11), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n461_), .A2(new_n466_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  AOI211_X1 g270(.A(new_n469_), .B(new_n457_), .C1(new_n461_), .C2(new_n466_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n474_), .B(new_n418_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n472_), .B1(new_n470_), .B2(new_n468_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n438_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n475_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(G230gat), .A3(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT12), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G230gat), .A2(G233gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n438_), .A2(KEYINPUT12), .A3(new_n476_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n475_), .A4(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G120gat), .B(G148gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT5), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G176gat), .B(G204gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n479_), .A2(new_n484_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n488_), .B(KEYINPUT69), .Z(new_n491_));
  AOI21_X1  g290(.A(new_n491_), .B1(new_n479_), .B2(new_n484_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT13), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(KEYINPUT70), .A3(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n495_), .A2(KEYINPUT70), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(KEYINPUT70), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n493_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n496_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G15gat), .B(G22gat), .ZN(new_n501_));
  INV_X1    g300(.A(G1gat), .ZN(new_n502_));
  INV_X1    g301(.A(G8gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT14), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G1gat), .B(G8gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  OR2_X1    g306(.A1(new_n507_), .A2(new_n398_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n398_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT76), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(KEYINPUT76), .A3(new_n509_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT77), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(KEYINPUT77), .A3(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n400_), .A2(new_n507_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(new_n514_), .A3(new_n508_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n518_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G113gat), .B(G141gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G169gat), .B(G197gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n523_), .B(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n525_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n518_), .A2(new_n519_), .A3(new_n521_), .A4(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n500_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G231gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n507_), .B(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(new_n474_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G127gat), .B(G155gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT16), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT17), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n535_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n539_), .B(new_n540_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n535_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT74), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n545_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n532_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n456_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT96), .ZN(new_n552_));
  OAI21_X1  g351(.A(G1gat), .B1(new_n552_), .B2(new_n328_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n395_), .A2(new_n532_), .ZN(new_n554_));
  OR3_X1    g353(.A1(new_n452_), .A2(new_n454_), .A3(KEYINPUT73), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT37), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT75), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n548_), .B(new_n558_), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n554_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT95), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n327_), .A2(new_n502_), .ZN(new_n563_));
  OR3_X1    g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT38), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n562_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n566_));
  AND3_X1   g365(.A1(new_n564_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n565_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n553_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT97), .ZN(G1324gat));
  NAND2_X1  g369(.A1(new_n390_), .A2(new_n392_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n456_), .A2(new_n572_), .A3(new_n550_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT98), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n573_), .A2(new_n574_), .A3(G8gat), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n574_), .B1(new_n573_), .B2(G8gat), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT39), .ZN(new_n577_));
  OR3_X1    g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n577_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n572_), .A2(new_n503_), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n578_), .B(new_n579_), .C1(new_n561_), .C2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT40), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(G1325gat));
  OAI21_X1  g382(.A(G15gat), .B1(new_n552_), .B2(new_n387_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT41), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT41), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n586_), .B(G15gat), .C1(new_n552_), .C2(new_n387_), .ZN(new_n587_));
  OR3_X1    g386(.A1(new_n561_), .A2(G15gat), .A3(new_n387_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n585_), .A2(new_n587_), .A3(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT99), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n585_), .A2(KEYINPUT99), .A3(new_n587_), .A4(new_n588_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(G1326gat));
  OAI21_X1  g392(.A(G22gat), .B1(new_n552_), .B2(new_n372_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT42), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n372_), .A2(G22gat), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n595_), .B1(new_n561_), .B2(new_n596_), .ZN(G1327gat));
  XNOR2_X1  g396(.A(new_n555_), .B(KEYINPUT37), .ZN(new_n598_));
  OAI21_X1  g397(.A(KEYINPUT43), .B1(new_n395_), .B2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT43), .ZN(new_n600_));
  INV_X1    g399(.A(new_n387_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n374_), .A2(new_n371_), .A3(new_n328_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n602_), .A2(new_n202_), .B1(new_n372_), .B2(new_n370_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n601_), .B1(new_n603_), .B2(new_n375_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n393_), .A2(new_n394_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n600_), .B(new_n557_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n599_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n607_), .A2(new_n531_), .A3(new_n559_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT44), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT100), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n548_), .B(KEYINPUT75), .ZN(new_n612_));
  AOI211_X1 g411(.A(new_n532_), .B(new_n612_), .C1(new_n599_), .C2(new_n606_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n611_), .B1(new_n613_), .B2(KEYINPUT44), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n608_), .A2(KEYINPUT100), .A3(new_n609_), .ZN(new_n615_));
  AOI211_X1 g414(.A(new_n328_), .B(new_n610_), .C1(new_n614_), .C2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(G29gat), .ZN(new_n617_));
  INV_X1    g416(.A(new_n455_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n612_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n554_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT101), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n554_), .A2(KEYINPUT101), .A3(new_n619_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n327_), .A2(new_n617_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT102), .ZN(new_n626_));
  OAI22_X1  g425(.A1(new_n616_), .A2(new_n617_), .B1(new_n624_), .B2(new_n626_), .ZN(G1328gat));
  INV_X1    g426(.A(KEYINPUT46), .ZN(new_n628_));
  INV_X1    g427(.A(G36gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n610_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(new_n572_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n622_), .A2(new_n629_), .A3(new_n572_), .A4(new_n623_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT45), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n628_), .B1(new_n631_), .B2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n610_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n615_), .ZN(new_n637_));
  AOI21_X1  g436(.A(KEYINPUT100), .B1(new_n608_), .B2(new_n609_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n572_), .B(new_n636_), .C1(new_n637_), .C2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(G36gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(new_n633_), .A3(KEYINPUT46), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n635_), .A2(new_n641_), .ZN(G1329gat));
  NAND2_X1  g441(.A1(new_n614_), .A2(new_n615_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n643_), .A2(G43gat), .A3(new_n601_), .A4(new_n636_), .ZN(new_n644_));
  INV_X1    g443(.A(G43gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n624_), .B2(new_n387_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT47), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT47), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n644_), .A2(new_n649_), .A3(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(G1330gat));
  INV_X1    g450(.A(G50gat), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n610_), .A2(new_n652_), .A3(new_n372_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n622_), .A2(new_n371_), .A3(new_n623_), .ZN(new_n654_));
  AOI22_X1  g453(.A1(new_n653_), .A2(new_n643_), .B1(new_n652_), .B2(new_n654_), .ZN(G1331gat));
  INV_X1    g454(.A(new_n500_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(new_n529_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n456_), .A2(new_n612_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT103), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n456_), .A2(KEYINPUT103), .A3(new_n612_), .A4(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(G57gat), .B1(new_n662_), .B2(new_n328_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n598_), .A2(new_n612_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n657_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n395_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n666_), .A2(new_n462_), .A3(new_n327_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n663_), .A2(new_n667_), .ZN(G1332gat));
  NAND3_X1  g467(.A1(new_n666_), .A2(new_n464_), .A3(new_n572_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n660_), .A2(new_n572_), .A3(new_n661_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT48), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(G64gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n670_), .B2(G64gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(G1333gat));
  INV_X1    g475(.A(G71gat), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n666_), .A2(new_n677_), .A3(new_n601_), .ZN(new_n678_));
  OAI21_X1  g477(.A(G71gat), .B1(new_n662_), .B2(new_n387_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n679_), .A2(KEYINPUT49), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(KEYINPUT49), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n678_), .B1(new_n680_), .B2(new_n681_), .ZN(G1334gat));
  OAI21_X1  g481(.A(G78gat), .B1(new_n662_), .B2(new_n372_), .ZN(new_n683_));
  XOR2_X1   g482(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n684_));
  OR2_X1    g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n684_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n372_), .A2(G78gat), .ZN(new_n687_));
  XOR2_X1   g486(.A(new_n687_), .B(KEYINPUT106), .Z(new_n688_));
  NAND2_X1  g487(.A1(new_n666_), .A2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n685_), .A2(new_n686_), .A3(new_n689_), .ZN(G1335gat));
  AOI211_X1 g489(.A(new_n612_), .B(new_n665_), .C1(new_n599_), .C2(new_n606_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G85gat), .B1(new_n692_), .B2(new_n328_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n619_), .B(new_n657_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT107), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n695_), .A2(new_n402_), .A3(new_n327_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n696_), .ZN(G1336gat));
  OAI21_X1  g496(.A(G92gat), .B1(new_n692_), .B2(new_n571_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n695_), .A2(new_n403_), .A3(new_n572_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1337gat));
  OAI21_X1  g499(.A(G99gat), .B1(new_n692_), .B2(new_n387_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n695_), .A2(new_n411_), .A3(new_n601_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n704_));
  XOR2_X1   g503(.A(new_n703_), .B(new_n704_), .Z(G1338gat));
  INV_X1    g504(.A(KEYINPUT52), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n607_), .A2(new_n371_), .A3(new_n559_), .A4(new_n657_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(G106gat), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n708_), .B1(new_n707_), .B2(G106gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n706_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n711_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(KEYINPUT52), .A3(new_n709_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n695_), .A2(new_n412_), .A3(new_n371_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n712_), .A2(new_n714_), .A3(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT53), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT53), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n712_), .A2(new_n714_), .A3(new_n715_), .A4(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1339gat));
  INV_X1    g519(.A(KEYINPUT117), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT54), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n500_), .A2(new_n529_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n560_), .B2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n723_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n664_), .A2(KEYINPUT54), .A3(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n724_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT113), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n515_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n520_), .A2(new_n515_), .A3(new_n508_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n525_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n728_), .B1(new_n729_), .B2(new_n731_), .ZN(new_n732_));
  OR3_X1    g531(.A1(new_n729_), .A2(new_n731_), .A3(new_n728_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n494_), .A2(new_n528_), .A3(new_n732_), .A4(new_n733_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n438_), .A2(KEYINPUT12), .A3(new_n476_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT12), .B1(new_n438_), .B2(new_n476_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n438_), .A2(new_n476_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n735_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n738_), .A2(KEYINPUT111), .A3(KEYINPUT55), .A4(new_n482_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT55), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n740_), .B1(new_n484_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n742_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n736_), .A2(new_n737_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n482_), .B1(new_n744_), .B2(new_n483_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n484_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n743_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(new_n491_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT56), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT56), .ZN(new_n752_));
  AOI211_X1 g551(.A(new_n752_), .B(new_n491_), .C1(new_n743_), .C2(new_n748_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n751_), .A2(new_n753_), .A3(KEYINPUT112), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n746_), .B1(new_n738_), .B2(new_n482_), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n742_), .A2(new_n739_), .B1(new_n755_), .B2(new_n484_), .ZN(new_n756_));
  OAI211_X1 g555(.A(KEYINPUT112), .B(new_n752_), .C1(new_n756_), .C2(new_n491_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n757_), .A2(new_n529_), .A3(new_n489_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n734_), .B1(new_n754_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n618_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT57), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT57), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(new_n762_), .A3(new_n618_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT58), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n752_), .B1(new_n756_), .B2(new_n491_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n749_), .A2(KEYINPUT56), .A3(new_n750_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n528_), .A2(new_n489_), .A3(new_n733_), .A4(new_n732_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n766_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT114), .B(new_n770_), .C1(new_n767_), .C2(new_n768_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n765_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n557_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n770_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT58), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT116), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n775_), .B1(new_n774_), .B2(new_n557_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n764_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n727_), .B1(new_n782_), .B2(new_n549_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n393_), .A2(new_n327_), .A3(new_n601_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n721_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n784_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n771_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT114), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n777_), .A2(new_n766_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT58), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT115), .B1(new_n790_), .B2(new_n598_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(new_n776_), .A3(new_n779_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n548_), .B1(new_n792_), .B2(new_n764_), .ZN(new_n793_));
  OAI211_X1 g592(.A(KEYINPUT117), .B(new_n786_), .C1(new_n793_), .C2(new_n727_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n785_), .A2(new_n529_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(G113gat), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n795_), .A2(KEYINPUT118), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT118), .B1(new_n795_), .B2(new_n796_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n782_), .A2(new_n559_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n727_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  XOR2_X1   g600(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n786_), .A3(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(KEYINPUT59), .B1(new_n783_), .B2(new_n784_), .ZN(new_n804_));
  AND4_X1   g603(.A1(G113gat), .A2(new_n803_), .A3(new_n529_), .A4(new_n804_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n797_), .A2(new_n798_), .A3(new_n805_), .ZN(G1340gat));
  INV_X1    g605(.A(KEYINPUT60), .ZN(new_n807_));
  XOR2_X1   g606(.A(KEYINPUT120), .B(G120gat), .Z(new_n808_));
  NAND3_X1  g607(.A1(new_n500_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n785_), .A2(new_n794_), .A3(new_n810_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n803_), .A2(new_n500_), .A3(new_n804_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n811_), .B1(new_n812_), .B2(new_n808_), .ZN(G1341gat));
  NAND3_X1  g612(.A1(new_n803_), .A2(new_n548_), .A3(new_n804_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(G127gat), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n559_), .A2(G127gat), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n785_), .A2(new_n794_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1342gat));
  NAND3_X1  g617(.A1(new_n803_), .A2(new_n557_), .A3(new_n804_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(G134gat), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n618_), .A2(G134gat), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n785_), .A2(new_n794_), .A3(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(G1343gat));
  NAND3_X1  g622(.A1(new_n387_), .A2(new_n327_), .A3(new_n371_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n783_), .A2(new_n572_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n529_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n500_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g628(.A1(new_n825_), .A2(new_n612_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(KEYINPUT61), .B(G155gat), .ZN(new_n831_));
  XNOR2_X1  g630(.A(new_n830_), .B(new_n831_), .ZN(G1346gat));
  NAND3_X1  g631(.A1(new_n825_), .A2(new_n297_), .A3(new_n455_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n825_), .A2(new_n557_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n833_), .B1(new_n835_), .B2(new_n297_), .ZN(G1347gat));
  NAND2_X1  g635(.A1(new_n572_), .A2(new_n394_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n371_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n801_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n226_), .A3(new_n529_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT62), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT121), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n801_), .A2(new_n842_), .A3(new_n529_), .A4(new_n838_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n612_), .B1(new_n792_), .B2(new_n764_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n529_), .B(new_n838_), .C1(new_n844_), .C2(new_n727_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT121), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n843_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n841_), .B1(new_n847_), .B2(G169gat), .ZN(new_n848_));
  AOI211_X1 g647(.A(KEYINPUT62), .B(new_n215_), .C1(new_n843_), .C2(new_n846_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n840_), .B1(new_n848_), .B2(new_n849_), .ZN(G1348gat));
  AOI21_X1  g649(.A(G176gat), .B1(new_n839_), .B2(new_n500_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n783_), .A2(new_n371_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n837_), .A2(new_n216_), .A3(new_n656_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n852_), .B2(new_n853_), .ZN(G1349gat));
  NAND4_X1  g653(.A1(new_n852_), .A2(new_n572_), .A3(new_n394_), .A4(new_n612_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n549_), .A2(new_n246_), .ZN(new_n856_));
  AOI22_X1  g655(.A1(new_n855_), .A2(new_n204_), .B1(new_n839_), .B2(new_n856_), .ZN(G1350gat));
  NAND2_X1  g656(.A1(new_n455_), .A2(new_n203_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT122), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n839_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n839_), .A2(new_n557_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n860_), .B1(new_n862_), .B2(new_n210_), .ZN(G1351gat));
  INV_X1    g662(.A(new_n783_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n387_), .A2(new_n328_), .A3(new_n371_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n572_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n867_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n864_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(G197gat), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n869_), .A2(KEYINPUT124), .A3(new_n870_), .A4(new_n530_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n870_), .B1(new_n869_), .B2(new_n530_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n869_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n875_), .A2(G197gat), .A3(new_n529_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n871_), .B1(new_n874_), .B2(new_n876_), .ZN(G1352gat));
  AOI21_X1  g676(.A(new_n656_), .B1(KEYINPUT125), .B2(G204gat), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n878_), .ZN(new_n879_));
  OR2_X1    g678(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1353gat));
  AOI21_X1  g680(.A(new_n549_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n864_), .A2(new_n868_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT126), .ZN(new_n884_));
  NOR2_X1   g683(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n885_));
  OR3_X1    g684(.A1(new_n883_), .A2(new_n884_), .A3(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n884_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n885_), .ZN(new_n888_));
  AND3_X1   g687(.A1(new_n886_), .A2(new_n887_), .A3(new_n888_), .ZN(G1354gat));
  NAND2_X1  g688(.A1(new_n875_), .A2(new_n455_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT127), .B(G218gat), .Z(new_n891_));
  NOR2_X1   g690(.A1(new_n598_), .A2(new_n891_), .ZN(new_n892_));
  AOI22_X1  g691(.A1(new_n890_), .A2(new_n891_), .B1(new_n875_), .B2(new_n892_), .ZN(G1355gat));
endmodule


