//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n912_, new_n914_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n967_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_;
  XNOR2_X1  g000(.A(G113gat), .B(G120gat), .ZN(new_n202_));
  INV_X1    g001(.A(G134gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G127gat), .ZN(new_n204_));
  INV_X1    g003(.A(G127gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G134gat), .ZN(new_n206_));
  AND3_X1   g005(.A1(new_n204_), .A2(new_n206_), .A3(KEYINPUT86), .ZN(new_n207_));
  AOI21_X1  g006(.A(KEYINPUT86), .B1(new_n204_), .B2(new_n206_), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n202_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT87), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT86), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n205_), .A2(G134gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n203_), .A2(G127gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n211_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n204_), .A2(new_n206_), .A3(KEYINPUT86), .ZN(new_n215_));
  XOR2_X1   g014(.A(G113gat), .B(G120gat), .Z(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  AND3_X1   g016(.A1(new_n209_), .A2(new_n210_), .A3(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n210_), .B1(new_n209_), .B2(new_n217_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT22), .B(G169gat), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT83), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n223_), .A2(KEYINPUT83), .A3(new_n224_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(G183gat), .A3(G190gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT81), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT81), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n235_), .A2(G183gat), .A3(G190gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n232_), .B1(new_n237_), .B2(new_n231_), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n227_), .A2(new_n228_), .B1(new_n230_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n233_), .A2(KEYINPUT23), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT80), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n233_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n231_), .A2(new_n237_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT79), .ZN(new_n245_));
  INV_X1    g044(.A(G169gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(new_n222_), .ZN(new_n247_));
  OAI21_X1  g046(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT24), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT82), .B1(new_n244_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n242_), .A2(new_n243_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n235_), .B1(G183gat), .B2(G190gat), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n233_), .A2(KEYINPUT81), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n231_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT82), .ZN(new_n256_));
  INV_X1    g055(.A(new_n249_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n250_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(G183gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT78), .B1(new_n260_), .B2(KEYINPUT25), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(G190gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT25), .B(G183gat), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n261_), .B(new_n262_), .C1(new_n263_), .C2(KEYINPUT78), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n247_), .A2(KEYINPUT24), .A3(new_n248_), .A4(new_n224_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n239_), .B1(new_n259_), .B2(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(KEYINPUT84), .B(KEYINPUT30), .Z(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n266_), .B1(new_n250_), .B2(new_n258_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n269_), .B1(new_n272_), .B2(new_n239_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(G15gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(G71gat), .B(G99gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT85), .B(G43gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n271_), .A2(new_n273_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n279_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n282_));
  NOR3_X1   g081(.A1(new_n281_), .A2(new_n282_), .A3(KEYINPUT31), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT31), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n271_), .A2(new_n273_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n279_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n284_), .B1(new_n287_), .B2(new_n280_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n220_), .B1(new_n283_), .B2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT31), .B1(new_n281_), .B2(new_n282_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(new_n284_), .A3(new_n280_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n220_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n289_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT27), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G226gat), .A2(G233gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT19), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT92), .ZN(new_n300_));
  OR2_X1    g099(.A1(new_n263_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n263_), .A2(new_n300_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n302_), .A3(new_n262_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT24), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(new_n246_), .A3(new_n222_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n303_), .A2(new_n265_), .A3(new_n238_), .A4(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G211gat), .B(G218gat), .ZN(new_n307_));
  INV_X1    g106(.A(G197gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT91), .B1(new_n308_), .B2(G204gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(KEYINPUT21), .A3(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G197gat), .B(G204gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n313_), .A2(KEYINPUT21), .A3(new_n307_), .A4(new_n309_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n307_), .A2(KEYINPUT21), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n312_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n224_), .B(new_n223_), .C1(new_n244_), .C2(new_n229_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n306_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT20), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT93), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n256_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n322_));
  AOI211_X1 g121(.A(KEYINPUT82), .B(new_n249_), .C1(new_n251_), .C2(new_n254_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n267_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n239_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n316_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n321_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n321_), .B(new_n327_), .C1(new_n272_), .C2(new_n239_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n299_), .B(new_n320_), .C1(new_n328_), .C2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G8gat), .B(G36gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT18), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G64gat), .B(G92gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  NAND2_X1  g134(.A1(new_n268_), .A2(new_n316_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n306_), .A2(new_n317_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT20), .B1(new_n338_), .B2(new_n316_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n298_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n331_), .A2(new_n335_), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n335_), .B1(new_n331_), .B2(new_n340_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n296_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT98), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI211_X1 g144(.A(KEYINPUT98), .B(new_n296_), .C1(new_n341_), .C2(new_n342_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n298_), .B(new_n320_), .C1(new_n328_), .C2(new_n330_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n335_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n299_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT97), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n331_), .A2(new_n335_), .A3(new_n340_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT97), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n347_), .A2(new_n349_), .A3(new_n353_), .A4(new_n348_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n351_), .A2(KEYINPUT27), .A3(new_n352_), .A4(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT94), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n207_), .A2(new_n208_), .A3(new_n202_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n216_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT87), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n209_), .A2(new_n217_), .A3(new_n210_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT88), .ZN(new_n361_));
  NOR2_X1   g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G155gat), .A2(G162gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(G141gat), .ZN(new_n366_));
  INV_X1    g165(.A(G148gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT2), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT2), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n369_), .A2(G141gat), .A3(G148gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n366_), .A2(new_n367_), .A3(KEYINPUT3), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(G141gat), .B2(G148gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n365_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G141gat), .B(G148gat), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n362_), .B1(KEYINPUT1), .B2(new_n364_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT1), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(G155gat), .A3(G162gat), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n377_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n361_), .B1(new_n376_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n377_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n364_), .A2(KEYINPUT1), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n363_), .A2(new_n384_), .A3(new_n380_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n368_), .A2(new_n370_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n386_), .B(KEYINPUT88), .C1(new_n387_), .C2(new_n365_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n359_), .A2(new_n360_), .A3(new_n382_), .A4(new_n388_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n356_), .B1(new_n389_), .B2(KEYINPUT4), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n382_), .A2(new_n388_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n220_), .A2(new_n391_), .A3(KEYINPUT94), .A4(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G225gat), .A2(G233gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n376_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n397_), .A2(new_n217_), .A3(new_n209_), .A4(new_n386_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n389_), .A2(new_n398_), .A3(KEYINPUT4), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n394_), .A2(new_n396_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n389_), .A2(new_n398_), .A3(new_n395_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT96), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n389_), .A2(new_n398_), .A3(KEYINPUT96), .A4(new_n395_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n400_), .A2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G1gat), .B(G29gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT0), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(G57gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT95), .B(G85gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n406_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n400_), .A2(new_n405_), .A3(new_n411_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G22gat), .B(G50gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT90), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n382_), .A2(new_n388_), .A3(KEYINPUT29), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G228gat), .A2(G233gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n316_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n417_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT29), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(new_n397_), .B2(new_n386_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n419_), .B1(new_n423_), .B2(new_n316_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G78gat), .B(G106gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n421_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n416_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n421_), .A2(new_n424_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n425_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n421_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n416_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  XOR2_X1   g233(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n391_), .A2(KEYINPUT29), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n382_), .A2(new_n388_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n435_), .B1(new_n438_), .B2(new_n422_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n429_), .A2(new_n434_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n440_), .B1(new_n429_), .B2(new_n434_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n413_), .B(new_n414_), .C1(new_n441_), .C2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n345_), .A2(new_n346_), .A3(new_n355_), .A4(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n347_), .A2(new_n349_), .A3(KEYINPUT32), .A4(new_n335_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n335_), .A2(KEYINPUT32), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n331_), .A2(new_n340_), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n414_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n411_), .B1(new_n400_), .B2(new_n405_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n446_), .B(new_n448_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT33), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n414_), .A2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n400_), .A2(KEYINPUT33), .A3(new_n405_), .A4(new_n411_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n394_), .A2(new_n395_), .A3(new_n399_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n389_), .A2(new_n398_), .A3(new_n396_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(new_n412_), .A3(new_n456_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n453_), .A2(new_n454_), .A3(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT93), .B1(new_n268_), .B2(new_n316_), .ZN(new_n459_));
  AOI211_X1 g258(.A(new_n298_), .B(new_n319_), .C1(new_n459_), .C2(new_n329_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n339_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n299_), .B1(new_n461_), .B2(new_n336_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n348_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n352_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n451_), .B1(new_n458_), .B2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n441_), .A2(new_n442_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n295_), .B1(new_n445_), .B2(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n449_), .A2(new_n450_), .ZN(new_n469_));
  AND4_X1   g268(.A1(new_n469_), .A2(new_n289_), .A3(new_n466_), .A4(new_n293_), .ZN(new_n470_));
  AND4_X1   g269(.A1(new_n346_), .A2(new_n470_), .A3(new_n355_), .A4(new_n345_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT12), .ZN(new_n473_));
  XNOR2_X1  g272(.A(KEYINPUT10), .B(G99gat), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT64), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(KEYINPUT64), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(G106gat), .B1(new_n476_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G99gat), .A2(G106gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT6), .ZN(new_n482_));
  INV_X1    g281(.A(G85gat), .ZN(new_n483_));
  INV_X1    g282(.A(G92gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G85gat), .A2(G92gat), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(KEYINPUT9), .A3(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n486_), .A2(KEYINPUT9), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n482_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n480_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n481_), .B(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT7), .ZN(new_n493_));
  INV_X1    g292(.A(G99gat), .ZN(new_n494_));
  INV_X1    g293(.A(G106gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n493_), .A2(new_n494_), .A3(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT66), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT66), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n496_), .A2(new_n500_), .A3(new_n497_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n492_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n485_), .A2(new_n486_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT65), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT8), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT65), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n503_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT8), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n507_), .B(new_n508_), .C1(new_n492_), .C2(new_n498_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n490_), .B1(new_n505_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G57gat), .B(G64gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G71gat), .B(G78gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(KEYINPUT11), .ZN(new_n513_));
  XOR2_X1   g312(.A(G71gat), .B(G78gat), .Z(new_n514_));
  INV_X1    g313(.A(G64gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(G57gat), .ZN(new_n516_));
  INV_X1    g315(.A(G57gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(G64gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n518_), .A3(KEYINPUT11), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n514_), .A2(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n511_), .A2(KEYINPUT11), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n513_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n473_), .B1(new_n510_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n501_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n500_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n482_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n508_), .B1(new_n526_), .B2(new_n507_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n492_), .A2(new_n498_), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n504_), .A2(new_n528_), .A3(KEYINPUT8), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n482_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n479_), .ZN(new_n531_));
  AOI21_X1  g330(.A(KEYINPUT64), .B1(new_n477_), .B2(new_n478_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n495_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(KEYINPUT67), .B1(new_n530_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT67), .ZN(new_n535_));
  NOR3_X1   g334(.A1(new_n480_), .A2(new_n489_), .A3(new_n535_), .ZN(new_n536_));
  OAI22_X1  g335(.A1(new_n527_), .A2(new_n529_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n522_), .A2(KEYINPUT68), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT68), .ZN(new_n539_));
  OAI211_X1 g338(.A(new_n539_), .B(new_n513_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(new_n473_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n537_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(G230gat), .ZN(new_n544_));
  INV_X1    g343(.A(G233gat), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n510_), .A2(new_n522_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n523_), .A2(new_n543_), .A3(new_n547_), .A4(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n510_), .A2(new_n522_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n522_), .ZN(new_n551_));
  AOI211_X1 g350(.A(new_n490_), .B(new_n551_), .C1(new_n505_), .C2(new_n509_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n546_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G120gat), .B(G148gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT5), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G176gat), .B(G204gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n555_), .B(new_n556_), .Z(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n549_), .A2(new_n553_), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT69), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n549_), .A2(new_n553_), .A3(KEYINPUT69), .A4(new_n558_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n549_), .A2(new_n553_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(new_n557_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT13), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n563_), .A2(KEYINPUT13), .A3(new_n565_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT70), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G229gat), .A2(G233gat), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G29gat), .B(G36gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G43gat), .B(G50gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G15gat), .B(G22gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(KEYINPUT72), .B(G1gat), .ZN(new_n578_));
  INV_X1    g377(.A(G8gat), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT14), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n577_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT73), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT73), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n584_), .B(new_n577_), .C1(new_n580_), .C2(new_n581_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G1gat), .B(G8gat), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n583_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n587_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n576_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n590_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n576_), .B(KEYINPUT15), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n592_), .A2(new_n588_), .A3(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n573_), .B1(new_n591_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n576_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n592_), .A2(new_n588_), .A3(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n591_), .A2(new_n598_), .A3(new_n573_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G113gat), .B(G141gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(G169gat), .B(G197gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n596_), .A2(new_n599_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n602_), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n591_), .A2(new_n598_), .A3(new_n573_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n604_), .B1(new_n605_), .B2(new_n595_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n589_), .A2(new_n590_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT74), .Z(new_n611_));
  OR2_X1    g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n609_), .A2(new_n611_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n522_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G127gat), .B(G155gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT16), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT17), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n612_), .A2(new_n613_), .A3(new_n551_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n619_), .A2(KEYINPUT17), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n615_), .A2(new_n620_), .A3(new_n621_), .A4(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n541_), .B(KEYINPUT75), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n614_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n614_), .A2(new_n624_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n620_), .B(KEYINPUT76), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n623_), .B1(new_n625_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT77), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT37), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT35), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n634_));
  NAND2_X1  g433(.A1(G232gat), .A2(G233gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI22_X1  g436(.A1(new_n510_), .A2(new_n576_), .B1(new_n633_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n537_), .A2(new_n593_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n637_), .A2(new_n633_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(G190gat), .B(G218gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(G134gat), .B(G162gat), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n645_), .A2(KEYINPUT36), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n640_), .A2(new_n641_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n642_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n645_), .B(KEYINPUT36), .Z(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n642_), .B2(new_n647_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n632_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n652_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(KEYINPUT37), .A3(new_n648_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n631_), .A2(new_n657_), .ZN(new_n658_));
  NOR4_X1   g457(.A1(new_n472_), .A2(new_n571_), .A3(new_n608_), .A4(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n469_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n660_), .A3(new_n578_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT38), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n445_), .A2(new_n467_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n294_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n345_), .A2(new_n355_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n346_), .A3(new_n470_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n570_), .A2(new_n608_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(KEYINPUT99), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT99), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n670_), .B1(new_n570_), .B2(new_n608_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n629_), .B(KEYINPUT77), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n649_), .A2(new_n652_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n667_), .A2(new_n672_), .A3(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G1gat), .B1(new_n676_), .B2(new_n469_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n662_), .A2(new_n677_), .ZN(G1324gat));
  NAND2_X1  g477(.A1(new_n665_), .A2(new_n346_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n659_), .A2(new_n579_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n679_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G8gat), .B1(new_n676_), .B2(new_n681_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(KEYINPUT39), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT101), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(KEYINPUT39), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT100), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n680_), .B1(new_n684_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT40), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n687_), .B(new_n688_), .ZN(G1325gat));
  OAI21_X1  g488(.A(G15gat), .B1(new_n676_), .B2(new_n294_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n690_), .A2(KEYINPUT41), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(KEYINPUT41), .ZN(new_n692_));
  INV_X1    g491(.A(G15gat), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n659_), .A2(new_n693_), .A3(new_n295_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n691_), .A2(new_n692_), .A3(new_n694_), .ZN(G1326gat));
  OAI21_X1  g494(.A(G22gat), .B1(new_n676_), .B2(new_n466_), .ZN(new_n696_));
  XOR2_X1   g495(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n697_));
  OR2_X1    g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n697_), .ZN(new_n699_));
  INV_X1    g498(.A(G22gat), .ZN(new_n700_));
  INV_X1    g499(.A(new_n466_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n659_), .A2(new_n700_), .A3(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n698_), .A2(new_n699_), .A3(new_n702_), .ZN(G1327gat));
  OAI211_X1 g502(.A(KEYINPUT43), .B(new_n656_), .C1(new_n468_), .C2(new_n471_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n631_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n657_), .B1(new_n664_), .B2(new_n666_), .ZN(new_n706_));
  XOR2_X1   g505(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n707_));
  OAI211_X1 g506(.A(new_n704_), .B(new_n705_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n707_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n711_), .B1(new_n472_), .B2(new_n657_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n712_), .A2(KEYINPUT104), .A3(new_n704_), .A4(new_n705_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT44), .B1(new_n710_), .B2(new_n713_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n712_), .A2(KEYINPUT44), .A3(new_n704_), .A4(new_n705_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n660_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G29gat), .B1(new_n714_), .B2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT105), .ZN(new_n718_));
  INV_X1    g517(.A(new_n674_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n631_), .A2(new_n719_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n667_), .A2(new_n668_), .A3(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(G29gat), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n660_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n718_), .A2(new_n723_), .ZN(G1328gat));
  NAND2_X1  g523(.A1(new_n710_), .A2(new_n713_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n715_), .A2(new_n679_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n727_), .A2(new_n728_), .A3(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT106), .B1(new_n714_), .B2(new_n729_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(G36gat), .A3(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(G36gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n721_), .A2(new_n734_), .A3(new_n679_), .ZN(new_n735_));
  XOR2_X1   g534(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n736_));
  XNOR2_X1  g535(.A(new_n735_), .B(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n733_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n733_), .A2(KEYINPUT46), .A3(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1329gat));
  NAND3_X1  g541(.A1(new_n715_), .A2(G43gat), .A3(new_n295_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n721_), .A2(new_n295_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  OAI22_X1  g544(.A1(new_n714_), .A2(new_n743_), .B1(G43gat), .B2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g546(.A(G50gat), .B1(new_n721_), .B2(new_n701_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n715_), .A2(G50gat), .A3(new_n701_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n727_), .B2(new_n749_), .ZN(G1331gat));
  INV_X1    g549(.A(new_n570_), .ZN(new_n751_));
  NOR2_X1   g550(.A1(new_n658_), .A2(new_n751_), .ZN(new_n752_));
  XNOR2_X1  g551(.A(new_n752_), .B(KEYINPUT108), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n472_), .A2(new_n607_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n517_), .A3(new_n660_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n571_), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n757_), .A2(new_n673_), .A3(new_n674_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n758_), .A2(new_n660_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n756_), .B1(new_n759_), .B2(new_n517_), .ZN(G1332gat));
  AOI21_X1  g559(.A(new_n515_), .B1(new_n758_), .B2(new_n679_), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT48), .Z(new_n762_));
  NAND3_X1  g561(.A1(new_n755_), .A2(new_n515_), .A3(new_n679_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(G1333gat));
  INV_X1    g563(.A(G71gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n765_), .B1(new_n758_), .B2(new_n295_), .ZN(new_n766_));
  XOR2_X1   g565(.A(new_n766_), .B(KEYINPUT49), .Z(new_n767_));
  NAND3_X1  g566(.A1(new_n755_), .A2(new_n765_), .A3(new_n295_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1334gat));
  INV_X1    g568(.A(G78gat), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n755_), .A2(new_n770_), .A3(new_n701_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n758_), .B2(new_n701_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n772_), .A2(new_n773_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n771_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT109), .B(new_n771_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1335gat));
  NAND3_X1  g579(.A1(new_n754_), .A2(new_n571_), .A3(new_n720_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n781_), .A2(G85gat), .A3(new_n469_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n712_), .A2(new_n704_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n631_), .A2(new_n751_), .A3(new_n607_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n660_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n782_), .B1(new_n786_), .B2(G85gat), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n787_), .B(KEYINPUT110), .ZN(G1336gat));
  NAND3_X1  g587(.A1(new_n785_), .A2(G92gat), .A3(new_n679_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n484_), .B1(new_n781_), .B2(new_n681_), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n790_), .A2(KEYINPUT111), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(KEYINPUT111), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n789_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  XOR2_X1   g592(.A(new_n793_), .B(KEYINPUT112), .Z(G1337gat));
  NAND2_X1  g593(.A1(new_n785_), .A2(new_n295_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(G99gat), .ZN(new_n796_));
  INV_X1    g595(.A(new_n781_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n797_), .B(new_n295_), .C1(new_n531_), .C2(new_n532_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799_));
  AOI22_X1  g598(.A1(new_n796_), .A2(new_n798_), .B1(KEYINPUT113), .B2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(KEYINPUT113), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(G1338gat));
  NAND3_X1  g601(.A1(new_n783_), .A2(new_n701_), .A3(new_n784_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n804_), .A3(G106gat), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT114), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT114), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n803_), .A2(new_n807_), .A3(new_n804_), .A4(G106gat), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n803_), .A2(G106gat), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT52), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n806_), .A2(new_n808_), .A3(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n797_), .A2(new_n495_), .A3(new_n701_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(G1339gat));
  NAND3_X1  g615(.A1(new_n591_), .A2(new_n594_), .A3(new_n573_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n591_), .A2(new_n598_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n602_), .B(new_n817_), .C1(new_n818_), .C2(new_n573_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n606_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n523_), .A2(new_n543_), .A3(KEYINPUT55), .A4(new_n548_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n546_), .A2(KEYINPUT116), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n549_), .A2(new_n826_), .ZN(new_n827_));
  AOI22_X1  g626(.A1(new_n537_), .A2(new_n542_), .B1(new_n510_), .B2(new_n522_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n828_), .A2(KEYINPUT55), .A3(new_n523_), .A4(new_n823_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n825_), .A2(new_n827_), .A3(new_n829_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n557_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT56), .B1(new_n830_), .B2(new_n557_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n821_), .B(KEYINPUT58), .C1(new_n831_), .C2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n656_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n830_), .A2(new_n557_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n557_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(KEYINPUT58), .B1(new_n839_), .B2(new_n821_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n834_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n563_), .A2(new_n607_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n843_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n820_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT57), .B(new_n719_), .C1(new_n844_), .C2(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n846_), .A2(KEYINPUT118), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n561_), .A2(new_n562_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n845_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n674_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n848_), .B1(new_n852_), .B2(KEYINPUT57), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n842_), .B1(new_n847_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n719_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT117), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT117), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n852_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(KEYINPUT57), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n673_), .B1(new_n854_), .B2(new_n859_), .ZN(new_n860_));
  NOR3_X1   g659(.A1(new_n673_), .A2(new_n607_), .A3(new_n656_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(KEYINPUT54), .A3(new_n751_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT54), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n631_), .A2(new_n608_), .A3(new_n657_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n570_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n860_), .A2(new_n867_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n294_), .A2(new_n701_), .A3(new_n469_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n681_), .A3(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT59), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n679_), .B1(new_n860_), .B2(new_n867_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n873_), .A2(KEYINPUT59), .A3(new_n869_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n872_), .A2(new_n874_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G113gat), .B1(new_n875_), .B2(new_n608_), .ZN(new_n876_));
  OR3_X1    g675(.A1(new_n870_), .A2(G113gat), .A3(new_n608_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1340gat));
  INV_X1    g677(.A(new_n571_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G120gat), .B1(new_n875_), .B2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n870_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT60), .ZN(new_n882_));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n570_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n884_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n881_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n880_), .A2(new_n886_), .ZN(G1341gat));
  OAI21_X1  g686(.A(G127gat), .B1(new_n875_), .B2(new_n673_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n881_), .A2(new_n205_), .A3(new_n631_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1342gat));
  NAND3_X1  g689(.A1(new_n881_), .A2(new_n203_), .A3(new_n674_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n657_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(new_n892_), .B2(new_n203_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(KEYINPUT119), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n895_), .B(new_n891_), .C1(new_n892_), .C2(new_n203_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1343gat));
  NOR3_X1   g696(.A1(new_n295_), .A2(new_n469_), .A3(new_n466_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n846_), .A2(KEYINPUT118), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n852_), .A2(new_n848_), .A3(KEYINPUT57), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n841_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n852_), .A2(new_n857_), .ZN(new_n903_));
  AOI211_X1 g702(.A(KEYINPUT117), .B(new_n674_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n902_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n631_), .B1(new_n901_), .B2(new_n905_), .ZN(new_n906_));
  OAI211_X1 g705(.A(new_n681_), .B(new_n898_), .C1(new_n906_), .C2(new_n866_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(KEYINPUT120), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n868_), .A2(new_n909_), .A3(new_n681_), .A4(new_n898_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n908_), .A2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n607_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n571_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g714(.A(KEYINPUT61), .B(G155gat), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT121), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n917_), .B1(new_n911_), .B2(new_n631_), .ZN(new_n918_));
  AOI211_X1 g717(.A(KEYINPUT121), .B(new_n673_), .C1(new_n908_), .C2(new_n910_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n916_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n909_), .B1(new_n873_), .B2(new_n898_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n907_), .A2(KEYINPUT120), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n631_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(KEYINPUT121), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n911_), .A2(new_n917_), .A3(new_n631_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n916_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n924_), .A2(new_n925_), .A3(new_n926_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n920_), .A2(new_n927_), .ZN(G1346gat));
  INV_X1    g727(.A(new_n911_), .ZN(new_n929_));
  OR3_X1    g728(.A1(new_n929_), .A2(G162gat), .A3(new_n719_), .ZN(new_n930_));
  OAI21_X1  g729(.A(G162gat), .B1(new_n929_), .B2(new_n657_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1347gat));
  AOI21_X1  g731(.A(new_n681_), .B1(new_n860_), .B2(new_n867_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n933_), .A2(new_n470_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n935_), .A2(new_n221_), .A3(new_n607_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n933_), .A2(new_n470_), .A3(new_n607_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n937_), .B1(new_n938_), .B2(G169gat), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT122), .ZN(new_n940_));
  AND2_X1   g739(.A1(new_n939_), .A2(new_n940_), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n938_), .A2(new_n937_), .A3(G169gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n942_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n936_), .B1(new_n941_), .B2(new_n943_), .ZN(G1348gat));
  OAI21_X1  g743(.A(G176gat), .B1(new_n934_), .B2(new_n879_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n570_), .A2(new_n222_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n934_), .B2(new_n946_), .ZN(G1349gat));
  AOI21_X1  g746(.A(new_n260_), .B1(new_n935_), .B2(new_n631_), .ZN(new_n948_));
  INV_X1    g747(.A(new_n948_), .ZN(new_n949_));
  INV_X1    g748(.A(KEYINPUT123), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n301_), .A2(new_n302_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n935_), .A2(new_n631_), .ZN(new_n952_));
  OAI211_X1 g751(.A(new_n949_), .B(new_n950_), .C1(new_n951_), .C2(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n952_), .A2(new_n951_), .ZN(new_n954_));
  OAI21_X1  g753(.A(KEYINPUT123), .B1(new_n954_), .B2(new_n948_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n953_), .A2(new_n955_), .ZN(G1350gat));
  OAI21_X1  g755(.A(G190gat), .B1(new_n934_), .B2(new_n657_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n674_), .A2(new_n262_), .ZN(new_n958_));
  XOR2_X1   g757(.A(new_n958_), .B(KEYINPUT124), .Z(new_n959_));
  OAI21_X1  g758(.A(new_n957_), .B1(new_n934_), .B2(new_n959_), .ZN(G1351gat));
  NOR2_X1   g759(.A1(new_n295_), .A2(new_n443_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n933_), .A2(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n962_), .A2(new_n608_), .ZN(new_n963_));
  XOR2_X1   g762(.A(KEYINPUT125), .B(G197gat), .Z(new_n964_));
  XNOR2_X1  g763(.A(new_n963_), .B(new_n964_), .ZN(G1352gat));
  INV_X1    g764(.A(new_n962_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n966_), .A2(new_n571_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g767(.A(new_n673_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n966_), .A2(new_n969_), .ZN(new_n970_));
  INV_X1    g769(.A(KEYINPUT127), .ZN(new_n971_));
  NOR2_X1   g770(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n972_));
  XOR2_X1   g771(.A(new_n972_), .B(KEYINPUT126), .Z(new_n973_));
  NAND3_X1  g772(.A1(new_n970_), .A2(new_n971_), .A3(new_n973_), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n974_), .B1(new_n970_), .B2(new_n973_), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n971_), .B1(new_n970_), .B2(new_n973_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n975_), .A2(new_n976_), .ZN(G1354gat));
  OAI21_X1  g776(.A(G218gat), .B1(new_n962_), .B2(new_n657_), .ZN(new_n978_));
  OR2_X1    g777(.A1(new_n719_), .A2(G218gat), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n978_), .B1(new_n962_), .B2(new_n979_), .ZN(G1355gat));
endmodule


