//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_, new_n889_, new_n890_, new_n891_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n928_, new_n929_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G43gat), .B(G50gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G29gat), .B(G36gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G43gat), .B(G50gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT15), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210_));
  INV_X1    g009(.A(G1gat), .ZN(new_n211_));
  INV_X1    g010(.A(G8gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G1gat), .B(G8gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n209_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n208_), .ZN(new_n218_));
  OR2_X1    g017(.A1(new_n216_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G229gat), .A2(G233gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n216_), .B(new_n218_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n220_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n221_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G113gat), .B(G141gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G169gat), .B(G197gat), .ZN(new_n227_));
  XOR2_X1   g026(.A(new_n226_), .B(new_n227_), .Z(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n225_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT78), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n221_), .A2(new_n224_), .A3(new_n228_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n225_), .A2(KEYINPUT78), .A3(new_n229_), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G141gat), .ZN(new_n237_));
  INV_X1    g036(.A(G148gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G141gat), .A2(G148gat), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G155gat), .A2(G162gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT83), .B1(new_n242_), .B2(KEYINPUT1), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT83), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT1), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n244_), .A2(new_n245_), .A3(G155gat), .A4(G162gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G155gat), .ZN(new_n248_));
  INV_X1    g047(.A(G162gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n249_), .A3(KEYINPUT82), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n242_), .A2(KEYINPUT1), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT82), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n252_), .B1(G155gat), .B2(G162gat), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n250_), .A2(new_n251_), .A3(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n241_), .B1(new_n247_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT84), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(KEYINPUT84), .B(new_n241_), .C1(new_n247_), .C2(new_n254_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT29), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n250_), .A2(new_n253_), .A3(new_n242_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT87), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT87), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n250_), .A2(new_n253_), .A3(new_n263_), .A4(new_n242_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT3), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(KEYINPUT85), .A3(new_n266_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT2), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n240_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n240_), .A2(new_n273_), .ZN(new_n276_));
  AOI22_X1  g075(.A1(KEYINPUT2), .A2(new_n276_), .B1(new_n239_), .B2(KEYINPUT3), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n272_), .A2(new_n275_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT88), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n265_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n279_), .B1(new_n265_), .B2(new_n278_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n259_), .B(new_n260_), .C1(new_n280_), .C2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT28), .ZN(new_n283_));
  AND2_X1   g082(.A1(new_n262_), .A2(new_n264_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n276_), .A2(KEYINPUT2), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n239_), .A2(KEYINPUT3), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(new_n275_), .A3(new_n286_), .ZN(new_n287_));
  NOR4_X1   g086(.A1(new_n268_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT85), .B1(new_n270_), .B2(new_n266_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT88), .B1(new_n284_), .B2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n265_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT28), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(new_n260_), .A4(new_n259_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n283_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G22gat), .B(G50gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n283_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G78gat), .B(G106gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT93), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G228gat), .A2(G233gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT21), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n308_), .B1(G197gat), .B2(G204gat), .ZN(new_n309_));
  INV_X1    g108(.A(G204gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT89), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT89), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(G204gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n309_), .B1(new_n314_), .B2(G197gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G211gat), .B(G218gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT90), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G197gat), .A2(G204gat), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(new_n314_), .B2(G197gat), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n318_), .B1(new_n320_), .B2(KEYINPUT21), .ZN(new_n321_));
  INV_X1    g120(.A(G197gat), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n322_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n323_));
  OAI211_X1 g122(.A(KEYINPUT90), .B(new_n308_), .C1(new_n323_), .C2(new_n319_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n317_), .B1(new_n321_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n319_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT89), .B(G204gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n326_), .B1(new_n327_), .B2(new_n322_), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n328_), .A2(new_n308_), .A3(new_n316_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n325_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n259_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT29), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n332_), .B2(KEYINPUT92), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT92), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n331_), .A2(new_n334_), .A3(KEYINPUT29), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n307_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT91), .B1(new_n325_), .B2(new_n329_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n317_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n324_), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT90), .B1(new_n328_), .B2(new_n308_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT91), .ZN(new_n342_));
  INV_X1    g141(.A(new_n329_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n337_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n307_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n346_), .B1(new_n331_), .B2(KEYINPUT29), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n306_), .B1(new_n336_), .B2(new_n349_), .ZN(new_n350_));
  AOI22_X1  g149(.A1(new_n292_), .A2(new_n293_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT92), .B1(new_n351_), .B2(new_n260_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n330_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n352_), .A2(new_n335_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(new_n346_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n355_), .A2(new_n305_), .A3(new_n348_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n303_), .B1(new_n350_), .B2(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n304_), .B1(new_n336_), .B2(new_n349_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(new_n356_), .A3(new_n303_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT94), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  AOI22_X1  g160(.A1(new_n354_), .A2(new_n346_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n302_), .B1(new_n362_), .B2(new_n305_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(KEYINPUT94), .A3(new_n358_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n357_), .B1(new_n361_), .B2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G1gat), .B(G29gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(G85gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT0), .B(G57gat), .ZN(new_n368_));
  XOR2_X1   g167(.A(new_n367_), .B(new_n368_), .Z(new_n369_));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(G127gat), .B(G134gat), .Z(new_n371_));
  XOR2_X1   g170(.A(G113gat), .B(G120gat), .Z(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  NAND3_X1  g172(.A1(new_n331_), .A2(KEYINPUT99), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n373_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n294_), .A2(new_n259_), .A3(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n374_), .A2(KEYINPUT4), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n331_), .A2(KEYINPUT99), .A3(new_n378_), .A4(new_n373_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n370_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n370_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n331_), .A2(new_n373_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n382_), .B2(new_n376_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n369_), .B1(new_n380_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT33), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT100), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT19), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n390_));
  INV_X1    g189(.A(G183gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT25), .ZN(new_n392_));
  INV_X1    g191(.A(G190gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT26), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n395_));
  AOI22_X1  g194(.A1(new_n390_), .A2(new_n392_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n396_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n391_), .A2(KEYINPUT25), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n393_), .A2(KEYINPUT26), .ZN(new_n399_));
  OAI211_X1 g198(.A(new_n398_), .B(new_n399_), .C1(new_n395_), .C2(new_n394_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G183gat), .A2(G190gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT23), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT24), .ZN(new_n404_));
  INV_X1    g203(.A(G169gat), .ZN(new_n405_));
  INV_X1    g204(.A(G176gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G169gat), .B(G176gat), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n403_), .B(new_n407_), .C1(new_n404_), .C2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n391_), .A2(new_n393_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n403_), .A2(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(new_n405_), .ZN(new_n413_));
  OAI22_X1  g212(.A1(new_n401_), .A2(new_n409_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n414_), .B1(new_n337_), .B2(new_n344_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n417_), .B(new_n403_), .C1(new_n408_), .C2(new_n416_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n398_), .A2(new_n392_), .ZN(new_n420_));
  AND3_X1   g219(.A1(new_n399_), .A2(KEYINPUT95), .A3(new_n394_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT95), .B1(new_n399_), .B2(new_n394_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n420_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  OR2_X1    g222(.A1(new_n413_), .A2(KEYINPUT97), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n413_), .A2(KEYINPUT97), .B1(new_n403_), .B2(new_n410_), .ZN(new_n425_));
  AOI22_X1  g224(.A1(new_n419_), .A2(new_n423_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT20), .B1(new_n330_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n389_), .B1(new_n415_), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G8gat), .B(G36gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT18), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G64gat), .B(G92gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n430_), .B(new_n431_), .Z(new_n432_));
  NAND3_X1  g231(.A1(new_n337_), .A2(new_n344_), .A3(new_n414_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT20), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(new_n330_), .B2(new_n426_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n389_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n428_), .A2(new_n432_), .A3(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n432_), .B1(new_n428_), .B2(new_n437_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT98), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n428_), .A2(new_n437_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n432_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT98), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n428_), .A2(new_n432_), .A3(new_n437_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n440_), .A2(new_n446_), .ZN(new_n447_));
  OAI211_X1 g246(.A(KEYINPUT33), .B(new_n369_), .C1(new_n380_), .C2(new_n383_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n369_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n382_), .A2(new_n376_), .A3(new_n381_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n377_), .A2(new_n379_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n449_), .B(new_n450_), .C1(new_n451_), .C2(new_n381_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n448_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT100), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n384_), .A2(new_n454_), .A3(new_n385_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n387_), .A2(new_n447_), .A3(new_n453_), .A4(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n383_), .B1(new_n451_), .B2(new_n381_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(new_n449_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n384_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n432_), .A2(KEYINPUT32), .ZN(new_n460_));
  OR3_X1    g259(.A1(new_n415_), .A2(new_n427_), .A3(new_n389_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n433_), .A2(new_n435_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(new_n389_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n460_), .B1(new_n461_), .B2(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n428_), .A2(new_n437_), .A3(new_n460_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n459_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n365_), .A2(new_n456_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n357_), .ZN(new_n469_));
  AND4_X1   g268(.A1(KEYINPUT94), .A2(new_n358_), .A3(new_n356_), .A4(new_n303_), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT94), .B1(new_n363_), .B2(new_n358_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n445_), .A2(KEYINPUT27), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n461_), .A2(new_n463_), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n432_), .B(KEYINPUT101), .Z(new_n475_));
  AOI21_X1  g274(.A(new_n473_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT27), .B1(new_n443_), .B2(new_n445_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n459_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n472_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G71gat), .B(G99gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(G43gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n414_), .B(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G227gat), .A2(G233gat), .ZN(new_n485_));
  INV_X1    g284(.A(G15gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n485_), .B(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT30), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n484_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT81), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n373_), .B(KEYINPUT31), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n493_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n468_), .A2(new_n481_), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n478_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n472_), .A2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n496_), .A2(new_n459_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n236_), .B1(new_n497_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT15), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n208_), .B(new_n503_), .ZN(new_n504_));
  XOR2_X1   g303(.A(G85gat), .B(G92gat), .Z(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT9), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT65), .B(G85gat), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT9), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n508_), .A3(G92gat), .ZN(new_n509_));
  OR2_X1    g308(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n510_));
  INV_X1    g309(.A(G106gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G99gat), .A2(G106gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT6), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT6), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(G99gat), .A3(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n506_), .A2(new_n509_), .A3(new_n513_), .A4(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT66), .ZN(new_n520_));
  INV_X1    g319(.A(G99gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n511_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT7), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT7), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n520_), .A2(new_n524_), .A3(new_n521_), .A4(new_n511_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n518_), .A3(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G85gat), .B(G92gat), .ZN(new_n528_));
  AND2_X1   g327(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n526_), .A2(new_n527_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n527_), .B1(new_n526_), .B2(new_n530_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n519_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n504_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n526_), .A2(new_n530_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n527_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n526_), .A2(new_n527_), .A3(new_n530_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n539_), .A2(new_n218_), .A3(new_n519_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G232gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT34), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n542_), .A2(KEYINPUT35), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n534_), .A2(new_n540_), .A3(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT74), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n534_), .A2(new_n540_), .A3(KEYINPUT74), .A4(new_n543_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n534_), .A2(new_n540_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n542_), .A2(KEYINPUT35), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n543_), .A2(new_n549_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n546_), .A2(new_n547_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G190gat), .B(G218gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT75), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G134gat), .B(G162gat), .ZN(new_n555_));
  XOR2_X1   g354(.A(new_n554_), .B(new_n555_), .Z(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n552_), .A2(KEYINPUT36), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT36), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n551_), .A2(KEYINPUT76), .A3(new_n561_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n561_), .B1(new_n551_), .B2(KEYINPUT76), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n558_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT37), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT37), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n558_), .B(new_n566_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n567_));
  INV_X1    g366(.A(G64gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(G57gat), .ZN(new_n569_));
  INV_X1    g368(.A(G57gat), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(G64gat), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n569_), .A2(new_n571_), .A3(KEYINPUT68), .ZN(new_n572_));
  AOI21_X1  g371(.A(KEYINPUT68), .B1(new_n569_), .B2(new_n571_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT11), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT68), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n570_), .A2(G64gat), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n568_), .A2(G57gat), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n575_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT11), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n569_), .A2(new_n571_), .A3(KEYINPUT68), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n578_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G71gat), .B(G78gat), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n574_), .A2(new_n581_), .A3(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(KEYINPUT11), .B(new_n582_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(new_n216_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(G231gat), .A2(G233gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(G127gat), .B(G155gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G183gat), .B(G211gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(KEYINPUT71), .A3(KEYINPUT17), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n590_), .A2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n597_), .B1(KEYINPUT17), .B2(new_n596_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n589_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n565_), .A2(new_n567_), .A3(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT13), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G230gat), .A2(G233gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(KEYINPUT64), .Z(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT69), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n584_), .A2(new_n585_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n607_), .B1(new_n608_), .B2(new_n533_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT70), .ZN(new_n610_));
  AND4_X1   g409(.A1(new_n506_), .A2(new_n509_), .A3(new_n513_), .A4(new_n518_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(KEYINPUT69), .A3(new_n586_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n609_), .A2(new_n610_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n608_), .A2(new_n533_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n610_), .B1(new_n609_), .B2(new_n613_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n606_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n586_), .A2(KEYINPUT71), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT71), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n584_), .A2(new_n620_), .A3(new_n585_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n619_), .A2(KEYINPUT12), .A3(new_n533_), .A4(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT12), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n623_), .B1(new_n612_), .B2(new_n586_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n539_), .A2(new_n586_), .A3(new_n519_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT72), .B1(new_n626_), .B2(new_n605_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT72), .ZN(new_n628_));
  AOI211_X1 g427(.A(new_n628_), .B(new_n606_), .C1(new_n612_), .C2(new_n586_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n625_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(G120gat), .B(G148gat), .Z(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n618_), .A2(new_n630_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n636_), .B1(new_n618_), .B2(new_n630_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n603_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n639_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n641_), .A2(KEYINPUT13), .A3(new_n637_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n602_), .A2(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n502_), .A2(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n211_), .A3(new_n459_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT38), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT102), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n647_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT104), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n500_), .A2(new_n365_), .A3(new_n478_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n496_), .ZN(new_n653_));
  AOI211_X1 g452(.A(new_n465_), .B(new_n464_), .C1(new_n458_), .C2(new_n384_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n384_), .A2(new_n454_), .A3(new_n385_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n454_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n448_), .A2(new_n452_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n440_), .B2(new_n446_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n654_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n653_), .B1(new_n660_), .B2(new_n365_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n652_), .B1(new_n661_), .B2(new_n481_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(new_n564_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n601_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n643_), .A2(new_n236_), .A3(new_n664_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n663_), .A2(KEYINPUT103), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(KEYINPUT103), .B1(new_n663_), .B2(new_n665_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G1gat), .B1(new_n668_), .B2(new_n479_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n649_), .A2(new_n651_), .A3(new_n669_), .ZN(G1324gat));
  NAND3_X1  g469(.A1(new_n645_), .A2(new_n212_), .A3(new_n498_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n663_), .A2(new_n498_), .A3(new_n665_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT39), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n672_), .A2(new_n673_), .A3(G8gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n672_), .B2(G8gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(G1325gat));
  OAI21_X1  g477(.A(G15gat), .B1(new_n668_), .B2(new_n496_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT41), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT41), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n681_), .B(G15gat), .C1(new_n668_), .C2(new_n496_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n645_), .A2(new_n486_), .A3(new_n653_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT105), .Z(new_n684_));
  NAND3_X1  g483(.A1(new_n680_), .A2(new_n682_), .A3(new_n684_), .ZN(G1326gat));
  INV_X1    g484(.A(G22gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n645_), .A2(new_n686_), .A3(new_n472_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n472_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n688_), .A2(new_n689_), .A3(G22gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n688_), .B2(G22gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(G1327gat));
  INV_X1    g491(.A(new_n643_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(new_n235_), .A3(new_n664_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n497_), .A2(new_n501_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n565_), .A2(new_n567_), .ZN(new_n698_));
  XOR2_X1   g497(.A(new_n698_), .B(KEYINPUT106), .Z(new_n699_));
  AOI21_X1  g498(.A(new_n696_), .B1(new_n697_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n696_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n497_), .B2(new_n501_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT44), .B(new_n695_), .C1(new_n700_), .C2(new_n702_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n698_), .B(KEYINPUT106), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT43), .B1(new_n662_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n702_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n694_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n703_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(G29gat), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n479_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n564_), .A2(new_n664_), .A3(KEYINPUT108), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT108), .B1(new_n564_), .B2(new_n664_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n693_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  AOI211_X1 g513(.A(new_n236_), .B(new_n714_), .C1(new_n497_), .C2(new_n501_), .ZN(new_n715_));
  AOI21_X1  g514(.A(G29gat), .B1(new_n715_), .B2(new_n459_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n711_), .A2(new_n716_), .ZN(G1328gat));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n718_), .A2(KEYINPUT109), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n498_), .B(new_n703_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G36gat), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n718_), .A2(KEYINPUT109), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT45), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n478_), .A2(G36gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n715_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n714_), .ZN(new_n727_));
  AND4_X1   g526(.A1(new_n724_), .A2(new_n502_), .A3(new_n727_), .A4(new_n725_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n723_), .B1(new_n726_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n720_), .B1(new_n722_), .B2(new_n730_), .ZN(new_n731_));
  AOI211_X1 g530(.A(new_n719_), .B(new_n729_), .C1(new_n721_), .C2(G36gat), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1329gat));
  INV_X1    g532(.A(G43gat), .ZN(new_n734_));
  INV_X1    g533(.A(new_n715_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(new_n496_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n653_), .A2(G43gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n709_), .B2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g538(.A1(new_n735_), .A2(G50gat), .A3(new_n365_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n472_), .B(new_n703_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n742_));
  AND3_X1   g541(.A1(new_n741_), .A2(new_n742_), .A3(G50gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n742_), .B1(new_n741_), .B2(G50gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1331gat));
  NOR3_X1   g544(.A1(new_n693_), .A2(new_n235_), .A3(new_n664_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n663_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n459_), .A2(G57gat), .ZN(new_n748_));
  OR3_X1    g547(.A1(new_n747_), .A2(KEYINPUT111), .A3(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n693_), .A2(new_n235_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n697_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n698_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n601_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n570_), .B1(new_n753_), .B2(new_n479_), .ZN(new_n754_));
  OAI21_X1  g553(.A(KEYINPUT111), .B1(new_n747_), .B2(new_n748_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n749_), .A2(new_n754_), .A3(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n756_), .B(new_n757_), .ZN(G1332gat));
  OAI21_X1  g557(.A(G64gat), .B1(new_n747_), .B2(new_n478_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT48), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n498_), .A2(new_n568_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n753_), .B2(new_n761_), .ZN(G1333gat));
  OAI21_X1  g561(.A(G71gat), .B1(new_n747_), .B2(new_n496_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT49), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n496_), .A2(G71gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n753_), .B2(new_n765_), .ZN(G1334gat));
  OAI21_X1  g565(.A(G78gat), .B1(new_n747_), .B2(new_n365_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT50), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n365_), .A2(G78gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n753_), .B2(new_n769_), .ZN(G1335gat));
  OR2_X1    g569(.A1(new_n712_), .A2(new_n713_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n751_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(G85gat), .B1(new_n772_), .B2(new_n459_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n750_), .A2(new_n664_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT113), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT113), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n750_), .A2(new_n776_), .A3(new_n664_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n778_), .B1(new_n700_), .B2(new_n702_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT114), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  OAI211_X1 g580(.A(KEYINPUT114), .B(new_n778_), .C1(new_n700_), .C2(new_n702_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n459_), .A2(new_n507_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n773_), .B1(new_n783_), .B2(new_n784_), .ZN(G1336gat));
  INV_X1    g584(.A(G92gat), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n772_), .A2(new_n786_), .A3(new_n498_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n478_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n786_), .ZN(G1337gat));
  NAND4_X1  g588(.A1(new_n772_), .A2(new_n653_), .A3(new_n510_), .A4(new_n512_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n496_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n521_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT51), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT51), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(new_n790_), .C1(new_n791_), .C2(new_n521_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(G1338gat));
  NAND3_X1  g595(.A1(new_n772_), .A2(new_n511_), .A3(new_n472_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n472_), .B(new_n778_), .C1(new_n700_), .C2(new_n702_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(G106gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n798_), .B2(G106gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n797_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT53), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT53), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n804_), .B(new_n797_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1339gat));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n644_), .B2(new_n236_), .ZN(new_n808_));
  NOR4_X1   g607(.A1(new_n602_), .A2(new_n643_), .A3(KEYINPUT54), .A4(new_n235_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n228_), .B1(new_n222_), .B2(new_n220_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n217_), .A2(new_n219_), .A3(new_n223_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n232_), .A2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n622_), .A2(new_n609_), .A3(new_n624_), .A4(new_n613_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n606_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n629_), .A2(new_n627_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n622_), .A2(new_n624_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n820_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n625_), .B(KEYINPUT55), .C1(new_n627_), .C2(new_n629_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n816_), .A2(KEYINPUT115), .A3(new_n606_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n819_), .A2(new_n823_), .A3(new_n824_), .A4(new_n825_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n826_), .A2(KEYINPUT56), .A3(new_n635_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT56), .B1(new_n826_), .B2(new_n635_), .ZN(new_n828_));
  NOR3_X1   g627(.A1(new_n827_), .A2(new_n828_), .A3(KEYINPUT116), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n235_), .A2(new_n637_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n826_), .A2(new_n635_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n815_), .B1(new_n829_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n564_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(KEYINPUT57), .A3(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n637_), .A2(new_n814_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n826_), .A2(KEYINPUT56), .A3(new_n635_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n834_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(KEYINPUT58), .B1(new_n842_), .B2(KEYINPUT117), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT117), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n827_), .A2(new_n828_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n844_), .B(new_n845_), .C1(new_n846_), .C2(new_n840_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n843_), .A2(new_n847_), .A3(new_n698_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849_));
  INV_X1    g648(.A(new_n815_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n834_), .A2(new_n835_), .A3(new_n841_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n830_), .B1(new_n828_), .B2(KEYINPUT116), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n849_), .B1(new_n853_), .B2(new_n564_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n839_), .A2(new_n848_), .A3(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n810_), .B1(new_n855_), .B2(new_n664_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n499_), .A2(new_n459_), .A3(new_n653_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(G113gat), .B1(new_n858_), .B2(new_n235_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n855_), .A2(new_n664_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n810_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n857_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT59), .B1(new_n863_), .B2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n856_), .A2(new_n866_), .A3(new_n857_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n860_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n863_), .A2(KEYINPUT59), .A3(new_n864_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n866_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(KEYINPUT118), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n868_), .A2(new_n871_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n236_), .A2(KEYINPUT119), .ZN(new_n873_));
  MUX2_X1   g672(.A(KEYINPUT119), .B(new_n873_), .S(G113gat), .Z(new_n874_));
  AOI21_X1  g673(.A(new_n859_), .B1(new_n872_), .B2(new_n874_), .ZN(G1340gat));
  XNOR2_X1  g674(.A(KEYINPUT120), .B(G120gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n876_), .B1(new_n693_), .B2(KEYINPUT60), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n858_), .B(new_n877_), .C1(KEYINPUT60), .C2(new_n876_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n693_), .B1(new_n869_), .B2(new_n870_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n876_), .ZN(G1341gat));
  INV_X1    g679(.A(G127gat), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n858_), .A2(new_n881_), .A3(new_n601_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n664_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n882_), .B1(new_n883_), .B2(new_n881_), .ZN(G1342gat));
  AOI21_X1  g683(.A(G134gat), .B1(new_n858_), .B2(new_n564_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT121), .B(G134gat), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n752_), .A2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n872_), .B2(new_n887_), .ZN(G1343gat));
  NOR4_X1   g687(.A1(new_n365_), .A2(new_n653_), .A3(new_n498_), .A4(new_n479_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n863_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n236_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(new_n237_), .ZN(G1344gat));
  NOR2_X1   g691(.A1(new_n890_), .A2(new_n693_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(new_n238_), .ZN(G1345gat));
  AND2_X1   g693(.A1(new_n863_), .A2(new_n889_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT123), .Z(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n895_), .A2(new_n601_), .A3(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n897_), .B1(new_n890_), .B2(new_n664_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(KEYINPUT122), .B(KEYINPUT124), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n899_), .A2(new_n902_), .A3(new_n900_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1346gat));
  AOI21_X1  g705(.A(G162gat), .B1(new_n895_), .B2(new_n564_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n890_), .A2(new_n249_), .A3(new_n704_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1347gat));
  NAND3_X1  g708(.A1(new_n500_), .A2(new_n365_), .A3(new_n498_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n856_), .A2(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT22), .B(G169gat), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n235_), .A2(new_n912_), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n913_), .B(KEYINPUT125), .Z(new_n914_));
  NAND2_X1  g713(.A1(new_n911_), .A2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n911_), .A2(new_n235_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(G169gat), .ZN(new_n918_));
  AOI211_X1 g717(.A(KEYINPUT62), .B(new_n405_), .C1(new_n911_), .C2(new_n235_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n915_), .B1(new_n918_), .B2(new_n919_), .ZN(G1348gat));
  XNOR2_X1  g719(.A(KEYINPUT126), .B(G176gat), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n406_), .A2(KEYINPUT126), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n911_), .A2(new_n643_), .ZN(new_n923_));
  MUX2_X1   g722(.A(new_n921_), .B(new_n922_), .S(new_n923_), .Z(G1349gat));
  NAND2_X1  g723(.A1(new_n911_), .A2(new_n601_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n420_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n926_), .B1(new_n391_), .B2(new_n925_), .ZN(G1350gat));
  OAI211_X1 g726(.A(new_n911_), .B(new_n564_), .C1(new_n421_), .C2(new_n422_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n856_), .A2(new_n752_), .A3(new_n910_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n928_), .B1(new_n929_), .B2(new_n393_), .ZN(G1351gat));
  NOR4_X1   g729(.A1(new_n365_), .A2(new_n653_), .A3(new_n478_), .A4(new_n459_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n863_), .A2(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n932_), .A2(new_n236_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(new_n322_), .ZN(G1352gat));
  NOR2_X1   g733(.A1(new_n932_), .A2(new_n693_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(G204gat), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n936_), .B1(new_n314_), .B2(new_n935_), .ZN(G1353gat));
  NOR2_X1   g736(.A1(new_n932_), .A2(new_n664_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  XOR2_X1   g739(.A(KEYINPUT63), .B(G211gat), .Z(new_n941_));
  NOR3_X1   g740(.A1(new_n932_), .A2(new_n664_), .A3(new_n941_), .ZN(new_n942_));
  OAI21_X1  g741(.A(KEYINPUT127), .B1(new_n940_), .B2(new_n942_), .ZN(new_n943_));
  OR3_X1    g742(.A1(new_n932_), .A2(new_n664_), .A3(new_n941_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945_));
  OAI211_X1 g744(.A(new_n944_), .B(new_n945_), .C1(new_n938_), .C2(new_n939_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n943_), .A2(new_n946_), .ZN(G1354gat));
  OAI21_X1  g746(.A(G218gat), .B1(new_n932_), .B2(new_n752_), .ZN(new_n948_));
  OR2_X1    g747(.A1(new_n838_), .A2(G218gat), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n932_), .B2(new_n949_), .ZN(G1355gat));
endmodule


