//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n608_, new_n609_, new_n610_, new_n611_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n869_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT7), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT6), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .A4(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT65), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G85gat), .ZN(new_n218_));
  INV_X1    g017(.A(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT65), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(new_n214_), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n212_), .A2(new_n213_), .A3(new_n217_), .A4(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT66), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n212_), .A2(KEYINPUT66), .A3(new_n217_), .A4(new_n222_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(KEYINPUT8), .A3(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G57gat), .B(G64gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n229_));
  XOR2_X1   g028(.A(G71gat), .B(G78gat), .Z(new_n230_));
  OR2_X1    g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n228_), .A2(KEYINPUT11), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n230_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n231_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  XOR2_X1   g033(.A(KEYINPUT10), .B(G99gat), .Z(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n205_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n220_), .A2(KEYINPUT9), .A3(new_n214_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n209_), .A2(new_n210_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n214_), .A2(KEYINPUT9), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .A4(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT8), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n223_), .A2(new_n224_), .A3(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n227_), .A2(new_n234_), .A3(new_n240_), .A4(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G230gat), .ZN(new_n244_));
  INV_X1    g043(.A(G233gat), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n243_), .A2(new_n247_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n223_), .A2(new_n224_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n226_), .A2(KEYINPUT8), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n240_), .B(new_n242_), .C1(new_n249_), .C2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT12), .ZN(new_n252_));
  INV_X1    g051(.A(new_n234_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n252_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n248_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT68), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n248_), .B(new_n258_), .C1(new_n254_), .C2(new_n255_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n251_), .A2(new_n253_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT67), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(new_n243_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n251_), .A2(KEYINPUT67), .A3(new_n253_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n262_), .A2(new_n246_), .A3(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n257_), .A2(new_n259_), .A3(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G120gat), .B(G148gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT5), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G176gat), .B(G204gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(new_n268_), .Z(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n257_), .A2(new_n271_), .A3(new_n259_), .A4(new_n264_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT13), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n270_), .A2(KEYINPUT13), .A3(new_n272_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G29gat), .B(G36gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G43gat), .B(G50gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G1gat), .B(G8gat), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n283_), .A2(KEYINPUT72), .ZN(new_n284_));
  INV_X1    g083(.A(G8gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G15gat), .B(G22gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(KEYINPUT72), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n284_), .A2(new_n286_), .A3(new_n287_), .A4(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n283_), .B(KEYINPUT72), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n286_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n282_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G229gat), .A2(G233gat), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n281_), .B(KEYINPUT15), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n292_), .A2(new_n289_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n296_), .A2(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n298_), .A2(new_n281_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n295_), .B1(new_n302_), .B2(new_n293_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G113gat), .B(G141gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G169gat), .B(G197gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n305_), .B(new_n306_), .Z(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n304_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n301_), .A2(new_n303_), .A3(new_n307_), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n309_), .A2(KEYINPUT74), .A3(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT74), .B1(new_n309_), .B2(new_n310_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n278_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT101), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G231gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n234_), .B(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(new_n299_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G127gat), .B(G155gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(G183gat), .B(G211gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT17), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n318_), .A2(new_n324_), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n323_), .A2(KEYINPUT17), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n318_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n315_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G190gat), .B(G218gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G134gat), .B(G162gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n332_), .B(KEYINPUT36), .Z(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G232gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT35), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  AND2_X1   g138(.A1(new_n251_), .A2(new_n297_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n227_), .A2(new_n281_), .A3(new_n240_), .A4(new_n242_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n338_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n339_), .B1(new_n340_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n251_), .A2(new_n297_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n339_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(new_n342_), .A4(new_n341_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n334_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n332_), .A2(KEYINPUT36), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(new_n347_), .A3(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT70), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n344_), .A2(KEYINPUT70), .A3(new_n347_), .A4(new_n349_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n348_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G127gat), .B(G134gat), .Z(new_n355_));
  XOR2_X1   g154(.A(G113gat), .B(G120gat), .Z(new_n356_));
  XOR2_X1   g155(.A(new_n355_), .B(new_n356_), .Z(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G227gat), .A2(G233gat), .ZN(new_n359_));
  INV_X1    g158(.A(G71gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(G99gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G15gat), .B(G43gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT80), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n362_), .B(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(KEYINPUT78), .B(KEYINPUT79), .Z(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G183gat), .A2(G190gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT23), .ZN(new_n369_));
  INV_X1    g168(.A(G169gat), .ZN(new_n370_));
  INV_X1    g169(.A(G176gat), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n369_), .B1(KEYINPUT24), .B2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(KEYINPUT24), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n373_), .B1(KEYINPUT76), .B2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT25), .B(G183gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(KEYINPUT26), .B(G190gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT75), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n375_), .A2(KEYINPUT76), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n376_), .A2(new_n381_), .A3(new_n382_), .ZN(new_n383_));
  OR2_X1    g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n369_), .A2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT22), .B(G169gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n371_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n374_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n388_), .A2(KEYINPUT77), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(KEYINPUT77), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n385_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n383_), .A2(new_n391_), .A3(KEYINPUT30), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT30), .B1(new_n383_), .B2(new_n391_), .ZN(new_n394_));
  OAI21_X1  g193(.A(KEYINPUT81), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n394_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT81), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n396_), .A2(new_n397_), .A3(new_n392_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n367_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n398_), .A2(new_n367_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT31), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n367_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(new_n393_), .A2(KEYINPUT81), .A3(new_n394_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n397_), .B1(new_n396_), .B2(new_n392_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT31), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n398_), .A2(new_n367_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT82), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n401_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n409_), .B1(new_n401_), .B2(new_n408_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n358_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n401_), .A2(new_n408_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT82), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n401_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n414_), .A2(new_n357_), .A3(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n412_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT93), .ZN(new_n418_));
  XNOR2_X1  g217(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G226gat), .A2(G233gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT89), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n377_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n378_), .B(KEYINPUT90), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n375_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n373_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT91), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n386_), .B(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(new_n371_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n369_), .A2(new_n384_), .B1(G169gat), .B2(G176gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n428_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G211gat), .B(G218gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT87), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G197gat), .B(G204gat), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT21), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n438_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n436_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT87), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n435_), .B(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n439_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n445_), .ZN(new_n446_));
  OAI211_X1 g245(.A(KEYINPUT20), .B(new_n421_), .C1(new_n434_), .C2(new_n446_), .ZN(new_n447_));
  AND2_X1   g246(.A1(new_n442_), .A2(new_n445_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n448_), .B1(new_n391_), .B2(new_n383_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n418_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n383_), .A2(new_n391_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n446_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n421_), .A2(KEYINPUT20), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n425_), .A2(new_n427_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n453_), .B1(new_n454_), .B2(new_n448_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n455_), .A3(KEYINPUT93), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n450_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n421_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n448_), .A2(new_n383_), .A3(new_n391_), .ZN(new_n459_));
  OAI21_X1  g258(.A(KEYINPUT20), .B1(new_n454_), .B2(new_n448_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n458_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT92), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G8gat), .B(G36gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT18), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G64gat), .B(G92gat), .ZN(new_n466_));
  XOR2_X1   g265(.A(new_n465_), .B(new_n466_), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n434_), .A2(new_n446_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n468_), .B(KEYINPUT20), .C1(new_n451_), .C2(new_n446_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(KEYINPUT92), .A3(new_n458_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n457_), .A2(new_n463_), .A3(new_n467_), .A4(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT99), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n450_), .A2(new_n456_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT99), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(new_n467_), .A4(new_n470_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT27), .ZN(new_n476_));
  XOR2_X1   g275(.A(KEYINPUT98), .B(KEYINPUT20), .Z(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n434_), .B2(new_n446_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n458_), .B1(new_n479_), .B2(new_n449_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n480_), .B1(new_n469_), .B2(new_n458_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n467_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n476_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n472_), .A2(new_n475_), .A3(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n457_), .A2(new_n463_), .A3(new_n470_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n482_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT27), .B1(new_n486_), .B2(new_n471_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT100), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n467_), .B1(new_n473_), .B2(new_n470_), .ZN(new_n489_));
  AND4_X1   g288(.A1(new_n467_), .A2(new_n457_), .A3(new_n463_), .A4(new_n470_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n476_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n472_), .A2(new_n475_), .A3(new_n483_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT100), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n488_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT83), .B(KEYINPUT84), .ZN(new_n496_));
  NOR2_X1   g295(.A1(G155gat), .A2(G162gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G155gat), .A2(G162gat), .ZN(new_n499_));
  XOR2_X1   g298(.A(new_n499_), .B(KEYINPUT1), .Z(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(G141gat), .ZN(new_n502_));
  INV_X1    g301(.A(G148gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(G141gat), .A2(G148gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  OR2_X1    g305(.A1(new_n504_), .A2(KEYINPUT3), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT2), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n505_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n504_), .A2(KEYINPUT3), .ZN(new_n511_));
  NAND4_X1  g310(.A1(new_n507_), .A2(new_n509_), .A3(new_n510_), .A4(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n498_), .A2(new_n499_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n506_), .A2(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n448_), .B1(new_n514_), .B2(KEYINPUT29), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  XNOR2_X1  g316(.A(G22gat), .B(G50gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT86), .ZN(new_n519_));
  OR3_X1    g318(.A1(new_n514_), .A2(KEYINPUT29), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G228gat), .A2(G233gat), .ZN(new_n521_));
  INV_X1    g320(.A(G78gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(new_n205_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n519_), .B1(new_n514_), .B2(KEYINPUT29), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n520_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n520_), .B2(new_n526_), .ZN(new_n528_));
  OR3_X1    g327(.A1(new_n517_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n517_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AND2_X1   g330(.A1(new_n498_), .A2(new_n500_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n504_), .A2(new_n505_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n513_), .B(KEYINPUT94), .C1(new_n532_), .C2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n358_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n506_), .A2(KEYINPUT94), .A3(new_n357_), .A4(new_n513_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT4), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G225gat), .A2(G233gat), .ZN(new_n539_));
  XOR2_X1   g338(.A(new_n539_), .B(KEYINPUT95), .Z(new_n540_));
  NOR2_X1   g339(.A1(new_n358_), .A2(KEYINPUT4), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n514_), .A2(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n538_), .A2(new_n540_), .A3(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n537_), .A2(new_n539_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G1gat), .B(G29gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(G85gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT0), .B(G57gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(new_n548_), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n545_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n543_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n417_), .A2(new_n495_), .A3(new_n531_), .A4(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n412_), .A2(new_n416_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n531_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n489_), .A2(new_n490_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n537_), .A2(KEYINPUT96), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT96), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n535_), .A2(new_n560_), .A3(new_n536_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n559_), .A2(new_n540_), .A3(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n538_), .A2(new_n539_), .A3(new_n542_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(new_n563_), .A3(new_n550_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT97), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n562_), .A2(new_n563_), .A3(KEYINPUT97), .A4(new_n550_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n543_), .A2(KEYINPUT33), .A3(new_n544_), .A4(new_n549_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT33), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n552_), .A2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n558_), .A2(new_n568_), .A3(new_n569_), .A4(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n481_), .A2(KEYINPUT32), .A3(new_n467_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n467_), .A2(KEYINPUT32), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n473_), .A2(new_n574_), .A3(new_n470_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n553_), .A2(new_n573_), .A3(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n557_), .B1(new_n572_), .B2(new_n576_), .ZN(new_n577_));
  AND4_X1   g376(.A1(new_n557_), .A2(new_n491_), .A3(new_n492_), .A4(new_n554_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n556_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n354_), .B1(new_n555_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n329_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n202_), .B1(new_n582_), .B2(new_n553_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT38), .ZN(new_n584_));
  INV_X1    g383(.A(new_n313_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n555_), .B2(new_n579_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n328_), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT37), .B1(new_n348_), .B2(KEYINPUT71), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n354_), .A2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n354_), .A2(new_n588_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n587_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(new_n277_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n586_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(new_n202_), .A3(new_n553_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n583_), .B1(new_n584_), .B2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n595_), .B1(new_n584_), .B2(new_n594_), .ZN(G1324gat));
  INV_X1    g395(.A(new_n495_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n593_), .A2(new_n285_), .A3(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(G8gat), .B1(new_n581_), .B2(new_n495_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n599_), .A2(KEYINPUT39), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(KEYINPUT39), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n598_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n598_), .B(new_n603_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(G1325gat));
  OAI21_X1  g406(.A(G15gat), .B1(new_n581_), .B2(new_n556_), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n608_), .B(KEYINPUT41), .Z(new_n609_));
  INV_X1    g408(.A(G15gat), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n593_), .A2(new_n610_), .A3(new_n417_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(G1326gat));
  XNOR2_X1  g411(.A(new_n531_), .B(KEYINPUT103), .ZN(new_n613_));
  OAI21_X1  g412(.A(G22gat), .B1(new_n581_), .B2(new_n613_), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT42), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n613_), .A2(G22gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT104), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n593_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(G1327gat));
  INV_X1    g418(.A(G29gat), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n315_), .A2(new_n587_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n354_), .A2(new_n588_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n354_), .A2(new_n588_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  AOI211_X1 g423(.A(KEYINPUT43), .B(new_n624_), .C1(new_n555_), .C2(new_n579_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT43), .ZN(new_n626_));
  INV_X1    g425(.A(new_n568_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n571_), .A2(new_n486_), .A3(new_n569_), .A4(new_n471_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n576_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n491_), .A2(new_n492_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n531_), .A2(new_n553_), .ZN(new_n631_));
  AOI22_X1  g430(.A1(new_n629_), .A2(new_n531_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n491_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n493_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n531_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n412_), .A2(new_n416_), .A3(new_n554_), .ZN(new_n636_));
  OAI22_X1  g435(.A1(new_n632_), .A2(new_n417_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n624_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n626_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n621_), .B1(new_n625_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT44), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(KEYINPUT44), .B(new_n621_), .C1(new_n625_), .C2(new_n639_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(new_n553_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT105), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n620_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n646_), .B1(new_n645_), .B2(new_n644_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n354_), .A2(new_n328_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n277_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n586_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(new_n620_), .A3(new_n553_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n647_), .A2(new_n652_), .ZN(G1328gat));
  NOR2_X1   g452(.A1(new_n495_), .A2(G36gat), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n637_), .A2(new_n313_), .A3(new_n649_), .A4(new_n654_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n655_), .A2(KEYINPUT45), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(KEYINPUT45), .ZN(new_n657_));
  OAI22_X1  g456(.A1(new_n656_), .A2(new_n657_), .B1(KEYINPUT106), .B2(KEYINPUT46), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n642_), .A2(new_n597_), .A3(new_n643_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n659_), .B2(G36gat), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT46), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n660_), .B(new_n663_), .ZN(G1329gat));
  INV_X1    g463(.A(G43gat), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n556_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n642_), .A2(new_n643_), .A3(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n665_), .B1(new_n650_), .B2(new_n556_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT107), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n642_), .A2(new_n669_), .A3(new_n643_), .A4(new_n666_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n671_), .A2(new_n672_), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n672_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1330gat));
  INV_X1    g475(.A(new_n613_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G50gat), .B1(new_n651_), .B2(new_n677_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n642_), .A2(new_n643_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n557_), .A2(G50gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(G1331gat));
  AOI21_X1  g480(.A(new_n313_), .B1(new_n555_), .B2(new_n579_), .ZN(new_n682_));
  AND4_X1   g481(.A1(new_n277_), .A2(new_n682_), .A3(new_n587_), .A4(new_n624_), .ZN(new_n683_));
  INV_X1    g482(.A(G57gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n683_), .A2(new_n684_), .A3(new_n553_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n580_), .A2(new_n585_), .A3(new_n277_), .A4(new_n587_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n686_), .A2(KEYINPUT109), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(KEYINPUT109), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(new_n553_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n685_), .B1(new_n690_), .B2(new_n684_), .ZN(G1332gat));
  NOR2_X1   g490(.A1(new_n495_), .A2(G64gat), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT110), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n683_), .A2(new_n693_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n687_), .A2(new_n597_), .A3(new_n688_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT48), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n695_), .A2(new_n696_), .A3(G64gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n695_), .B2(G64gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(G1333gat));
  NAND3_X1  g498(.A1(new_n683_), .A2(new_n360_), .A3(new_n417_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n687_), .A2(new_n417_), .A3(new_n688_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT49), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n701_), .A2(new_n702_), .A3(G71gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n701_), .B2(G71gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n700_), .B1(new_n703_), .B2(new_n704_), .ZN(G1334gat));
  NAND3_X1  g504(.A1(new_n683_), .A2(new_n522_), .A3(new_n677_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n687_), .A2(new_n677_), .A3(new_n688_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT50), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(G78gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n707_), .B2(G78gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(G1335gat));
  NOR2_X1   g510(.A1(new_n278_), .A2(new_n648_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n682_), .A2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n713_), .A2(new_n218_), .A3(new_n553_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n277_), .A2(new_n585_), .A3(new_n328_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n637_), .A2(new_n638_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT43), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n637_), .A2(new_n626_), .A3(new_n638_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(KEYINPUT111), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT111), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n720_), .B1(new_n625_), .B2(new_n639_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n715_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n722_), .A2(new_n553_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n714_), .B1(new_n723_), .B2(new_n218_), .ZN(G1336gat));
  AOI21_X1  g523(.A(G92gat), .B1(new_n713_), .B2(new_n597_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT112), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n495_), .A2(new_n219_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n722_), .B2(new_n727_), .ZN(G1337gat));
  AOI21_X1  g527(.A(new_n204_), .B1(new_n722_), .B2(new_n417_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n417_), .A2(new_n235_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n713_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  OR3_X1    g531(.A1(new_n729_), .A2(KEYINPUT51), .A3(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(KEYINPUT51), .B1(new_n729_), .B2(new_n732_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1338gat));
  INV_X1    g534(.A(KEYINPUT114), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n715_), .A2(new_n531_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n736_), .B1(new_n738_), .B2(new_n205_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n625_), .A2(new_n639_), .ZN(new_n740_));
  OAI211_X1 g539(.A(KEYINPUT114), .B(G106gat), .C1(new_n740_), .C2(new_n737_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n739_), .A2(KEYINPUT52), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT52), .ZN(new_n743_));
  OAI211_X1 g542(.A(new_n736_), .B(new_n743_), .C1(new_n738_), .C2(new_n205_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n682_), .A2(new_n205_), .A3(new_n557_), .A4(new_n712_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT113), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(new_n744_), .A3(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT53), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n742_), .A2(new_n749_), .A3(new_n744_), .A4(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(G1339gat));
  INV_X1    g550(.A(KEYINPUT118), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n313_), .A2(G113gat), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT117), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT116), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n299_), .A2(new_n282_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n293_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n307_), .B1(new_n759_), .B2(new_n294_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n300_), .A2(new_n758_), .A3(new_n295_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n310_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n272_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n257_), .A2(new_n766_), .A3(new_n259_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n243_), .A2(new_n247_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n260_), .A2(KEYINPUT12), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n768_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n243_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n772_));
  AOI22_X1  g571(.A1(KEYINPUT55), .A2(new_n771_), .B1(new_n772_), .B2(new_n246_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n767_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT56), .B1(new_n774_), .B2(new_n269_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT56), .ZN(new_n776_));
  AOI211_X1 g575(.A(new_n776_), .B(new_n271_), .C1(new_n767_), .C2(new_n773_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n765_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT58), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  OAI211_X1 g579(.A(KEYINPUT58), .B(new_n765_), .C1(new_n775_), .C2(new_n777_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n638_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT115), .B1(new_n273_), .B2(new_n764_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n784_), .B(new_n763_), .C1(new_n270_), .C2(new_n272_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n313_), .A2(new_n272_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n787_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n354_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n782_), .B1(new_n789_), .B2(KEYINPUT57), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n273_), .A2(new_n764_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n784_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n273_), .A2(KEYINPUT115), .A3(new_n764_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n788_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n354_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n794_), .A2(KEYINPUT57), .A3(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n328_), .B1(new_n790_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n592_), .B2(new_n585_), .ZN(new_n800_));
  NOR4_X1   g599(.A1(new_n591_), .A2(new_n277_), .A3(KEYINPUT54), .A4(new_n313_), .ZN(new_n801_));
  OR2_X1    g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n798_), .A2(new_n802_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n635_), .A2(new_n556_), .A3(new_n554_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT59), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT59), .ZN(new_n806_));
  INV_X1    g605(.A(new_n804_), .ZN(new_n807_));
  AOI211_X1 g606(.A(new_n806_), .B(new_n807_), .C1(new_n798_), .C2(new_n802_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n756_), .B1(new_n805_), .B2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n800_), .A2(new_n801_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n794_), .A2(new_n795_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n813_), .A2(new_n796_), .A3(new_n782_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n810_), .B1(new_n814_), .B2(new_n328_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n806_), .B1(new_n815_), .B2(new_n807_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n624_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n811_), .A2(new_n812_), .B1(new_n781_), .B2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n587_), .B1(new_n818_), .B2(new_n796_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT59), .B(new_n804_), .C1(new_n819_), .C2(new_n810_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n816_), .A2(KEYINPUT116), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n755_), .B1(new_n809_), .B2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n815_), .A2(new_n807_), .ZN(new_n823_));
  AOI21_X1  g622(.A(G113gat), .B1(new_n823_), .B2(new_n313_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n752_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n816_), .A2(KEYINPUT116), .A3(new_n820_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT116), .B1(new_n816_), .B2(new_n820_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n754_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n824_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n828_), .A2(KEYINPUT118), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n825_), .A2(new_n830_), .ZN(G1340gat));
  INV_X1    g630(.A(G120gat), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(KEYINPUT60), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n278_), .B2(KEYINPUT60), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n834_), .B2(KEYINPUT119), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n823_), .B(new_n835_), .C1(KEYINPUT119), .C2(new_n834_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n278_), .B1(new_n816_), .B2(new_n820_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n832_), .ZN(G1341gat));
  AND2_X1   g637(.A1(new_n587_), .A2(G127gat), .ZN(new_n839_));
  OAI22_X1  g638(.A1(new_n826_), .A2(new_n827_), .B1(KEYINPUT120), .B2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(new_n587_), .A3(new_n823_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n842_), .B(new_n839_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(G127gat), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n841_), .A2(new_n844_), .ZN(G1342gat));
  INV_X1    g644(.A(KEYINPUT122), .ZN(new_n846_));
  INV_X1    g645(.A(G134gat), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n624_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n809_), .B2(new_n821_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n803_), .A2(new_n354_), .A3(new_n804_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n847_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT121), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(new_n854_), .A3(new_n847_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n846_), .B1(new_n850_), .B2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n848_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n858_));
  AND3_X1   g657(.A1(new_n851_), .A2(new_n854_), .A3(new_n847_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n854_), .B1(new_n851_), .B2(new_n847_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n858_), .A2(KEYINPUT122), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n857_), .A2(new_n862_), .ZN(G1343gat));
  NOR3_X1   g662(.A1(new_n815_), .A2(new_n417_), .A3(new_n531_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n597_), .A2(new_n554_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n866_), .A2(new_n585_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(new_n502_), .ZN(G1344gat));
  NOR2_X1   g667(.A1(new_n866_), .A2(new_n278_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n503_), .ZN(G1345gat));
  NAND3_X1  g669(.A1(new_n864_), .A2(new_n587_), .A3(new_n865_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT123), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n864_), .A2(new_n873_), .A3(new_n587_), .A4(new_n865_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT61), .B(G155gat), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n872_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1346gat));
  INV_X1    g677(.A(G162gat), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n866_), .A2(new_n879_), .A3(new_n624_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n866_), .B2(new_n795_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(KEYINPUT124), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n883_), .B(new_n879_), .C1(new_n866_), .C2(new_n795_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n880_), .B1(new_n882_), .B2(new_n884_), .ZN(G1347gat));
  INV_X1    g684(.A(KEYINPUT62), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n495_), .A2(new_n553_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n417_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT125), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n889_), .A2(new_n803_), .A3(new_n613_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n585_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n886_), .B1(new_n891_), .B2(new_n370_), .ZN(new_n892_));
  OAI211_X1 g691(.A(KEYINPUT62), .B(G169gat), .C1(new_n890_), .C2(new_n585_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n430_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n892_), .A2(new_n893_), .A3(new_n894_), .ZN(G1348gat));
  INV_X1    g694(.A(new_n890_), .ZN(new_n896_));
  AOI21_X1  g695(.A(G176gat), .B1(new_n896_), .B2(new_n277_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n815_), .A2(new_n557_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n889_), .A2(G176gat), .A3(new_n277_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(G1349gat));
  NOR3_X1   g699(.A1(new_n890_), .A2(new_n423_), .A3(new_n328_), .ZN(new_n901_));
  INV_X1    g700(.A(G183gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n898_), .A2(new_n889_), .A3(new_n587_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n896_), .A2(new_n424_), .A3(new_n354_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G190gat), .B1(new_n890_), .B2(new_n624_), .ZN(new_n906_));
  AND2_X1   g705(.A1(new_n906_), .A2(KEYINPUT126), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n906_), .A2(KEYINPUT126), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n905_), .B1(new_n907_), .B2(new_n908_), .ZN(G1351gat));
  NOR2_X1   g708(.A1(new_n417_), .A2(new_n531_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n803_), .A2(new_n910_), .A3(new_n887_), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n911_), .A2(KEYINPUT127), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(KEYINPUT127), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n585_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(G197gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1352gat));
  AOI21_X1  g715(.A(new_n278_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n917_));
  INV_X1    g716(.A(G204gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1353gat));
  OR2_X1    g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n912_), .A2(new_n913_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n587_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(KEYINPUT63), .B(G211gat), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n328_), .B(new_n923_), .C1(new_n912_), .C2(new_n913_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n922_), .A2(new_n924_), .ZN(G1354gat));
  INV_X1    g724(.A(G218gat), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n921_), .A2(new_n926_), .A3(new_n354_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n624_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n928_), .B2(new_n926_), .ZN(G1355gat));
endmodule


