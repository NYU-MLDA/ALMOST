//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n788_, new_n789_, new_n790_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n940_, new_n941_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_;
  NOR2_X1   g000(.A1(G211gat), .A2(G218gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT95), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G211gat), .A2(G218gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n205_), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT95), .B1(new_n207_), .B2(new_n202_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n208_), .A3(KEYINPUT21), .ZN(new_n209_));
  INV_X1    g008(.A(G197gat), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(G204gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT92), .B1(new_n210_), .B2(G204gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n209_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n213_), .ZN(new_n217_));
  AND2_X1   g016(.A1(KEYINPUT93), .A2(KEYINPUT21), .ZN(new_n218_));
  NOR2_X1   g017(.A1(KEYINPUT93), .A2(KEYINPUT21), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n217_), .A2(new_n211_), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G204gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(G197gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n213_), .A2(new_n223_), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n224_), .A2(KEYINPUT21), .B1(new_n203_), .B2(new_n205_), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n221_), .A2(new_n225_), .A3(KEYINPUT94), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT94), .B1(new_n221_), .B2(new_n225_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n216_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT96), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n216_), .B(KEYINPUT96), .C1(new_n226_), .C2(new_n227_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G141gat), .B(G148gat), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT89), .ZN(new_n235_));
  INV_X1    g034(.A(G155gat), .ZN(new_n236_));
  INV_X1    g035(.A(G162gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT89), .B1(G155gat), .B2(G162gat), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G155gat), .A2(G162gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT1), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT1), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(G155gat), .A3(G162gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n234_), .B1(new_n240_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n247_));
  INV_X1    g046(.A(G141gat), .ZN(new_n248_));
  INV_X1    g047(.A(G148gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G141gat), .A2(G148gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT2), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n250_), .A2(new_n253_), .A3(new_n254_), .A4(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n241_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n257_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n246_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT29), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G228gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT91), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n232_), .A2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(G78gat), .B(G106gat), .Z(new_n267_));
  AOI21_X1  g066(.A(new_n263_), .B1(new_n228_), .B2(new_n261_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n266_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n267_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n264_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n271_), .B1(new_n272_), .B2(new_n268_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT97), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n268_), .B1(new_n232_), .B2(new_n265_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n275_), .B1(new_n276_), .B2(new_n267_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n260_), .A2(KEYINPUT29), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(G22gat), .B(G50gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n260_), .A2(KEYINPUT29), .ZN(new_n282_));
  INV_X1    g081(.A(new_n279_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n280_), .A2(new_n281_), .A3(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n281_), .B1(new_n280_), .B2(new_n284_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n274_), .B1(new_n277_), .B2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n285_), .A2(new_n286_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n270_), .A2(new_n289_), .A3(new_n273_), .A4(new_n275_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(G127gat), .A2(G134gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G127gat), .A2(G134gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G120gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G113gat), .ZN(new_n296_));
  INV_X1    g095(.A(G113gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G120gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n296_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n292_), .A2(new_n296_), .A3(new_n298_), .A4(new_n293_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XOR2_X1   g101(.A(KEYINPUT88), .B(G43gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(G71gat), .B(G99gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n304_), .B(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G183gat), .ZN(new_n308_));
  INV_X1    g107(.A(G190gat), .ZN(new_n309_));
  NOR3_X1   g108(.A1(new_n308_), .A2(new_n309_), .A3(KEYINPUT23), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT23), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(G183gat), .B2(G190gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n313_), .A2(KEYINPUT87), .ZN(new_n314_));
  OAI21_X1  g113(.A(KEYINPUT23), .B1(new_n308_), .B2(new_n309_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT87), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n311_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(G183gat), .B2(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G169gat), .A2(G176gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(G169gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT22), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT86), .ZN(new_n324_));
  INV_X1    g123(.A(G176gat), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n322_), .A2(KEYINPUT22), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n324_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n323_), .A2(KEYINPUT86), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n321_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT26), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(KEYINPUT85), .A3(G190gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n308_), .A2(KEYINPUT25), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n309_), .A2(KEYINPUT26), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n331_), .A2(new_n332_), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT84), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(G183gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n330_), .A2(G190gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT85), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n335_), .A2(new_n337_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n334_), .B(new_n340_), .C1(new_n335_), .C2(new_n337_), .ZN(new_n341_));
  OR3_X1    g140(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n342_));
  NOR2_X1   g141(.A1(G169gat), .A2(G176gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n320_), .A2(KEYINPUT24), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n342_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n345_), .B1(new_n311_), .B2(new_n315_), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n319_), .A2(new_n329_), .B1(new_n341_), .B2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT30), .B(G15gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n348_), .B(KEYINPUT31), .Z(new_n349_));
  NOR2_X1   g148(.A1(new_n347_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G227gat), .A2(G233gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n347_), .A2(new_n349_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n352_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n307_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n356_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(new_n354_), .A3(new_n306_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n256_), .A2(new_n258_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n242_), .A2(new_n244_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n238_), .A2(new_n239_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n233_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n302_), .B1(new_n361_), .B2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n301_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n296_), .A2(new_n298_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n368_), .A2(new_n246_), .A3(new_n259_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n365_), .A2(new_n369_), .A3(KEYINPUT4), .ZN(new_n370_));
  NAND2_X1  g169(.A1(G225gat), .A2(G233gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n260_), .A2(new_n373_), .A3(new_n302_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n370_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT99), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT99), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n370_), .A2(new_n377_), .A3(new_n372_), .A4(new_n374_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n365_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n376_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(KEYINPUT100), .B(KEYINPUT0), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G57gat), .B(G85gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n380_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n385_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n376_), .A2(new_n387_), .A3(new_n378_), .A4(new_n379_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n291_), .A2(new_n360_), .A3(new_n389_), .ZN(new_n390_));
  XOR2_X1   g189(.A(G64gat), .B(G92gat), .Z(new_n391_));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n391_), .B(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n347_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT19), .ZN(new_n399_));
  AND4_X1   g198(.A1(new_n338_), .A2(new_n332_), .A3(new_n333_), .A4(new_n337_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(new_n345_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n318_), .A2(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n326_), .A2(new_n323_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(new_n325_), .ZN(new_n404_));
  OAI22_X1  g203(.A1(new_n310_), .A2(new_n313_), .B1(G183gat), .B2(G190gat), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n320_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n402_), .A2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT20), .B1(new_n228_), .B2(new_n407_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n397_), .A2(new_n399_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n399_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n230_), .A2(new_n347_), .A3(new_n231_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT20), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n412_), .B1(new_n228_), .B2(new_n407_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n410_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n396_), .B1(new_n409_), .B2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n411_), .A2(new_n413_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(new_n399_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n347_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n221_), .A2(new_n225_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT94), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n221_), .A2(new_n225_), .A3(KEYINPUT94), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT96), .B1(new_n423_), .B2(new_n216_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n231_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n418_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n408_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n410_), .A3(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n417_), .A2(new_n395_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n415_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT27), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n410_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n411_), .A2(new_n410_), .A3(new_n413_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n396_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(KEYINPUT27), .A3(new_n429_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n432_), .A2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n390_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT104), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n360_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n388_), .A2(KEYINPUT33), .ZN(new_n442_));
  INV_X1    g241(.A(new_n379_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n443_), .B1(new_n375_), .B2(KEYINPUT99), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT33), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n444_), .A2(new_n445_), .A3(new_n387_), .A4(new_n378_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n370_), .A2(new_n371_), .A3(new_n374_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n365_), .A2(new_n369_), .A3(new_n372_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n385_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT101), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n447_), .A2(new_n429_), .A3(new_n415_), .A4(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n395_), .A2(KEYINPUT32), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n455_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n386_), .A2(new_n388_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n417_), .A2(new_n454_), .A3(new_n428_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n453_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT102), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(new_n291_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n288_), .A2(new_n389_), .A3(new_n290_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n432_), .A3(new_n436_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  AOI22_X1  g264(.A1(new_n453_), .A2(new_n459_), .B1(new_n290_), .B2(new_n288_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n466_), .A2(new_n461_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n441_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT103), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n409_), .A2(new_n414_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n431_), .B1(new_n470_), .B2(new_n395_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n435_), .A2(new_n471_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n466_), .A2(new_n461_), .B1(new_n472_), .B2(new_n463_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n460_), .A2(new_n291_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT102), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT103), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(new_n477_), .A3(new_n441_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n440_), .B1(new_n469_), .B2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G183gat), .B(G211gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(G127gat), .B(G155gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  AOI21_X1  g283(.A(KEYINPUT81), .B1(new_n484_), .B2(KEYINPUT17), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G15gat), .B(G22gat), .ZN(new_n486_));
  INV_X1    g285(.A(G1gat), .ZN(new_n487_));
  INV_X1    g286(.A(G8gat), .ZN(new_n488_));
  OAI21_X1  g287(.A(KEYINPUT14), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G8gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n485_), .B(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G231gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT69), .B(G71gat), .ZN(new_n496_));
  INV_X1    g295(.A(G78gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G57gat), .B(G64gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT11), .ZN(new_n500_));
  OR2_X1    g299(.A1(new_n498_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n498_), .A2(KEYINPUT11), .A3(new_n499_), .ZN(new_n502_));
  AND2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n495_), .A2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n504_), .B1(KEYINPUT17), .B2(new_n484_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n495_), .A2(new_n503_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n508_));
  INV_X1    g307(.A(G99gat), .ZN(new_n509_));
  INV_X1    g308(.A(G106gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT6), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n511_), .A2(new_n514_), .A3(new_n515_), .A4(new_n516_), .ZN(new_n517_));
  XOR2_X1   g316(.A(G85gat), .B(G92gat), .Z(new_n518_));
  XNOR2_X1  g317(.A(KEYINPUT67), .B(KEYINPUT8), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT68), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n518_), .ZN(new_n522_));
  AOI22_X1  g321(.A1(new_n520_), .A2(new_n521_), .B1(new_n522_), .B2(KEYINPUT8), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n520_), .A2(new_n521_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT9), .ZN(new_n526_));
  INV_X1    g325(.A(G85gat), .ZN(new_n527_));
  INV_X1    g326(.A(G92gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n526_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT66), .ZN(new_n530_));
  NAND3_X1  g329(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n531_));
  AOI22_X1  g330(.A1(new_n529_), .A2(KEYINPUT65), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n531_), .B1(G85gat), .B2(G92gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT66), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n532_), .B(new_n534_), .C1(KEYINPUT65), .C2(new_n529_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n514_), .A2(new_n515_), .ZN(new_n536_));
  XOR2_X1   g335(.A(KEYINPUT10), .B(G99gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT64), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n535_), .B(new_n536_), .C1(new_n538_), .C2(G106gat), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n525_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G29gat), .B(G36gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G43gat), .B(G50gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(KEYINPUT73), .B(KEYINPUT15), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n543_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n525_), .A2(new_n539_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G232gat), .A2(G233gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n550_), .B(KEYINPUT34), .Z(new_n551_));
  INV_X1    g350(.A(KEYINPUT35), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n551_), .A2(new_n552_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n553_), .B1(new_n554_), .B2(KEYINPUT76), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n555_), .B1(KEYINPUT76), .B2(new_n554_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n544_), .A2(new_n549_), .A3(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(G190gat), .B(G218gat), .Z(new_n558_));
  XNOR2_X1  g357(.A(G134gat), .B(G162gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT36), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n562_), .B(KEYINPUT75), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n546_), .B1(new_n539_), .B2(new_n525_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT74), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n564_), .A2(new_n565_), .B1(new_n540_), .B2(new_n543_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n549_), .A2(KEYINPUT74), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n554_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n557_), .B(new_n563_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT77), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n560_), .B(KEYINPUT36), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n569_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n557_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT78), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n574_), .A2(new_n575_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(KEYINPUT77), .A3(new_n563_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT78), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n580_), .B(new_n573_), .C1(new_n574_), .C2(new_n575_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n572_), .A2(new_n577_), .A3(new_n579_), .A4(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT37), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT37), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n570_), .A2(new_n576_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(KEYINPUT79), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT79), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n583_), .A2(new_n589_), .A3(new_n586_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NOR3_X1   g390(.A1(new_n479_), .A2(new_n507_), .A3(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n548_), .A2(new_n503_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n501_), .A2(new_n502_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n595_), .A2(new_n525_), .A3(new_n539_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n593_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n594_), .A2(KEYINPUT12), .A3(new_n596_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT12), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n548_), .A2(new_n503_), .A3(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n597_), .B1(new_n601_), .B2(new_n593_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G120gat), .B(G148gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(new_n222_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(KEYINPUT5), .B(G176gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n604_), .B(new_n605_), .Z(new_n606_));
  OR2_X1    g405(.A1(new_n606_), .A2(KEYINPUT70), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n602_), .A2(new_n607_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT71), .B(KEYINPUT13), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n610_), .B1(KEYINPUT71), .B2(KEYINPUT13), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n615_), .A2(KEYINPUT72), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(KEYINPUT72), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G113gat), .B(G141gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G169gat), .B(G197gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n492_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(new_n543_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT82), .ZN(new_n624_));
  INV_X1    g423(.A(new_n543_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n492_), .A2(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n624_), .B(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G229gat), .A2(G233gat), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n630_), .A2(KEYINPUT83), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n547_), .A2(new_n492_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n628_), .A3(new_n623_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT83), .ZN(new_n634_));
  AOI22_X1  g433(.A1(new_n627_), .A2(new_n629_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n621_), .B1(new_n631_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n633_), .A2(new_n634_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n630_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n621_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n638_), .B(new_n639_), .C1(KEYINPUT83), .C2(new_n630_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n618_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n592_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n487_), .A3(new_n457_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT38), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n440_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n477_), .B1(new_n476_), .B2(new_n441_), .ZN(new_n650_));
  AOI211_X1 g449(.A(KEYINPUT103), .B(new_n360_), .C1(new_n473_), .C2(new_n475_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n642_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n570_), .A2(new_n576_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT105), .Z(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(new_n507_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G1gat), .B1(new_n658_), .B2(new_n389_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n646_), .A2(new_n647_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n648_), .A2(new_n659_), .A3(new_n660_), .ZN(G1324gat));
  OAI21_X1  g460(.A(G8gat), .B1(new_n658_), .B2(new_n472_), .ZN(new_n662_));
  XOR2_X1   g461(.A(KEYINPUT107), .B(KEYINPUT39), .Z(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n662_), .A2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n472_), .A2(G8gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n645_), .A2(KEYINPUT106), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT106), .ZN(new_n668_));
  INV_X1    g467(.A(new_n666_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n668_), .B1(new_n644_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n667_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n662_), .A2(new_n664_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n665_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n665_), .A2(new_n671_), .A3(KEYINPUT40), .A4(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1325gat));
  OAI21_X1  g476(.A(G15gat), .B1(new_n658_), .B2(new_n441_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n678_), .A2(KEYINPUT41), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(KEYINPUT41), .ZN(new_n680_));
  OR3_X1    g479(.A1(new_n644_), .A2(G15gat), .A3(new_n441_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n679_), .A2(new_n680_), .A3(new_n681_), .ZN(G1326gat));
  OAI21_X1  g481(.A(G22gat), .B1(new_n658_), .B2(new_n291_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT42), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n291_), .A2(G22gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n644_), .B2(new_n685_), .ZN(G1327gat));
  INV_X1    g485(.A(new_n507_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n687_), .A2(new_n655_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n654_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(G29gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n690_), .A3(new_n457_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT108), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n692_), .B1(new_n591_), .B2(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n589_), .B1(new_n583_), .B2(new_n586_), .ZN(new_n695_));
  AOI211_X1 g494(.A(KEYINPUT79), .B(new_n585_), .C1(new_n582_), .C2(KEYINPUT37), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n694_), .B1(new_n479_), .B2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n693_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT43), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n652_), .A2(new_n591_), .A3(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n698_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n653_), .A2(new_n507_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT44), .B1(new_n702_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706_));
  AOI211_X1 g505(.A(new_n706_), .B(new_n703_), .C1(new_n698_), .C2(new_n701_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n705_), .A2(new_n707_), .A3(new_n389_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n691_), .B1(new_n708_), .B2(new_n690_), .ZN(G1328gat));
  INV_X1    g508(.A(KEYINPUT46), .ZN(new_n710_));
  INV_X1    g509(.A(G36gat), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n705_), .A2(new_n707_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n712_), .B2(new_n437_), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n654_), .A2(new_n711_), .A3(new_n437_), .A4(new_n688_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT45), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n710_), .B1(new_n713_), .B2(new_n716_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n705_), .A2(new_n707_), .A3(new_n472_), .ZN(new_n718_));
  OAI211_X1 g517(.A(KEYINPUT46), .B(new_n715_), .C1(new_n718_), .C2(new_n711_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1329gat));
  INV_X1    g519(.A(new_n705_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n702_), .A2(KEYINPUT44), .A3(new_n704_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n721_), .A2(G43gat), .A3(new_n360_), .A4(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n654_), .A2(new_n360_), .A3(new_n688_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n725_));
  INV_X1    g524(.A(G43gat), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n725_), .B1(new_n724_), .B2(new_n726_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n723_), .A2(new_n729_), .A3(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n723_), .B2(new_n729_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(G1330gat));
  INV_X1    g532(.A(G50gat), .ZN(new_n734_));
  INV_X1    g533(.A(new_n291_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n689_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n705_), .A2(new_n707_), .A3(new_n291_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n737_), .B2(new_n734_), .ZN(G1331gat));
  INV_X1    g537(.A(new_n618_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n739_), .A2(new_n479_), .A3(new_n641_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n657_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT112), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n740_), .A2(KEYINPUT112), .A3(new_n657_), .ZN(new_n744_));
  INV_X1    g543(.A(G57gat), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n389_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n743_), .A2(new_n744_), .A3(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT113), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n747_), .A2(new_n748_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n615_), .A2(new_n641_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n592_), .A2(new_n751_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n752_), .A2(KEYINPUT111), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n389_), .B1(new_n752_), .B2(KEYINPUT111), .ZN(new_n754_));
  AOI21_X1  g553(.A(G57gat), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n749_), .A2(new_n750_), .A3(new_n755_), .ZN(G1332gat));
  OR3_X1    g555(.A1(new_n752_), .A2(G64gat), .A3(new_n472_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n743_), .A2(new_n437_), .A3(new_n744_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT48), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(G64gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(G64gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(G1333gat));
  OR3_X1    g561(.A1(new_n752_), .A2(G71gat), .A3(new_n441_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n743_), .A2(new_n360_), .A3(new_n744_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT49), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n764_), .A2(new_n765_), .A3(G71gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n764_), .B2(G71gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(G1334gat));
  NAND3_X1  g567(.A1(new_n743_), .A2(new_n735_), .A3(new_n744_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n769_), .A2(new_n770_), .A3(G78gat), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n769_), .B2(G78gat), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n735_), .A2(new_n497_), .ZN(new_n773_));
  OAI22_X1  g572(.A1(new_n771_), .A2(new_n772_), .B1(new_n752_), .B2(new_n773_), .ZN(G1335gat));
  NAND2_X1  g573(.A1(new_n740_), .A2(new_n688_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n527_), .B1(new_n775_), .B2(new_n389_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT114), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n751_), .A2(new_n507_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n698_), .B2(new_n701_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n780_), .A2(G85gat), .A3(new_n457_), .ZN(new_n781_));
  OAI211_X1 g580(.A(KEYINPUT114), .B(new_n527_), .C1(new_n775_), .C2(new_n389_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n778_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n778_), .A2(KEYINPUT115), .A3(new_n781_), .A4(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1336gat));
  INV_X1    g586(.A(new_n775_), .ZN(new_n788_));
  AOI21_X1  g587(.A(G92gat), .B1(new_n788_), .B2(new_n437_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n472_), .A2(new_n528_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n780_), .B2(new_n790_), .ZN(G1337gat));
  NOR3_X1   g590(.A1(new_n775_), .A2(new_n441_), .A3(new_n538_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n509_), .B1(new_n780_), .B2(new_n360_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT51), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n794_), .B(new_n796_), .ZN(G1338gat));
  NAND3_X1  g596(.A1(new_n788_), .A2(new_n510_), .A3(new_n735_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT52), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n780_), .A2(new_n735_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(G106gat), .ZN(new_n801_));
  AOI211_X1 g600(.A(KEYINPUT52), .B(new_n510_), .C1(new_n780_), .C2(new_n735_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n798_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT53), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n805_), .B(new_n798_), .C1(new_n801_), .C2(new_n802_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(G1339gat));
  AND2_X1   g606(.A1(new_n602_), .A2(new_n606_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n636_), .B2(new_n640_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n810_), .B1(new_n601_), .B2(new_n593_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n593_), .ZN(new_n812_));
  AOI211_X1 g611(.A(KEYINPUT55), .B(new_n812_), .C1(new_n598_), .C2(new_n600_), .ZN(new_n813_));
  OAI22_X1  g612(.A1(new_n811_), .A2(new_n813_), .B1(new_n593_), .B2(new_n601_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n606_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n814_), .A2(KEYINPUT117), .A3(KEYINPUT56), .A4(new_n815_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n809_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT56), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n601_), .A2(new_n593_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n601_), .A2(new_n593_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT55), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n601_), .A2(new_n810_), .A3(new_n593_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n819_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n818_), .B1(new_n823_), .B2(new_n606_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n814_), .A2(KEYINPUT56), .A3(new_n815_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n817_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n627_), .A2(new_n628_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n632_), .A2(new_n629_), .A3(new_n623_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n829_), .A2(new_n621_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n640_), .A2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n611_), .A2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT57), .B(new_n655_), .C1(new_n828_), .C2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n833_), .B1(new_n817_), .B2(new_n827_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n655_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n835_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n832_), .A2(new_n808_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n826_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT56), .B1(new_n814_), .B2(new_n815_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n839_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT58), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n839_), .B(KEYINPUT58), .C1(new_n840_), .C2(new_n841_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n844_), .B(new_n845_), .C1(new_n695_), .C2(new_n696_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n834_), .A2(new_n838_), .A3(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n507_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n641_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n588_), .A2(new_n590_), .A3(new_n849_), .A4(new_n687_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT54), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n697_), .A2(new_n852_), .A3(new_n687_), .A4(new_n849_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n848_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n472_), .A2(new_n457_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n441_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n855_), .A2(new_n291_), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(G113gat), .B1(new_n859_), .B2(new_n641_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n735_), .B1(new_n848_), .B2(new_n854_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n857_), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(KEYINPUT118), .A2(KEYINPUT59), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n863_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n861_), .B2(new_n857_), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT119), .B1(new_n865_), .B2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n858_), .A2(new_n867_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n871_), .A2(new_n872_), .A3(new_n864_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n642_), .A2(new_n297_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n860_), .B1(new_n874_), .B2(new_n875_), .ZN(G1340gat));
  OAI21_X1  g675(.A(new_n295_), .B1(new_n615_), .B2(KEYINPUT60), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n859_), .B(new_n877_), .C1(KEYINPUT60), .C2(new_n295_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n739_), .B1(new_n871_), .B2(new_n864_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880_));
  OAI21_X1  g679(.A(G120gat), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n880_), .B(new_n618_), .C1(new_n865_), .C2(new_n869_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n878_), .B1(new_n881_), .B2(new_n883_), .ZN(G1341gat));
  NAND2_X1  g683(.A1(new_n687_), .A2(G127gat), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(KEYINPUT122), .ZN(new_n886_));
  INV_X1    g685(.A(G127gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n858_), .B2(new_n507_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT121), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n889_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n874_), .A2(new_n886_), .B1(new_n890_), .B2(new_n891_), .ZN(G1342gat));
  AOI21_X1  g691(.A(G134gat), .B1(new_n859_), .B2(new_n656_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n591_), .A2(G134gat), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n874_), .B2(new_n894_), .ZN(G1343gat));
  AOI21_X1  g694(.A(new_n360_), .B1(new_n848_), .B2(new_n854_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n856_), .A2(new_n291_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n642_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(new_n248_), .ZN(G1344gat));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n739_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(new_n249_), .ZN(G1345gat));
  NOR2_X1   g701(.A1(new_n898_), .A2(new_n507_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT61), .B(G155gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906_));
  INV_X1    g705(.A(new_n898_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n656_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n906_), .B1(new_n908_), .B2(new_n237_), .ZN(new_n909_));
  AOI211_X1 g708(.A(KEYINPUT123), .B(G162gat), .C1(new_n907_), .C2(new_n656_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n898_), .A2(new_n237_), .A3(new_n697_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n909_), .A2(new_n910_), .A3(new_n911_), .ZN(G1347gat));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n855_), .A2(new_n291_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n437_), .A2(new_n360_), .A3(new_n389_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT124), .ZN(new_n916_));
  OR2_X1    g715(.A1(new_n914_), .A2(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n642_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n913_), .B1(new_n918_), .B2(new_n322_), .ZN(new_n919_));
  OAI211_X1 g718(.A(KEYINPUT62), .B(G169gat), .C1(new_n917_), .C2(new_n642_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n403_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n919_), .A2(new_n920_), .A3(new_n921_), .ZN(G1348gat));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n916_), .B1(new_n914_), .B2(new_n923_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n861_), .A2(KEYINPUT125), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n739_), .A2(new_n325_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n924_), .A2(new_n925_), .A3(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n927_), .A2(new_n928_), .ZN(new_n929_));
  NAND4_X1  g728(.A1(new_n924_), .A2(KEYINPUT126), .A3(new_n925_), .A4(new_n926_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n325_), .B1(new_n917_), .B2(new_n615_), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n929_), .A2(new_n930_), .A3(new_n931_), .ZN(G1349gat));
  NAND3_X1  g731(.A1(new_n924_), .A2(new_n687_), .A3(new_n925_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n917_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n507_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n935_));
  AOI22_X1  g734(.A1(new_n933_), .A2(new_n308_), .B1(new_n934_), .B2(new_n935_), .ZN(G1350gat));
  OAI21_X1  g735(.A(G190gat), .B1(new_n917_), .B2(new_n697_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n656_), .A2(new_n338_), .A3(new_n333_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n917_), .B2(new_n938_), .ZN(G1351gat));
  AND3_X1   g738(.A1(new_n896_), .A2(new_n463_), .A3(new_n437_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n641_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n618_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g743(.A(new_n507_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n940_), .A2(new_n945_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n947_));
  XOR2_X1   g746(.A(new_n946_), .B(new_n947_), .Z(G1354gat));
  NAND2_X1  g747(.A1(new_n940_), .A2(new_n656_), .ZN(new_n949_));
  XOR2_X1   g748(.A(KEYINPUT127), .B(G218gat), .Z(new_n950_));
  NOR2_X1   g749(.A1(new_n697_), .A2(new_n950_), .ZN(new_n951_));
  AOI22_X1  g750(.A1(new_n949_), .A2(new_n950_), .B1(new_n940_), .B2(new_n951_), .ZN(G1355gat));
endmodule


