//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n957_, new_n958_, new_n959_,
    new_n961_, new_n962_, new_n964_, new_n965_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n980_, new_n981_;
  XOR2_X1   g000(.A(G211gat), .B(G218gat), .Z(new_n202_));
  NOR2_X1   g001(.A1(G197gat), .A2(G204gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205_));
  NAND4_X1  g004(.A1(new_n202_), .A2(KEYINPUT21), .A3(new_n204_), .A4(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(KEYINPUT21), .A3(new_n205_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208_));
  AND2_X1   g007(.A1(G197gat), .A2(G204gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(new_n209_), .B2(new_n203_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n206_), .A2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT3), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(KEYINPUT2), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n218_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(G155gat), .B2(G162gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT85), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n224_), .A2(new_n225_), .A3(new_n219_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n225_), .B1(new_n224_), .B2(new_n219_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n219_), .A2(KEYINPUT1), .ZN(new_n228_));
  NOR3_X1   g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT84), .B1(G141gat), .B2(G148gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NOR3_X1   g030(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n216_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(KEYINPUT86), .B1(new_n229_), .B2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n219_), .B1(new_n220_), .B2(KEYINPUT1), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(KEYINPUT85), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n224_), .A2(new_n225_), .A3(new_n219_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n228_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT86), .ZN(new_n240_));
  INV_X1    g039(.A(new_n233_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n222_), .B1(new_n234_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT29), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n213_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G228gat), .A2(G233gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n246_), .B(KEYINPUT89), .Z(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  AND2_X1   g048(.A1(new_n206_), .A2(new_n212_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n218_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n228_), .B1(new_n235_), .B2(KEYINPUT85), .ZN(new_n252_));
  AOI211_X1 g051(.A(KEYINPUT86), .B(new_n233_), .C1(new_n252_), .C2(new_n237_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n240_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n251_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n250_), .B1(new_n255_), .B2(KEYINPUT29), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n247_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G78gat), .B(G106gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n249_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT90), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND4_X1  g060(.A1(new_n249_), .A2(new_n257_), .A3(KEYINPUT90), .A4(new_n258_), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n244_), .B(new_n251_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n263_));
  XOR2_X1   g062(.A(KEYINPUT87), .B(KEYINPUT28), .Z(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n234_), .A2(new_n242_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n264_), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n266_), .A2(new_n244_), .A3(new_n251_), .A4(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G22gat), .B(G50gat), .Z(new_n269_));
  AND3_X1   g068(.A1(new_n265_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n258_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n256_), .A2(new_n247_), .ZN(new_n274_));
  AOI211_X1 g073(.A(new_n250_), .B(new_n248_), .C1(new_n255_), .C2(KEYINPUT29), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n261_), .A2(new_n262_), .A3(new_n272_), .A4(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT88), .B1(new_n270_), .B2(new_n271_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n265_), .A2(new_n268_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n269_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT88), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n265_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n274_), .A2(new_n275_), .A3(new_n273_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n258_), .B1(new_n249_), .B2(new_n257_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n278_), .B(new_n284_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT27), .ZN(new_n288_));
  INV_X1    g087(.A(G169gat), .ZN(new_n289_));
  INV_X1    g088(.A(G176gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(KEYINPUT24), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G183gat), .A2(G190gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT23), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT23), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(G183gat), .A3(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT24), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n293_), .A2(new_n298_), .A3(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(KEYINPUT79), .A2(KEYINPUT26), .ZN(new_n303_));
  NOR2_X1   g102(.A1(KEYINPUT79), .A2(KEYINPUT26), .ZN(new_n304_));
  OAI21_X1  g103(.A(G190gat), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT80), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  OAI211_X1 g106(.A(KEYINPUT80), .B(G190gat), .C1(new_n303_), .C2(new_n304_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G190gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT26), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT25), .ZN(new_n312_));
  OR2_X1    g111(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(KEYINPUT78), .A2(G183gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n312_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n311_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n302_), .B1(new_n309_), .B2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n295_), .A2(new_n297_), .A3(KEYINPUT81), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT81), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n294_), .A2(new_n324_), .A3(KEYINPUT23), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n313_), .A2(new_n314_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n327_), .A2(G190gat), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n322_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n318_), .A2(new_n250_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT20), .ZN(new_n331_));
  OR2_X1    g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n296_), .B1(G183gat), .B2(G190gat), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n294_), .A2(KEYINPUT23), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n322_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(KEYINPUT91), .A2(KEYINPUT24), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(KEYINPUT91), .A2(KEYINPUT24), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n291_), .B(new_n292_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT26), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G190gat), .ZN(new_n342_));
  AND2_X1   g141(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n311_), .B(new_n342_), .C1(new_n343_), .C2(new_n316_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n339_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n345_), .A2(new_n299_), .A3(new_n337_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n340_), .A2(new_n344_), .A3(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n336_), .B1(new_n347_), .B2(new_n326_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n331_), .B1(new_n348_), .B2(new_n213_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n330_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT92), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G226gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT19), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n350_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT20), .B1(new_n348_), .B2(new_n213_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n318_), .A2(new_n329_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n213_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n353_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n356_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n354_), .A2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G8gat), .B(G36gat), .Z(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G64gat), .B(G92gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n359_), .B1(new_n330_), .B2(new_n349_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n368_), .A2(new_n351_), .ZN(new_n369_));
  NOR3_X1   g168(.A1(new_n361_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n250_), .B1(new_n318_), .B2(new_n329_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n371_), .A2(new_n355_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n351_), .A2(new_n368_), .B1(new_n372_), .B2(new_n359_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n350_), .A2(new_n353_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT92), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n366_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n288_), .B1(new_n370_), .B2(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n359_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n350_), .A2(new_n353_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n367_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(KEYINPUT100), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n373_), .A2(new_n366_), .A3(new_n375_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT100), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n383_), .B(new_n367_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n381_), .A2(KEYINPUT27), .A3(new_n382_), .A4(new_n384_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n277_), .A2(new_n287_), .A3(new_n377_), .A4(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387_));
  INV_X1    g186(.A(G15gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT30), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n357_), .B(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(G134gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G127gat), .ZN(new_n393_));
  INV_X1    g192(.A(G127gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(G134gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G120gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(G113gat), .ZN(new_n398_));
  INV_X1    g197(.A(G113gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(G120gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  AOI22_X1  g202(.A1(new_n393_), .A2(new_n395_), .B1(new_n398_), .B2(new_n400_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT82), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n404_), .A2(new_n405_), .A3(KEYINPUT83), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT83), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n396_), .A2(new_n401_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(new_n408_), .B2(KEYINPUT82), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n403_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT83), .B1(new_n404_), .B2(new_n405_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n408_), .A2(KEYINPUT82), .A3(new_n407_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(new_n402_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n391_), .B(new_n414_), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G71gat), .B(G99gat), .ZN(new_n416_));
  INV_X1    g215(.A(G43gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(KEYINPUT31), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n415_), .B(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n403_), .A2(new_n408_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n251_), .B(new_n422_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n423_), .B(KEYINPUT4), .C1(new_n243_), .C2(new_n414_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n414_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n255_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n428_), .B(KEYINPUT94), .Z(new_n429_));
  NAND3_X1  g228(.A1(new_n424_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  OAI211_X1 g229(.A(new_n423_), .B(new_n428_), .C1(new_n243_), .C2(new_n414_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT96), .ZN(new_n433_));
  XOR2_X1   g232(.A(G1gat), .B(G29gat), .Z(new_n434_));
  XOR2_X1   g233(.A(new_n433_), .B(new_n434_), .Z(new_n435_));
  XNOR2_X1  g234(.A(G57gat), .B(G85gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n433_), .B(new_n434_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n436_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n437_), .A2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n430_), .A2(new_n431_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n442_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n421_), .A2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n386_), .A2(new_n446_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n430_), .A2(new_n431_), .A3(new_n442_), .ZN(new_n448_));
  XOR2_X1   g247(.A(KEYINPUT98), .B(KEYINPUT33), .Z(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT99), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n437_), .A2(new_n440_), .A3(KEYINPUT33), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n430_), .A2(new_n431_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT97), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT97), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n430_), .A2(new_n453_), .A3(new_n456_), .A4(new_n431_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n424_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n459_));
  OAI211_X1 g258(.A(new_n423_), .B(new_n429_), .C1(new_n243_), .C2(new_n414_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n441_), .A3(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n367_), .B1(new_n361_), .B2(new_n369_), .ZN(new_n462_));
  AND3_X1   g261(.A1(new_n461_), .A2(new_n462_), .A3(new_n382_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n448_), .A2(KEYINPUT99), .A3(new_n449_), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n452_), .A2(new_n458_), .A3(new_n463_), .A4(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n277_), .A2(new_n287_), .ZN(new_n466_));
  OAI211_X1 g265(.A(KEYINPUT32), .B(new_n366_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n366_), .A2(KEYINPUT32), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n373_), .A2(new_n375_), .A3(new_n468_), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n467_), .B(new_n469_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n465_), .A2(new_n466_), .A3(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n445_), .A2(new_n377_), .A3(new_n385_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n277_), .A2(new_n287_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n421_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n447_), .B1(new_n471_), .B2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G29gat), .B(G36gat), .Z(new_n476_));
  XOR2_X1   g275(.A(G43gat), .B(G50gat), .Z(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G29gat), .B(G36gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G43gat), .B(G50gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  AND3_X1   g280(.A1(new_n478_), .A2(KEYINPUT15), .A3(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(KEYINPUT15), .B1(new_n478_), .B2(new_n481_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G15gat), .B(G22gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G1gat), .A2(G8gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT14), .ZN(new_n487_));
  INV_X1    g286(.A(G1gat), .ZN(new_n488_));
  INV_X1    g287(.A(G8gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  AOI22_X1  g289(.A1(new_n485_), .A2(new_n487_), .B1(new_n486_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n485_), .A2(new_n486_), .A3(new_n490_), .A4(new_n487_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n484_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n478_), .A2(new_n481_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G229gat), .A2(G233gat), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NOR3_X1   g299(.A1(new_n495_), .A2(new_n498_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT75), .ZN(new_n502_));
  INV_X1    g301(.A(new_n493_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n481_), .B(new_n478_), .C1(new_n503_), .C2(new_n491_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n504_), .A2(new_n497_), .A3(KEYINPUT74), .ZN(new_n505_));
  AOI21_X1  g304(.A(KEYINPUT74), .B1(new_n504_), .B2(new_n497_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n502_), .B1(new_n507_), .B2(new_n499_), .ZN(new_n508_));
  OAI211_X1 g307(.A(KEYINPUT75), .B(new_n500_), .C1(new_n505_), .C2(new_n506_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n501_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G113gat), .B(G141gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G169gat), .B(G197gat), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n511_), .B(new_n512_), .Z(new_n513_));
  OR2_X1    g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT76), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n510_), .A2(new_n515_), .A3(new_n513_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n510_), .B2(new_n513_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n514_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT77), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OAI211_X1 g319(.A(KEYINPUT77), .B(new_n514_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n475_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G85gat), .A2(G92gat), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(G85gat), .A2(G92gat), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G99gat), .A2(G106gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT6), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT6), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n531_), .A2(G99gat), .A3(G106gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  OR3_X1    g333(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n528_), .B1(new_n534_), .B2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT8), .B1(new_n528_), .B2(KEYINPUT65), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  OAI221_X1 g339(.A(new_n528_), .B1(KEYINPUT65), .B2(KEYINPUT8), .C1(new_n534_), .C2(new_n537_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n542_));
  NOR2_X1   g341(.A1(KEYINPUT9), .A2(G92gat), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n542_), .B1(new_n528_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(G85gat), .ZN(new_n545_));
  INV_X1    g344(.A(G92gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n543_), .B1(new_n547_), .B2(new_n525_), .ZN(new_n548_));
  XOR2_X1   g347(.A(KEYINPUT64), .B(KEYINPUT9), .Z(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n551_));
  NOR2_X1   g350(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(G106gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n544_), .A2(new_n550_), .A3(new_n533_), .A4(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n540_), .A2(new_n541_), .A3(new_n556_), .A4(new_n496_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT69), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n540_), .A2(new_n541_), .A3(new_n556_), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n557_), .A2(new_n558_), .B1(new_n559_), .B2(new_n484_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT70), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n548_), .A2(new_n549_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT10), .B(G99gat), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n533_), .B1(new_n563_), .B2(G106gat), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n565_), .A2(new_n550_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n566_), .A2(KEYINPUT69), .A3(new_n496_), .A4(new_n541_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n560_), .A2(new_n561_), .A3(new_n567_), .A4(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n557_), .A2(new_n558_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n559_), .A2(new_n484_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n567_), .A2(new_n573_), .A3(new_n561_), .A4(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n570_), .ZN(new_n576_));
  AOI21_X1  g375(.A(KEYINPUT35), .B1(new_n560_), .B2(new_n567_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n572_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT71), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G190gat), .B(G218gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n578_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n584_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n580_), .A2(new_n586_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n587_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n578_), .B(new_n579_), .C1(new_n589_), .C2(new_n585_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(KEYINPUT72), .B(KEYINPUT37), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n588_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(G57gat), .B(G64gat), .Z(new_n597_));
  INV_X1    g396(.A(KEYINPUT11), .ZN(new_n598_));
  INV_X1    g397(.A(G71gat), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(G78gat), .ZN(new_n600_));
  INV_X1    g399(.A(G78gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(G71gat), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n597_), .A2(new_n598_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(KEYINPUT66), .B1(new_n597_), .B2(new_n598_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G57gat), .B(G64gat), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT66), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n605_), .A2(new_n606_), .A3(KEYINPUT11), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(new_n604_), .A3(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n600_), .A2(new_n602_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n609_), .B1(new_n605_), .B2(KEYINPUT11), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n605_), .A2(new_n606_), .A3(KEYINPUT11), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n606_), .B1(new_n605_), .B2(KEYINPUT11), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n610_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n608_), .A2(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n566_), .A2(new_n541_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G230gat), .A2(G233gat), .ZN(new_n616_));
  AOI21_X1  g415(.A(KEYINPUT68), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(KEYINPUT68), .A3(new_n616_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  AND2_X1   g419(.A1(new_n608_), .A2(new_n613_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n621_), .A2(new_n559_), .A3(KEYINPUT12), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(KEYINPUT12), .B1(new_n621_), .B2(new_n559_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n620_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n621_), .A2(new_n559_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT67), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n615_), .A2(KEYINPUT67), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n621_), .A2(new_n559_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n629_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n616_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n626_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G120gat), .B(G148gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT5), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n637_), .B(new_n638_), .Z(new_n639_));
  NAND2_X1  g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n639_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n626_), .A2(new_n634_), .A3(new_n641_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n640_), .A2(KEYINPUT13), .A3(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT13), .B1(new_n640_), .B2(new_n642_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT73), .Z(new_n647_));
  XNOR2_X1  g446(.A(new_n494_), .B(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(new_n614_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT17), .ZN(new_n650_));
  XNOR2_X1  g449(.A(G127gat), .B(G155gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT16), .ZN(new_n652_));
  XOR2_X1   g451(.A(G183gat), .B(G211gat), .Z(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n649_), .A2(new_n650_), .A3(new_n654_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(KEYINPUT17), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n649_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n655_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n596_), .A2(new_n645_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n524_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n445_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(new_n488_), .A3(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT38), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n386_), .A2(new_n446_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n470_), .A2(new_n277_), .A3(new_n287_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n452_), .A2(new_n463_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n458_), .A2(new_n464_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n667_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n472_), .A2(new_n473_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n421_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n666_), .B1(new_n670_), .B2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n591_), .B(KEYINPUT102), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT103), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT101), .ZN(new_n678_));
  INV_X1    g477(.A(new_n645_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n523_), .B2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n522_), .A2(new_n645_), .A3(KEYINPUT101), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n677_), .A2(new_n658_), .A3(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(G1gat), .B1(new_n683_), .B2(new_n445_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n665_), .A2(new_n684_), .ZN(G1324gat));
  AND2_X1   g484(.A1(new_n377_), .A2(new_n385_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n683_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT104), .B1(new_n688_), .B2(G8gat), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT104), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n687_), .A2(new_n690_), .A3(new_n489_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT39), .ZN(new_n692_));
  OR3_X1    g491(.A1(new_n689_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n689_), .A2(new_n692_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n686_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n662_), .A2(new_n489_), .A3(new_n695_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n693_), .A2(KEYINPUT40), .A3(new_n694_), .A4(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT40), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n694_), .A2(new_n696_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n689_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n697_), .A2(new_n701_), .ZN(G1325gat));
  OAI21_X1  g501(.A(G15gat), .B1(new_n683_), .B2(new_n672_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT41), .Z(new_n704_));
  NAND3_X1  g503(.A1(new_n662_), .A2(new_n388_), .A3(new_n421_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1326gat));
  OAI21_X1  g505(.A(G22gat), .B1(new_n683_), .B2(new_n466_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT42), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n466_), .A2(G22gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n661_), .B2(new_n709_), .ZN(G1327gat));
  INV_X1    g509(.A(new_n591_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n711_), .A2(new_n658_), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n524_), .A2(new_n645_), .A3(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G29gat), .B1(new_n713_), .B2(new_n663_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n658_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n680_), .A2(new_n715_), .A3(new_n681_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n471_), .A2(new_n474_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n596_), .B1(new_n718_), .B2(new_n666_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT105), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n722_));
  OAI211_X1 g521(.A(new_n722_), .B(KEYINPUT43), .C1(new_n475_), .C2(new_n596_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n725_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n726_));
  NOR4_X1   g525(.A1(new_n475_), .A2(KEYINPUT106), .A3(new_n596_), .A4(KEYINPUT43), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT44), .B(new_n717_), .C1(new_n724_), .C2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT107), .ZN(new_n730_));
  INV_X1    g529(.A(new_n596_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n674_), .A2(new_n720_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(KEYINPUT106), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n719_), .A2(new_n725_), .A3(new_n720_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n721_), .A2(new_n723_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n716_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n737_), .A2(new_n738_), .A3(KEYINPUT44), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n717_), .B1(new_n724_), .B2(new_n728_), .ZN(new_n741_));
  AOI22_X1  g540(.A1(new_n730_), .A2(new_n739_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n663_), .A2(G29gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n714_), .B1(new_n742_), .B2(new_n743_), .ZN(G1328gat));
  INV_X1    g543(.A(G36gat), .ZN(new_n745_));
  OR2_X1    g544(.A1(new_n686_), .A2(KEYINPUT109), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n686_), .A2(KEYINPUT109), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n713_), .A2(new_n745_), .A3(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT110), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT45), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n695_), .B1(new_n737_), .B2(KEYINPUT44), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n730_), .B2(new_n739_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n753_), .A2(new_n754_), .A3(new_n745_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n686_), .B1(new_n741_), .B2(new_n740_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n738_), .B1(new_n737_), .B2(KEYINPUT44), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n733_), .A2(new_n734_), .B1(new_n721_), .B2(new_n723_), .ZN(new_n758_));
  NOR4_X1   g557(.A1(new_n758_), .A2(KEYINPUT107), .A3(new_n740_), .A4(new_n716_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n756_), .B1(new_n757_), .B2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT108), .B1(new_n760_), .B2(G36gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n751_), .B1(new_n755_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(KEYINPUT46), .B(new_n751_), .C1(new_n755_), .C2(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1329gat));
  NAND3_X1  g565(.A1(new_n742_), .A2(G43gat), .A3(new_n421_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n713_), .A2(new_n421_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(G43gat), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g569(.A(G50gat), .B1(new_n713_), .B2(new_n473_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n473_), .A2(G50gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n742_), .B2(new_n772_), .ZN(G1331gat));
  AND4_X1   g572(.A1(new_n677_), .A2(new_n658_), .A3(new_n523_), .A4(new_n679_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n774_), .A2(G57gat), .A3(new_n663_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT112), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n674_), .A2(new_n523_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT111), .ZN(new_n778_));
  NOR4_X1   g577(.A1(new_n778_), .A2(new_n715_), .A3(new_n645_), .A4(new_n731_), .ZN(new_n779_));
  AOI21_X1  g578(.A(G57gat), .B1(new_n779_), .B2(new_n663_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n776_), .A2(new_n780_), .ZN(G1332gat));
  INV_X1    g580(.A(G64gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n774_), .B2(new_n748_), .ZN(new_n783_));
  XOR2_X1   g582(.A(new_n783_), .B(KEYINPUT48), .Z(new_n784_));
  NAND3_X1  g583(.A1(new_n779_), .A2(new_n782_), .A3(new_n748_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(G1333gat));
  AOI21_X1  g585(.A(new_n599_), .B1(new_n774_), .B2(new_n421_), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT49), .Z(new_n788_));
  NAND3_X1  g587(.A1(new_n779_), .A2(new_n599_), .A3(new_n421_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1334gat));
  AOI21_X1  g589(.A(new_n601_), .B1(new_n774_), .B2(new_n473_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT50), .Z(new_n792_));
  NAND3_X1  g591(.A1(new_n779_), .A2(new_n601_), .A3(new_n473_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(G1335gat));
  NOR4_X1   g593(.A1(new_n758_), .A2(new_n658_), .A3(new_n522_), .A4(new_n645_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(G85gat), .B1(new_n797_), .B2(new_n445_), .ZN(new_n798_));
  NOR4_X1   g597(.A1(new_n778_), .A2(new_n711_), .A3(new_n658_), .A4(new_n645_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n799_), .A2(new_n545_), .A3(new_n663_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1336gat));
  INV_X1    g600(.A(new_n748_), .ZN(new_n802_));
  OAI21_X1  g601(.A(G92gat), .B1(new_n797_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n799_), .A2(new_n546_), .A3(new_n695_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(G1337gat));
  INV_X1    g604(.A(G99gat), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n795_), .B(KEYINPUT113), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n421_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n799_), .A2(new_n421_), .A3(new_n553_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT51), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(G99gat), .B1(new_n797_), .B2(new_n672_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT51), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n813_), .A3(new_n809_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n811_), .A2(new_n814_), .ZN(G1338gat));
  NAND3_X1  g614(.A1(new_n799_), .A2(new_n554_), .A3(new_n473_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n554_), .B1(new_n795_), .B2(new_n473_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n817_), .A2(new_n818_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n816_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT53), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n823_), .B(new_n816_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(G1339gat));
  NOR3_X1   g624(.A1(new_n386_), .A2(new_n672_), .A3(new_n445_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  OR2_X1    g626(.A1(new_n516_), .A2(new_n517_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n513_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n497_), .A2(new_n500_), .ZN(new_n830_));
  OAI221_X1 g629(.A(new_n829_), .B1(new_n495_), .B2(new_n830_), .C1(new_n507_), .C2(new_n500_), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n828_), .A2(new_n642_), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT12), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n631_), .A2(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n629_), .A2(new_n630_), .A3(new_n834_), .A4(new_n622_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n633_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT116), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n835_), .A2(new_n838_), .A3(new_n633_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n837_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n626_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n619_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n625_), .B(KEYINPUT55), .C1(new_n844_), .C2(new_n617_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n620_), .A2(KEYINPUT117), .A3(KEYINPUT55), .A4(new_n625_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n639_), .B1(new_n843_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT56), .ZN(new_n851_));
  INV_X1    g650(.A(new_n849_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n837_), .A2(new_n839_), .B1(new_n626_), .B2(new_n841_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n641_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT56), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n832_), .A2(new_n851_), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(KEYINPUT119), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(KEYINPUT119), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n832_), .A2(new_n851_), .A3(new_n856_), .A4(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(new_n731_), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863_));
  INV_X1    g662(.A(new_n642_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n864_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n855_), .B1(new_n854_), .B2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n850_), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n865_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n640_), .A2(new_n642_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n828_), .A2(new_n870_), .A3(new_n831_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n863_), .B1(new_n872_), .B2(new_n711_), .ZN(new_n873_));
  AOI211_X1 g672(.A(KEYINPUT57), .B(new_n591_), .C1(new_n869_), .C2(new_n871_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n862_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT120), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n862_), .B(new_n877_), .C1(new_n873_), .C2(new_n874_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n876_), .A2(new_n715_), .A3(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n659_), .A2(new_n522_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT114), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT114), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n880_), .A2(new_n884_), .A3(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT115), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n888_));
  OAI211_X1 g687(.A(KEYINPUT115), .B(KEYINPUT54), .C1(new_n659_), .C2(new_n522_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n886_), .A2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n827_), .B1(new_n879_), .B2(new_n891_), .ZN(new_n892_));
  AOI21_X1  g691(.A(G113gat), .B1(new_n892_), .B2(new_n522_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n875_), .A2(new_n715_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n891_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n895_), .A2(new_n896_), .A3(new_n826_), .ZN(new_n897_));
  OAI211_X1 g696(.A(KEYINPUT121), .B(new_n897_), .C1(new_n892_), .C2(new_n896_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n883_), .A2(new_n885_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n658_), .B1(new_n875_), .B2(KEYINPUT120), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n878_), .ZN(new_n902_));
  OAI21_X1  g701(.A(KEYINPUT59), .B1(new_n902_), .B2(new_n827_), .ZN(new_n903_));
  AOI21_X1  g702(.A(KEYINPUT121), .B1(new_n903_), .B2(new_n897_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n899_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n523_), .A2(new_n399_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n893_), .B1(new_n905_), .B2(new_n906_), .ZN(G1340gat));
  OAI21_X1  g706(.A(new_n397_), .B1(new_n645_), .B2(KEYINPUT60), .ZN(new_n908_));
  OAI211_X1 g707(.A(new_n892_), .B(new_n908_), .C1(KEYINPUT60), .C2(new_n397_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n903_), .A2(new_n679_), .A3(new_n897_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n911_), .B2(new_n397_), .ZN(G1341gat));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n902_), .A2(new_n715_), .A3(new_n827_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(G127gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n892_), .A2(new_n658_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n916_), .A2(KEYINPUT122), .A3(new_n394_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n715_), .A2(new_n394_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n905_), .B2(new_n919_), .ZN(G1342gat));
  INV_X1    g719(.A(new_n675_), .ZN(new_n921_));
  AOI21_X1  g720(.A(G134gat), .B1(new_n892_), .B2(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n596_), .A2(new_n392_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n905_), .B2(new_n923_), .ZN(G1343gat));
  NOR3_X1   g723(.A1(new_n902_), .A2(new_n466_), .A3(new_n421_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n748_), .A2(new_n445_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n925_), .A2(new_n522_), .A3(new_n926_), .ZN(new_n927_));
  XNOR2_X1  g726(.A(KEYINPUT123), .B(G141gat), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1344gat));
  NAND3_X1  g728(.A1(new_n925_), .A2(new_n679_), .A3(new_n926_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g730(.A1(new_n925_), .A2(new_n658_), .A3(new_n926_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(KEYINPUT61), .B(G155gat), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1346gat));
  INV_X1    g733(.A(G162gat), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n925_), .A2(new_n935_), .A3(new_n921_), .A4(new_n926_), .ZN(new_n936_));
  AND3_X1   g735(.A1(new_n925_), .A2(new_n731_), .A3(new_n926_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n937_), .B2(new_n935_), .ZN(G1347gat));
  NOR3_X1   g737(.A1(new_n802_), .A2(new_n473_), .A3(new_n446_), .ZN(new_n939_));
  AND2_X1   g738(.A1(new_n895_), .A2(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n522_), .ZN(new_n941_));
  OAI21_X1  g740(.A(KEYINPUT62), .B1(new_n941_), .B2(KEYINPUT22), .ZN(new_n942_));
  OAI21_X1  g741(.A(G169gat), .B1(new_n941_), .B2(KEYINPUT62), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n944_), .B1(new_n289_), .B2(new_n942_), .ZN(G1348gat));
  NAND2_X1  g744(.A1(new_n879_), .A2(new_n891_), .ZN(new_n946_));
  AND2_X1   g745(.A1(new_n946_), .A2(new_n939_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n645_), .A2(new_n290_), .ZN(new_n948_));
  AND3_X1   g747(.A1(new_n947_), .A2(KEYINPUT124), .A3(new_n948_), .ZN(new_n949_));
  AOI21_X1  g748(.A(KEYINPUT124), .B1(new_n947_), .B2(new_n948_), .ZN(new_n950_));
  AOI21_X1  g749(.A(G176gat), .B1(new_n940_), .B2(new_n679_), .ZN(new_n951_));
  NOR3_X1   g750(.A1(new_n949_), .A2(new_n950_), .A3(new_n951_), .ZN(G1349gat));
  NOR2_X1   g751(.A1(new_n343_), .A2(new_n316_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n940_), .A2(new_n953_), .A3(new_n658_), .ZN(new_n954_));
  AND3_X1   g753(.A1(new_n946_), .A2(new_n658_), .A3(new_n939_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n954_), .B1(new_n955_), .B2(new_n327_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT125), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n956_), .A2(new_n957_), .ZN(new_n958_));
  OAI211_X1 g757(.A(KEYINPUT125), .B(new_n954_), .C1(new_n955_), .C2(new_n327_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1350gat));
  NAND4_X1  g759(.A1(new_n940_), .A2(new_n311_), .A3(new_n342_), .A4(new_n921_), .ZN(new_n961_));
  AND2_X1   g760(.A1(new_n940_), .A2(new_n731_), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n961_), .B1(new_n962_), .B2(new_n310_), .ZN(G1351gat));
  NOR2_X1   g762(.A1(new_n802_), .A2(new_n663_), .ZN(new_n964_));
  NAND3_X1  g763(.A1(new_n925_), .A2(new_n522_), .A3(new_n964_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g765(.A1(new_n925_), .A2(new_n964_), .ZN(new_n967_));
  INV_X1    g766(.A(KEYINPUT126), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n968_), .A2(G204gat), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n967_), .A2(new_n679_), .A3(new_n969_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n925_), .A2(new_n964_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n971_), .A2(new_n645_), .ZN(new_n972_));
  XNOR2_X1  g771(.A(KEYINPUT126), .B(G204gat), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n970_), .B1(new_n972_), .B2(new_n973_), .ZN(G1353gat));
  AOI21_X1  g773(.A(new_n715_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n925_), .A2(new_n964_), .A3(new_n975_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n977_));
  XNOR2_X1  g776(.A(new_n977_), .B(KEYINPUT127), .ZN(new_n978_));
  XNOR2_X1  g777(.A(new_n976_), .B(new_n978_), .ZN(G1354gat));
  OR3_X1    g778(.A1(new_n971_), .A2(G218gat), .A3(new_n675_), .ZN(new_n980_));
  OAI21_X1  g779(.A(G218gat), .B1(new_n971_), .B2(new_n596_), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n980_), .A2(new_n981_), .ZN(G1355gat));
endmodule


