//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n951_, new_n953_, new_n954_, new_n956_,
    new_n957_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n982_, new_n983_,
    new_n985_, new_n986_, new_n987_, new_n989_, new_n990_, new_n991_,
    new_n992_, new_n994_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1001_, new_n1002_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT69), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G134gat), .B(G162gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT36), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT15), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G29gat), .B(G36gat), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(KEYINPUT67), .ZN(new_n209_));
  INV_X1    g008(.A(G36gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G29gat), .ZN(new_n211_));
  INV_X1    g010(.A(G29gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G36gat), .ZN(new_n213_));
  AND3_X1   g012(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT67), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT68), .B1(new_n209_), .B2(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G43gat), .B(G50gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(new_n213_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT67), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n208_), .A2(KEYINPUT67), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT68), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n215_), .A2(new_n216_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n216_), .B1(new_n215_), .B2(new_n222_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n207_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n215_), .A2(new_n222_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n216_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(KEYINPUT15), .A3(new_n223_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G99gat), .A2(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT6), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT6), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(G99gat), .A3(G106gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n236_));
  INV_X1    g035(.A(G106gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G85gat), .ZN(new_n240_));
  INV_X1    g039(.A(G92gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G85gat), .A2(G92gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(KEYINPUT9), .A3(new_n243_), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n243_), .A2(KEYINPUT9), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n235_), .A2(new_n239_), .A3(new_n244_), .A4(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n242_), .A2(new_n243_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT7), .ZN(new_n248_));
  INV_X1    g047(.A(G99gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n249_), .A3(new_n237_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  AOI211_X1 g051(.A(KEYINPUT8), .B(new_n247_), .C1(new_n252_), .C2(new_n235_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT8), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n235_), .A2(new_n251_), .A3(new_n250_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n247_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n254_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n246_), .B1(new_n253_), .B2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n226_), .A2(new_n230_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n229_), .A2(new_n223_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n246_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n232_), .A2(new_n234_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n250_), .A2(new_n251_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n256_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT8), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n255_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n261_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT35), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G232gat), .A2(G233gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(KEYINPUT34), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  AOI22_X1  g070(.A1(new_n260_), .A2(new_n267_), .B1(new_n268_), .B2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n268_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n259_), .A2(new_n272_), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n274_), .B1(new_n259_), .B2(new_n272_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n206_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n259_), .A2(new_n272_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n273_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n259_), .A2(new_n272_), .A3(new_n274_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT36), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n205_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT70), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n279_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n277_), .A2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT72), .B1(new_n285_), .B2(KEYINPUT37), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n277_), .A2(KEYINPUT71), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n288_), .B(new_n206_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n289_), .A3(new_n284_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n286_), .B1(KEYINPUT37), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT72), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n290_), .A2(new_n292_), .A3(KEYINPUT37), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT73), .B(G8gat), .ZN(new_n295_));
  INV_X1    g094(.A(G1gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT14), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G15gat), .B(G22gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT74), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G1gat), .B(G8gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n299_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n301_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G57gat), .B(G64gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G71gat), .B(G78gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(KEYINPUT11), .ZN(new_n311_));
  INV_X1    g110(.A(new_n310_), .ZN(new_n312_));
  INV_X1    g111(.A(G64gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(G57gat), .ZN(new_n314_));
  INV_X1    g113(.A(G57gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(G64gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n316_), .A3(KEYINPUT11), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n309_), .A2(KEYINPUT11), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n311_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n308_), .A2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G231gat), .A2(G233gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n322_), .B(KEYINPUT75), .Z(new_n323_));
  AOI21_X1  g122(.A(new_n320_), .B1(new_n302_), .B2(new_n306_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n321_), .A2(new_n323_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n323_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n320_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n307_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n327_), .B1(new_n329_), .B2(new_n324_), .ZN(new_n330_));
  XOR2_X1   g129(.A(G127gat), .B(G155gat), .Z(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT16), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G183gat), .B(G211gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT17), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n326_), .A2(new_n330_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT77), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n326_), .A2(new_n330_), .A3(KEYINPUT77), .A4(new_n335_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n326_), .A2(new_n330_), .ZN(new_n341_));
  XOR2_X1   g140(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n342_));
  NOR2_X1   g141(.A1(new_n334_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n340_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n294_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n348_), .A2(KEYINPUT78), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(KEYINPUT78), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT13), .ZN(new_n351_));
  INV_X1    g150(.A(G230gat), .ZN(new_n352_));
  INV_X1    g151(.A(G233gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n267_), .B2(new_n320_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT65), .B1(new_n267_), .B2(new_n320_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT12), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n258_), .A2(new_n328_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(KEYINPUT65), .A3(KEYINPUT12), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n356_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  OAI211_X1 g161(.A(new_n246_), .B(new_n320_), .C1(new_n253_), .C2(new_n257_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT64), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(new_n360_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n362_), .B1(new_n354_), .B2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G120gat), .B(G148gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT5), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G176gat), .B(G204gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT66), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n366_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n366_), .A2(new_n370_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n351_), .B1(new_n373_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n373_), .A2(new_n351_), .A3(new_n374_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n308_), .A2(new_n230_), .A3(new_n226_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n307_), .A2(new_n260_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G229gat), .A2(G233gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n381_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n380_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n307_), .A2(new_n260_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n383_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G113gat), .B(G141gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G169gat), .B(G197gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n387_), .B(new_n388_), .Z(new_n389_));
  NAND3_X1  g188(.A1(new_n382_), .A2(new_n386_), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n389_), .B1(new_n382_), .B2(new_n386_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n378_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G228gat), .A2(G233gat), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT86), .ZN(new_n398_));
  INV_X1    g197(.A(G155gat), .ZN(new_n399_));
  INV_X1    g198(.A(G162gat), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(KEYINPUT84), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT84), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(G155gat), .B2(G162gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G155gat), .A2(G162gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n407_));
  NOR3_X1   g206(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT85), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(G141gat), .A2(G148gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT2), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT2), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n414_), .A2(G141gat), .A3(G148gat), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n413_), .A2(new_n415_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n406_), .B1(new_n411_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n412_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(G141gat), .A2(G148gat), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n405_), .A2(KEYINPUT1), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT1), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n423_), .A2(G155gat), .A3(G162gat), .ZN(new_n424_));
  AND2_X1   g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n421_), .B1(new_n404_), .B2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT29), .B1(new_n417_), .B2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(G197gat), .A2(G204gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(G197gat), .A2(G204gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n429_), .A2(KEYINPUT21), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT21), .ZN(new_n432_));
  AND2_X1   g231(.A1(G197gat), .A2(G204gat), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n432_), .B1(new_n433_), .B2(new_n428_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G211gat), .B(G218gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n431_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n435_), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n433_), .A2(new_n428_), .A3(new_n432_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n398_), .B1(new_n427_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT29), .ZN(new_n442_));
  AOI22_X1  g241(.A1(new_n401_), .A2(new_n403_), .B1(G155gat), .B2(G162gat), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT3), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n419_), .A2(new_n409_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n414_), .B1(G141gat), .B2(G148gat), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n412_), .A2(KEYINPUT2), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n443_), .B1(new_n448_), .B2(new_n410_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n401_), .A2(new_n403_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n422_), .A2(new_n424_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n420_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n442_), .B1(new_n449_), .B2(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n436_), .A2(new_n439_), .ZN(new_n454_));
  NOR3_X1   g253(.A1(new_n453_), .A2(KEYINPUT86), .A3(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n397_), .B1(new_n441_), .B2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G78gat), .B(G106gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT86), .B1(new_n453_), .B2(new_n454_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n419_), .A2(new_n444_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT85), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n413_), .A2(new_n415_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n460_), .A2(new_n461_), .A3(new_n407_), .A4(new_n445_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n425_), .A2(new_n404_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n462_), .A2(new_n443_), .B1(new_n463_), .B2(new_n420_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n398_), .B(new_n440_), .C1(new_n464_), .C2(new_n442_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n458_), .A2(new_n465_), .A3(G228gat), .A4(G233gat), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n456_), .A2(new_n457_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT88), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n457_), .B(KEYINPUT87), .Z(new_n470_));
  NOR3_X1   g269(.A1(new_n441_), .A2(new_n455_), .A3(new_n397_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n458_), .A2(new_n465_), .B1(G228gat), .B2(G233gat), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n470_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n464_), .A2(new_n442_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(KEYINPUT28), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n474_), .A2(KEYINPUT28), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G22gat), .B(G50gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NOR3_X1   g278(.A1(new_n476_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n474_), .A2(KEYINPUT28), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n478_), .B1(new_n481_), .B2(new_n475_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n456_), .A2(KEYINPUT88), .A3(new_n466_), .A4(new_n457_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n469_), .A2(new_n473_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n471_), .A2(new_n470_), .A3(new_n472_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n470_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n487_), .B1(new_n456_), .B2(new_n466_), .ZN(new_n488_));
  OAI22_X1  g287(.A1(new_n486_), .A2(new_n488_), .B1(new_n480_), .B2(new_n482_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G8gat), .B(G36gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT18), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G64gat), .B(G92gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(G190gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT26), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT26), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G190gat), .ZN(new_n499_));
  INV_X1    g298(.A(G183gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT25), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT25), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(G183gat), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n497_), .A2(new_n499_), .A3(new_n501_), .A4(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G169gat), .ZN(new_n505_));
  INV_X1    g304(.A(G176gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G169gat), .A2(G176gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(KEYINPUT24), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n504_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT91), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n504_), .A2(KEYINPUT91), .A3(new_n509_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G183gat), .A2(G190gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT23), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT23), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n516_), .A2(G183gat), .A3(G190gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  OR3_X1    g317(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n512_), .A2(new_n513_), .A3(new_n520_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n518_), .B1(G183gat), .B2(G190gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n505_), .A2(KEYINPUT22), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT22), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(G169gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n525_), .A3(new_n506_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n508_), .B(KEYINPUT92), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n522_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n454_), .B1(new_n521_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n531_));
  NAND2_X1  g330(.A1(KEYINPUT79), .A2(G190gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(KEYINPUT26), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT80), .ZN(new_n534_));
  AND3_X1   g333(.A1(new_n499_), .A2(new_n501_), .A3(new_n503_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT80), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n531_), .A2(new_n536_), .A3(KEYINPUT26), .A4(new_n532_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n534_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n509_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n531_), .A2(new_n500_), .A3(new_n532_), .ZN(new_n541_));
  AOI22_X1  g340(.A1(new_n541_), .A2(new_n518_), .B1(G169gat), .B2(G176gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n526_), .A2(KEYINPUT81), .ZN(new_n543_));
  XNOR2_X1  g342(.A(KEYINPUT22), .B(G169gat), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT81), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n506_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n542_), .A2(new_n543_), .A3(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n540_), .A2(new_n454_), .A3(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G226gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT90), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n530_), .A2(KEYINPUT20), .A3(new_n548_), .A4(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT20), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n540_), .A2(new_n547_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n555_), .B2(new_n440_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n513_), .A2(new_n520_), .ZN(new_n557_));
  AOI21_X1  g356(.A(KEYINPUT91), .B1(new_n504_), .B2(new_n509_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n454_), .B(new_n528_), .C1(new_n557_), .C2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n551_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT95), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n553_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n551_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n543_), .A2(new_n546_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n564_), .A2(new_n542_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT20), .B1(new_n565_), .B2(new_n454_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n559_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n563_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(KEYINPUT95), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n495_), .B1(new_n562_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n552_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n548_), .A2(KEYINPUT20), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n571_), .B1(new_n572_), .B2(new_n529_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n555_), .A2(new_n440_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n574_), .A2(KEYINPUT20), .A3(new_n551_), .A4(new_n559_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n573_), .A2(new_n494_), .A3(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT27), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n573_), .A2(new_n575_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n495_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n573_), .A2(new_n494_), .A3(new_n575_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n570_), .A2(new_n578_), .B1(new_n582_), .B2(new_n577_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G127gat), .B(G134gat), .Z(new_n584_));
  INV_X1    g383(.A(G120gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(G113gat), .ZN(new_n586_));
  INV_X1    g385(.A(G113gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(G120gat), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n586_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n584_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G127gat), .B(G134gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G113gat), .B(G120gat), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n590_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n449_), .A2(new_n452_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT83), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n584_), .A2(new_n589_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n591_), .A2(new_n592_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n596_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n596_), .B1(new_n584_), .B2(new_n589_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  OAI211_X1 g401(.A(KEYINPUT4), .B(new_n595_), .C1(new_n602_), .C2(new_n464_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G225gat), .A2(G233gat), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n600_), .B1(new_n594_), .B2(new_n596_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n449_), .A2(new_n452_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT4), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n606_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n603_), .A2(new_n605_), .A3(new_n609_), .ZN(new_n610_));
  OAI211_X1 g409(.A(new_n595_), .B(new_n604_), .C1(new_n602_), .C2(new_n464_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G1gat), .B(G29gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(G85gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT0), .B(G57gat), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n613_), .B(new_n614_), .Z(new_n615_));
  AND3_X1   g414(.A1(new_n610_), .A2(new_n611_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n490_), .A2(new_n583_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n494_), .A2(KEYINPUT32), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n572_), .A2(new_n529_), .ZN(new_n621_));
  AOI22_X1  g420(.A1(new_n568_), .A2(KEYINPUT95), .B1(new_n621_), .B2(new_n552_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n560_), .A2(new_n561_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n620_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n573_), .A2(new_n620_), .A3(new_n575_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n625_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT93), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n494_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n628_), .B1(new_n576_), .B2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n580_), .A2(KEYINPUT93), .A3(new_n581_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n610_), .A2(new_n611_), .A3(new_n615_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n595_), .B1(new_n602_), .B2(new_n464_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n615_), .B1(new_n637_), .B2(new_n605_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n603_), .A2(new_n604_), .A3(new_n609_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n635_), .A2(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n610_), .A2(KEYINPUT33), .A3(new_n611_), .A4(new_n615_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT94), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n609_), .A2(new_n605_), .ZN(new_n644_));
  AOI22_X1  g443(.A1(new_n644_), .A2(new_n603_), .B1(new_n637_), .B2(new_n604_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT94), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(KEYINPUT33), .A4(new_n615_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n641_), .B1(new_n643_), .B2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n627_), .B1(new_n632_), .B2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n619_), .B1(new_n649_), .B2(new_n490_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(G71gat), .B(G99gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(G43gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n555_), .B(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT82), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n602_), .A2(KEYINPUT31), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n602_), .A2(KEYINPUT31), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n655_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(G227gat), .A2(G233gat), .ZN(new_n659_));
  INV_X1    g458(.A(G15gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT30), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n658_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n658_), .A2(new_n663_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n654_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n666_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n668_), .A2(new_n653_), .A3(new_n664_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT96), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n570_), .A2(new_n578_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n577_), .B1(new_n576_), .B2(new_n629_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n673_), .A2(new_n485_), .A3(new_n489_), .A4(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n670_), .A2(new_n618_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n485_), .A2(new_n489_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n618_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n669_), .B2(new_n667_), .ZN(new_n680_));
  NAND4_X1  g479(.A1(new_n678_), .A2(new_n680_), .A3(KEYINPUT96), .A4(new_n583_), .ZN(new_n681_));
  AOI22_X1  g480(.A1(new_n650_), .A2(new_n671_), .B1(new_n677_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  AND4_X1   g482(.A1(new_n349_), .A2(new_n350_), .A3(new_n396_), .A4(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(new_n296_), .A3(new_n679_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT38), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n285_), .ZN(new_n688_));
  NOR4_X1   g487(.A1(new_n682_), .A2(new_n395_), .A3(new_n688_), .A4(new_n345_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n296_), .B1(new_n689_), .B2(new_n679_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n685_), .A2(new_n686_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(KEYINPUT97), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(KEYINPUT97), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n691_), .B1(new_n693_), .B2(new_n694_), .ZN(G1324gat));
  INV_X1    g494(.A(new_n583_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n684_), .A2(new_n295_), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n689_), .A2(new_n696_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT39), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n698_), .A2(new_n699_), .A3(G8gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n698_), .B2(G8gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g502(.A1(new_n684_), .A2(new_n660_), .A3(new_n670_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n689_), .A2(new_n670_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(G15gat), .ZN(new_n706_));
  XNOR2_X1  g505(.A(KEYINPUT98), .B(KEYINPUT41), .ZN(new_n707_));
  OR2_X1    g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n707_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n704_), .A2(new_n708_), .A3(new_n709_), .ZN(G1326gat));
  INV_X1    g509(.A(G22gat), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n684_), .A2(new_n711_), .A3(new_n490_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n689_), .A2(new_n490_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G22gat), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n714_), .A2(KEYINPUT42), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(KEYINPUT42), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(G1327gat));
  NOR2_X1   g516(.A1(new_n346_), .A2(new_n285_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n683_), .A2(new_n396_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(G29gat), .B1(new_n720_), .B2(new_n679_), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n490_), .A2(new_n583_), .A3(new_n618_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n624_), .A2(new_n626_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n647_), .A2(new_n643_), .ZN(new_n724_));
  AOI22_X1  g523(.A1(new_n633_), .A2(new_n634_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n724_), .A2(new_n630_), .A3(new_n631_), .A4(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n490_), .B1(new_n723_), .B2(new_n726_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n671_), .B1(new_n722_), .B2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n677_), .A2(new_n681_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(KEYINPUT100), .A3(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n290_), .A2(new_n292_), .A3(KEYINPUT37), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n290_), .A2(KEYINPUT37), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n732_), .B2(new_n286_), .ZN(new_n733_));
  AND2_X1   g532(.A1(KEYINPUT100), .A2(KEYINPUT43), .ZN(new_n734_));
  OAI211_X1 g533(.A(new_n730_), .B(new_n733_), .C1(new_n682_), .C2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT99), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT43), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(KEYINPUT43), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n738_), .B1(new_n682_), .B2(new_n294_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n395_), .A2(new_n346_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n735_), .A2(new_n737_), .A3(new_n739_), .A4(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n737_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n729_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n723_), .A2(new_n726_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(new_n678_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n670_), .B1(new_n747_), .B2(new_n619_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n733_), .B1(new_n745_), .B2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n744_), .B1(new_n749_), .B2(new_n738_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n750_), .A2(KEYINPUT44), .A3(new_n735_), .A4(new_n740_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n743_), .A2(new_n751_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n618_), .A2(new_n212_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n721_), .B1(new_n752_), .B2(new_n753_), .ZN(G1328gat));
  NOR3_X1   g553(.A1(new_n719_), .A2(G36gat), .A3(new_n583_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n743_), .A2(new_n696_), .A3(new_n751_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n758_), .A2(KEYINPUT101), .A3(G36gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT101), .B1(new_n758_), .B2(G36gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n757_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT46), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  OAI211_X1 g562(.A(KEYINPUT46), .B(new_n757_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1329gat));
  NAND3_X1  g564(.A1(new_n752_), .A2(G43gat), .A3(new_n670_), .ZN(new_n766_));
  INV_X1    g565(.A(G43gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n767_), .B1(new_n719_), .B2(new_n671_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g569(.A(G50gat), .B1(new_n720_), .B2(new_n490_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n490_), .A2(G50gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n752_), .B2(new_n772_), .ZN(G1331gat));
  INV_X1    g572(.A(new_n378_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n349_), .A2(new_n350_), .A3(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT103), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n682_), .A2(new_n394_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n349_), .A2(KEYINPUT103), .A3(new_n350_), .A4(new_n774_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n777_), .A2(new_n679_), .A3(new_n778_), .A4(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT104), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n315_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n780_), .B2(new_n315_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n393_), .A2(new_n344_), .A3(new_n340_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n683_), .A2(new_n285_), .A3(new_n774_), .A4(new_n785_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n786_), .A2(KEYINPUT105), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(KEYINPUT105), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n787_), .A2(G57gat), .A3(new_n679_), .A4(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT106), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n782_), .A2(new_n783_), .A3(new_n790_), .ZN(G1332gat));
  AND3_X1   g590(.A1(new_n777_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n792_), .A2(new_n313_), .A3(new_n696_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n787_), .A2(new_n696_), .A3(new_n788_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT48), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n794_), .A2(new_n795_), .A3(G64gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n794_), .B2(G64gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n793_), .B1(new_n796_), .B2(new_n797_), .ZN(G1333gat));
  INV_X1    g597(.A(G71gat), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n792_), .A2(new_n799_), .A3(new_n670_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n787_), .A2(new_n670_), .A3(new_n788_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT49), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n801_), .A2(new_n802_), .A3(G71gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n801_), .B2(G71gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(G1334gat));
  NOR2_X1   g604(.A1(new_n678_), .A2(G78gat), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n806_), .B(KEYINPUT107), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n792_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n787_), .A2(new_n490_), .A3(new_n788_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT50), .ZN(new_n810_));
  AND3_X1   g609(.A1(new_n809_), .A2(new_n810_), .A3(G78gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n810_), .B1(new_n809_), .B2(G78gat), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n808_), .B1(new_n811_), .B2(new_n812_), .ZN(G1335gat));
  NOR3_X1   g612(.A1(new_n378_), .A2(new_n346_), .A3(new_n394_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n750_), .A2(new_n735_), .A3(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(G85gat), .B1(new_n815_), .B2(new_n618_), .ZN(new_n816_));
  AND3_X1   g615(.A1(new_n778_), .A2(new_n774_), .A3(new_n718_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n240_), .A3(new_n679_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1336gat));
  OAI21_X1  g618(.A(G92gat), .B1(new_n815_), .B2(new_n583_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(new_n241_), .A3(new_n696_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1337gat));
  OAI21_X1  g621(.A(G99gat), .B1(new_n815_), .B2(new_n671_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n670_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT108), .B1(new_n817_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(new_n826_));
  XOR2_X1   g625(.A(KEYINPUT109), .B(KEYINPUT51), .Z(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(G1338gat));
  XNOR2_X1  g627(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n829_));
  INV_X1    g628(.A(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n750_), .A2(new_n490_), .A3(new_n735_), .A4(new_n814_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n237_), .B1(new_n832_), .B2(KEYINPUT111), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT111), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n831_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(KEYINPUT52), .A3(new_n835_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n678_), .A2(G106gat), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n817_), .A2(new_n837_), .ZN(new_n838_));
  XOR2_X1   g637(.A(new_n838_), .B(KEYINPUT110), .Z(new_n839_));
  NAND2_X1  g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT52), .B1(new_n833_), .B2(new_n835_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n830_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n833_), .A2(new_n835_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n845_), .A2(new_n836_), .A3(new_n839_), .A4(new_n829_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n842_), .A2(new_n846_), .ZN(G1339gat));
  XNOR2_X1  g646(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT114), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n785_), .A2(new_n378_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n733_), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n848_), .A2(new_n849_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n294_), .A2(new_n378_), .A3(new_n785_), .A4(new_n853_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n373_), .A2(new_n374_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT116), .ZN(new_n857_));
  OR2_X1    g656(.A1(new_n307_), .A2(new_n260_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n383_), .B1(new_n858_), .B2(new_n380_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n857_), .B1(new_n859_), .B2(new_n389_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n381_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n389_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(KEYINPUT116), .A3(new_n862_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n379_), .A2(new_n380_), .A3(new_n383_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n860_), .A2(new_n863_), .A3(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n856_), .A2(new_n865_), .A3(new_n390_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT115), .B1(new_n362_), .B2(KEYINPUT55), .ZN(new_n867_));
  AOI21_X1  g666(.A(KEYINPUT12), .B1(new_n360_), .B2(KEYINPUT65), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT65), .ZN(new_n869_));
  AOI211_X1 g668(.A(new_n869_), .B(new_n358_), .C1(new_n258_), .C2(new_n328_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n355_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT55), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n362_), .A2(KEYINPUT55), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n364_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n354_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n867_), .A2(new_n874_), .A3(new_n875_), .A4(new_n877_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n878_), .A2(KEYINPUT56), .A3(new_n371_), .ZN(new_n879_));
  AOI21_X1  g678(.A(KEYINPUT56), .B1(new_n878_), .B2(new_n371_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n374_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n866_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n883_), .A2(KEYINPUT57), .A3(new_n285_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n285_), .ZN(new_n885_));
  XOR2_X1   g684(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n878_), .A2(KEYINPUT56), .A3(new_n371_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n878_), .A2(new_n371_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT56), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n878_), .A2(KEYINPUT118), .A3(KEYINPUT56), .A4(new_n371_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n891_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n865_), .A2(new_n390_), .A3(new_n374_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n733_), .ZN(new_n901_));
  AND3_X1   g700(.A1(new_n896_), .A2(KEYINPUT58), .A3(new_n897_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n884_), .B(new_n888_), .C1(new_n901_), .C2(new_n902_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n855_), .B1(new_n903_), .B2(new_n345_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n675_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n671_), .A2(new_n618_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  OAI21_X1  g706(.A(KEYINPUT59), .B1(new_n904_), .B2(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n393_), .A2(new_n587_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(KEYINPUT121), .ZN(new_n910_));
  AOI21_X1  g709(.A(KEYINPUT58), .B1(new_n896_), .B2(new_n897_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n902_), .A2(new_n911_), .A3(new_n294_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n886_), .B1(new_n883_), .B2(new_n285_), .ZN(new_n913_));
  OAI21_X1  g712(.A(KEYINPUT120), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT120), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n915_), .B(new_n888_), .C1(new_n901_), .C2(new_n902_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n914_), .A2(new_n884_), .A3(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n855_), .B1(new_n917_), .B2(new_n345_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n907_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n908_), .B(new_n910_), .C1(new_n918_), .C2(new_n921_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n904_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n923_), .A2(new_n394_), .A3(new_n919_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n587_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n922_), .A2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(KEYINPUT122), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n922_), .A2(new_n925_), .A3(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n927_), .A2(new_n929_), .ZN(G1340gat));
  OAI21_X1  g729(.A(new_n908_), .B1(new_n918_), .B2(new_n921_), .ZN(new_n931_));
  OAI21_X1  g730(.A(G120gat), .B1(new_n931_), .B2(new_n378_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n904_), .A2(new_n907_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n585_), .B1(new_n378_), .B2(KEYINPUT60), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n935_), .B1(KEYINPUT60), .B2(new_n585_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n932_), .B1(new_n934_), .B2(new_n936_), .ZN(G1341gat));
  AOI21_X1  g736(.A(G127gat), .B1(new_n933_), .B2(new_n346_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n931_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n346_), .A2(G127gat), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(KEYINPUT123), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n938_), .B1(new_n939_), .B2(new_n941_), .ZN(G1342gat));
  OAI21_X1  g741(.A(G134gat), .B1(new_n931_), .B2(new_n294_), .ZN(new_n943_));
  OR2_X1    g742(.A1(new_n285_), .A2(G134gat), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n934_), .B2(new_n944_), .ZN(G1343gat));
  NAND4_X1  g744(.A1(new_n490_), .A2(new_n583_), .A3(new_n679_), .A4(new_n671_), .ZN(new_n946_));
  XOR2_X1   g745(.A(new_n946_), .B(KEYINPUT124), .Z(new_n947_));
  NAND2_X1  g746(.A1(new_n923_), .A2(new_n947_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n948_), .A2(new_n393_), .ZN(new_n949_));
  XOR2_X1   g748(.A(new_n949_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g749(.A1(new_n948_), .A2(new_n378_), .ZN(new_n951_));
  XOR2_X1   g750(.A(new_n951_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g751(.A1(new_n948_), .A2(new_n345_), .ZN(new_n953_));
  XOR2_X1   g752(.A(KEYINPUT61), .B(G155gat), .Z(new_n954_));
  XNOR2_X1  g753(.A(new_n953_), .B(new_n954_), .ZN(G1346gat));
  OAI21_X1  g754(.A(G162gat), .B1(new_n948_), .B2(new_n294_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n688_), .A2(new_n400_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n948_), .B2(new_n957_), .ZN(G1347gat));
  NOR3_X1   g757(.A1(new_n676_), .A2(new_n490_), .A3(new_n583_), .ZN(new_n959_));
  INV_X1    g758(.A(new_n884_), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n888_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n960_), .B1(new_n961_), .B2(KEYINPUT120), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n346_), .B1(new_n962_), .B2(new_n916_), .ZN(new_n963_));
  OAI211_X1 g762(.A(new_n394_), .B(new_n959_), .C1(new_n963_), .C2(new_n855_), .ZN(new_n964_));
  XOR2_X1   g763(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n965_));
  INV_X1    g764(.A(new_n965_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n505_), .B1(new_n966_), .B2(KEYINPUT126), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n964_), .A2(new_n967_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n966_), .A2(KEYINPUT126), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n968_), .A2(new_n969_), .ZN(new_n970_));
  INV_X1    g769(.A(new_n959_), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n918_), .A2(new_n971_), .ZN(new_n972_));
  NAND3_X1  g771(.A1(new_n972_), .A2(new_n394_), .A3(new_n544_), .ZN(new_n973_));
  OAI211_X1 g772(.A(new_n964_), .B(new_n967_), .C1(KEYINPUT126), .C2(new_n966_), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n970_), .A2(new_n973_), .A3(new_n974_), .ZN(G1348gat));
  AOI21_X1  g774(.A(G176gat), .B1(new_n972_), .B2(new_n774_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n904_), .A2(new_n971_), .ZN(new_n977_));
  NAND3_X1  g776(.A1(new_n977_), .A2(G176gat), .A3(new_n774_), .ZN(new_n978_));
  NAND2_X1  g777(.A1(new_n978_), .A2(KEYINPUT127), .ZN(new_n979_));
  OR2_X1    g778(.A1(new_n978_), .A2(KEYINPUT127), .ZN(new_n980_));
  AOI21_X1  g779(.A(new_n976_), .B1(new_n979_), .B2(new_n980_), .ZN(G1349gat));
  AOI21_X1  g780(.A(G183gat), .B1(new_n977_), .B2(new_n346_), .ZN(new_n982_));
  AOI21_X1  g781(.A(new_n345_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n983_));
  AOI21_X1  g782(.A(new_n982_), .B1(new_n972_), .B2(new_n983_), .ZN(G1350gat));
  OAI21_X1  g783(.A(new_n959_), .B1(new_n963_), .B2(new_n855_), .ZN(new_n985_));
  OAI21_X1  g784(.A(G190gat), .B1(new_n985_), .B2(new_n294_), .ZN(new_n986_));
  NAND3_X1  g785(.A1(new_n688_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n987_));
  OAI21_X1  g786(.A(new_n986_), .B1(new_n985_), .B2(new_n987_), .ZN(G1351gat));
  NOR4_X1   g787(.A1(new_n678_), .A2(new_n583_), .A3(new_n679_), .A4(new_n670_), .ZN(new_n989_));
  NAND2_X1  g788(.A1(new_n923_), .A2(new_n989_), .ZN(new_n990_));
  INV_X1    g789(.A(new_n990_), .ZN(new_n991_));
  NAND2_X1  g790(.A1(new_n991_), .A2(new_n394_), .ZN(new_n992_));
  XNOR2_X1  g791(.A(new_n992_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g792(.A1(new_n991_), .A2(new_n774_), .ZN(new_n994_));
  XNOR2_X1  g793(.A(new_n994_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g794(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n996_));
  AND2_X1   g795(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n997_));
  NOR4_X1   g796(.A1(new_n990_), .A2(new_n345_), .A3(new_n996_), .A4(new_n997_), .ZN(new_n998_));
  NAND2_X1  g797(.A1(new_n991_), .A2(new_n346_), .ZN(new_n999_));
  AOI21_X1  g798(.A(new_n998_), .B1(new_n999_), .B2(new_n996_), .ZN(G1354gat));
  OR3_X1    g799(.A1(new_n990_), .A2(G218gat), .A3(new_n285_), .ZN(new_n1001_));
  OAI21_X1  g800(.A(G218gat), .B1(new_n990_), .B2(new_n294_), .ZN(new_n1002_));
  NAND2_X1  g801(.A1(new_n1001_), .A2(new_n1002_), .ZN(G1355gat));
endmodule


