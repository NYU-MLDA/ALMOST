//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n629_, new_n630_,
    new_n631_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n837_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(G169gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  AND2_X1   g006(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n208_));
  NOR2_X1   g007(.A1(KEYINPUT82), .A2(KEYINPUT25), .ZN(new_n209_));
  OAI21_X1  g008(.A(G183gat), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n210_), .B(KEYINPUT83), .Z(new_n211_));
  INV_X1    g010(.A(KEYINPUT26), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n213_), .B1(KEYINPUT25), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G190gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(KEYINPUT26), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n218_), .A2(KEYINPUT84), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(KEYINPUT84), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n215_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n211_), .A2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n224_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(KEYINPUT85), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT24), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n203_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n207_), .B1(new_n222_), .B2(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G197gat), .B(G204gat), .Z(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(KEYINPUT21), .ZN(new_n235_));
  XOR2_X1   g034(.A(G211gat), .B(G218gat), .Z(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT89), .ZN(new_n238_));
  INV_X1    g037(.A(G197gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(G204gat), .ZN(new_n240_));
  OAI211_X1 g039(.A(KEYINPUT21), .B(new_n240_), .C1(new_n234_), .C2(new_n238_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n237_), .A2(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n234_), .A2(new_n236_), .A3(KEYINPUT21), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT20), .B1(new_n233_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT92), .ZN(new_n247_));
  INV_X1    g046(.A(new_n213_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT91), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n218_), .A3(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(KEYINPUT91), .B1(new_n213_), .B2(new_n217_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(KEYINPUT25), .B(G183gat), .Z(new_n253_));
  OAI211_X1 g052(.A(new_n247_), .B(new_n227_), .C1(new_n252_), .C2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n253_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n227_), .ZN(new_n256_));
  OAI21_X1  g055(.A(KEYINPUT92), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n254_), .A2(new_n257_), .A3(new_n231_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n246_), .B1(new_n258_), .B2(new_n207_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G226gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT19), .ZN(new_n261_));
  OR3_X1    g060(.A1(new_n245_), .A2(new_n259_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT20), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n263_), .B1(new_n233_), .B2(new_n244_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n258_), .A2(new_n207_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT96), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n244_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n258_), .A2(KEYINPUT96), .A3(new_n207_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n265_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n261_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n262_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G8gat), .B(G36gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT18), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n274_), .B(new_n275_), .Z(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n272_), .A2(new_n277_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n264_), .B(new_n271_), .C1(new_n244_), .C2(new_n266_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n261_), .B1(new_n245_), .B2(new_n259_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT27), .B1(new_n281_), .B2(new_n277_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n276_), .ZN(new_n283_));
  OAI22_X1  g082(.A1(new_n278_), .A2(new_n282_), .B1(new_n283_), .B2(KEYINPUT27), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G78gat), .B(G106gat), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT29), .ZN(new_n287_));
  INV_X1    g086(.A(G141gat), .ZN(new_n288_));
  INV_X1    g087(.A(G148gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT86), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n290_), .B1(new_n291_), .B2(KEYINPUT3), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT87), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(KEYINPUT2), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT2), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n294_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT3), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n299_), .A2(new_n288_), .A3(new_n289_), .A4(KEYINPUT86), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n292_), .A2(new_n296_), .A3(new_n298_), .A4(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(G155gat), .B(G162gat), .Z(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT88), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n306_));
  AND3_X1   g105(.A1(new_n290_), .A2(new_n293_), .A3(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n303_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n301_), .A2(KEYINPUT88), .A3(new_n302_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n287_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n310_), .A2(new_n246_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G228gat), .A2(G233gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OAI211_X1 g112(.A(G228gat), .B(G233gat), .C1(new_n310_), .C2(new_n246_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n286_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n313_), .A2(new_n314_), .A3(new_n286_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n308_), .A2(new_n309_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n319_), .A2(KEYINPUT29), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G22gat), .B(G50gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT28), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n320_), .B(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(new_n315_), .B2(KEYINPUT90), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n318_), .A2(new_n324_), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n316_), .A2(KEYINPUT90), .A3(new_n317_), .A4(new_n323_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n284_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT97), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G225gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT94), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G127gat), .B(G134gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G113gat), .B(G120gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n319_), .A2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n308_), .A2(new_n336_), .A3(new_n309_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(KEYINPUT4), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n336_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT4), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n333_), .B1(new_n340_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n339_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n333_), .B1(new_n345_), .B2(new_n341_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G1gat), .B(G29gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(G85gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT0), .B(G57gat), .ZN(new_n350_));
  XOR2_X1   g149(.A(new_n349_), .B(new_n350_), .Z(new_n351_));
  OR4_X1    g150(.A1(new_n330_), .A2(new_n344_), .A3(new_n347_), .A4(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n351_), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n340_), .A2(new_n343_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n353_), .B(new_n346_), .C1(new_n354_), .C2(new_n333_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n351_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n355_), .A2(new_n356_), .A3(new_n330_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G71gat), .B(G99gat), .ZN(new_n360_));
  INV_X1    g159(.A(G43gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n233_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(new_n336_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G227gat), .A2(G233gat), .ZN(new_n365_));
  INV_X1    g164(.A(G15gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT30), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT31), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n364_), .B(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n359_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n329_), .A2(new_n371_), .ZN(new_n372_));
  NOR3_X1   g171(.A1(new_n284_), .A2(new_n359_), .A3(new_n327_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT98), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT95), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n279_), .A2(new_n280_), .A3(new_n375_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n376_), .B(new_n262_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n276_), .A2(KEYINPUT32), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n281_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n378_), .A2(new_n375_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n374_), .B1(new_n383_), .B2(new_n358_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT93), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n283_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n281_), .B(new_n277_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT93), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n344_), .A2(new_n347_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n389_), .A2(new_n353_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n354_), .A2(new_n333_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n345_), .A2(new_n341_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n351_), .B1(new_n392_), .B2(new_n332_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n390_), .A2(KEYINPUT33), .B1(new_n391_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT33), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n356_), .A2(new_n395_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n386_), .A2(new_n388_), .A3(new_n394_), .A4(new_n396_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n377_), .A2(new_n378_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n398_), .A2(KEYINPUT98), .A3(new_n352_), .A4(new_n357_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n384_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n373_), .B1(new_n400_), .B2(new_n327_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n370_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n372_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT70), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G57gat), .B(G64gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT11), .ZN(new_n406_));
  XOR2_X1   g205(.A(G71gat), .B(G78gat), .Z(new_n407_));
  OR2_X1    g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n405_), .A2(KEYINPUT11), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n407_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT7), .ZN(new_n413_));
  INV_X1    g212(.A(G99gat), .ZN(new_n414_));
  INV_X1    g213(.A(G106gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT67), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G99gat), .A2(G106gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT6), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT6), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(G99gat), .A3(G106gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .A4(KEYINPUT67), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n418_), .A2(new_n423_), .A3(new_n424_), .A4(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT68), .ZN(new_n427_));
  AND2_X1   g226(.A1(G85gat), .A2(G92gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(G85gat), .A2(G92gat), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n426_), .A2(new_n427_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n427_), .B1(new_n426_), .B2(new_n430_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT8), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n426_), .A2(new_n430_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n435_), .A2(KEYINPUT68), .A3(new_n433_), .ZN(new_n436_));
  INV_X1    g235(.A(G92gat), .ZN(new_n437_));
  OAI22_X1  g236(.A1(new_n428_), .A2(new_n429_), .B1(KEYINPUT9), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(G85gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n437_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT9), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G85gat), .A2(G92gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n438_), .A2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT66), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT66), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n438_), .A2(new_n443_), .A3(new_n446_), .ZN(new_n447_));
  OR2_X1    g246(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n415_), .A3(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n450_), .A2(KEYINPUT65), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n450_), .A2(KEYINPUT65), .B1(new_n420_), .B2(new_n422_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n445_), .A2(new_n447_), .A3(new_n451_), .A4(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n436_), .A2(new_n453_), .ZN(new_n454_));
  OAI211_X1 g253(.A(KEYINPUT12), .B(new_n412_), .C1(new_n434_), .C2(new_n454_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n451_), .A2(new_n452_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n447_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n446_), .B1(new_n438_), .B2(new_n443_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n456_), .A2(new_n459_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n435_), .A2(KEYINPUT68), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n426_), .A2(new_n427_), .A3(new_n430_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(KEYINPUT8), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n411_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n464_));
  XOR2_X1   g263(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n455_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n460_), .A2(new_n463_), .A3(new_n411_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G230gat), .A2(G233gat), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n469_), .B(KEYINPUT64), .Z(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n404_), .B1(new_n467_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n470_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n468_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n473_), .B1(new_n474_), .B2(new_n464_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n434_), .A2(new_n454_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n473_), .B1(new_n476_), .B2(new_n411_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n412_), .B1(new_n434_), .B2(new_n454_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n465_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n477_), .A2(new_n479_), .A3(KEYINPUT70), .A4(new_n455_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n472_), .A2(new_n475_), .A3(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G120gat), .B(G148gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G176gat), .B(G204gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n481_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n486_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n472_), .A2(new_n475_), .A3(new_n480_), .A4(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT13), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G29gat), .B(G36gat), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n493_), .A2(KEYINPUT72), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(KEYINPUT72), .ZN(new_n495_));
  XOR2_X1   g294(.A(G43gat), .B(G50gat), .Z(new_n496_));
  OR3_X1    g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n496_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT15), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n497_), .A2(new_n498_), .A3(KEYINPUT15), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G1gat), .B(G8gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT75), .ZN(new_n504_));
  INV_X1    g303(.A(G22gat), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n366_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G15gat), .A2(G22gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G1gat), .A2(G8gat), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n506_), .A2(new_n507_), .B1(KEYINPUT14), .B2(new_n508_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n504_), .B(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n501_), .A2(new_n502_), .A3(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(new_n504_), .B(new_n509_), .Z(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n499_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G229gat), .A2(G233gat), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT79), .B1(new_n514_), .B2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n512_), .B(new_n499_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n516_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT79), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n511_), .A2(new_n513_), .A3(new_n520_), .A4(new_n515_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n517_), .A2(new_n519_), .A3(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G113gat), .B(G141gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT80), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT81), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G169gat), .B(G197gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n525_), .B(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n522_), .A2(new_n528_), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n517_), .A2(new_n519_), .A3(new_n521_), .A4(new_n527_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n492_), .A2(new_n532_), .ZN(new_n533_));
  AND2_X1   g332(.A1(new_n403_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G232gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT34), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n536_), .A2(KEYINPUT35), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n501_), .A2(new_n502_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n476_), .A2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n537_), .B1(new_n539_), .B2(KEYINPUT73), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n476_), .A2(new_n538_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n476_), .A2(new_n499_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n536_), .A2(KEYINPUT35), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n540_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n541_), .A2(KEYINPUT73), .A3(new_n537_), .A4(new_n542_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G190gat), .B(G218gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G134gat), .B(G162gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n550_), .A2(KEYINPUT36), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n547_), .A2(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n550_), .B(KEYINPUT36), .Z(new_n553_));
  NAND3_X1  g352(.A1(new_n545_), .A2(new_n546_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT37), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n554_), .B2(KEYINPUT74), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n555_), .A2(new_n557_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n552_), .B(new_n554_), .C1(KEYINPUT74), .C2(new_n556_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT78), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G231gat), .A2(G233gat), .ZN(new_n563_));
  XOR2_X1   g362(.A(new_n411_), .B(new_n563_), .Z(new_n564_));
  OR2_X1    g363(.A1(new_n564_), .A2(new_n512_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n512_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(G127gat), .B(G155gat), .Z(new_n568_));
  XNOR2_X1  g367(.A(G183gat), .B(G211gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n567_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT77), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n565_), .B(new_n566_), .C1(new_n573_), .C2(new_n572_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n576_), .B1(new_n575_), .B2(new_n577_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n562_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n575_), .A2(new_n577_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT77), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(KEYINPUT78), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n561_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n534_), .A2(KEYINPUT99), .A3(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n403_), .A2(new_n587_), .A3(new_n533_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT99), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n358_), .A2(G1gat), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n588_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n593_), .A2(KEYINPUT100), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(KEYINPUT100), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(KEYINPUT38), .A3(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n403_), .A2(new_n555_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n582_), .A2(new_n583_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n492_), .A2(new_n598_), .A3(new_n532_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(G1gat), .B1(new_n600_), .B2(new_n358_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n596_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT38), .B1(new_n594_), .B2(new_n595_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n602_), .A2(new_n603_), .ZN(G1324gat));
  XNOR2_X1  g403(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(G8gat), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n588_), .A2(new_n607_), .A3(new_n284_), .A4(new_n591_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT101), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n403_), .A2(new_n555_), .A3(new_n284_), .A4(new_n599_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(G8gat), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n611_), .A2(KEYINPUT102), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(KEYINPUT102), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(KEYINPUT39), .A3(new_n613_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n613_), .A2(KEYINPUT39), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n606_), .B1(new_n609_), .B2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n608_), .B(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n619_), .A2(new_n615_), .A3(new_n614_), .A4(new_n605_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n617_), .A2(new_n620_), .ZN(G1325gat));
  AND2_X1   g420(.A1(new_n588_), .A2(new_n591_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n366_), .A3(new_n402_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n623_), .A2(KEYINPUT104), .ZN(new_n624_));
  OAI21_X1  g423(.A(G15gat), .B1(new_n600_), .B2(new_n370_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT41), .Z(new_n626_));
  NAND2_X1  g425(.A1(new_n623_), .A2(KEYINPUT104), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n624_), .A2(new_n626_), .A3(new_n627_), .ZN(G1326gat));
  OAI21_X1  g427(.A(G22gat), .B1(new_n600_), .B2(new_n327_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT42), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n622_), .A2(new_n505_), .A3(new_n328_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(G1327gat));
  NAND2_X1  g431(.A1(new_n403_), .A2(new_n561_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT43), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n403_), .A2(KEYINPUT43), .A3(new_n561_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n635_), .A2(new_n586_), .A3(new_n533_), .A4(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT44), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n585_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n640_), .A2(KEYINPUT44), .A3(new_n533_), .A4(new_n636_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n359_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(G29gat), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n585_), .A2(new_n555_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n534_), .A2(KEYINPUT105), .A3(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n403_), .A2(new_n533_), .A3(new_n645_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n358_), .A2(G29gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT106), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n644_), .A2(new_n653_), .ZN(G1328gat));
  NAND3_X1  g453(.A1(new_n639_), .A2(new_n284_), .A3(new_n641_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(G36gat), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT107), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n284_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n284_), .A2(new_n657_), .ZN(new_n659_));
  AOI21_X1  g458(.A(G36gat), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n646_), .A2(new_n649_), .A3(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT45), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n656_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT46), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n656_), .A2(new_n662_), .A3(KEYINPUT46), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(G1329gat));
  NAND2_X1  g466(.A1(new_n650_), .A2(new_n402_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(new_n361_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n639_), .A2(G43gat), .A3(new_n402_), .A4(new_n641_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1330gat));
  AOI21_X1  g473(.A(G50gat), .B1(new_n650_), .B2(new_n328_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n328_), .A2(G50gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n642_), .B2(new_n676_), .ZN(G1331gat));
  NOR2_X1   g476(.A1(new_n491_), .A2(new_n531_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n403_), .A2(new_n678_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n679_), .A2(new_n587_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(new_n359_), .ZN(new_n681_));
  INV_X1    g480(.A(G57gat), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n683_), .A2(KEYINPUT109), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(KEYINPUT109), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n597_), .A2(new_n585_), .A3(new_n678_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n358_), .A2(new_n682_), .ZN(new_n687_));
  AOI22_X1  g486(.A1(new_n684_), .A2(new_n685_), .B1(new_n686_), .B2(new_n687_), .ZN(G1332gat));
  INV_X1    g487(.A(G64gat), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n658_), .A2(new_n659_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n686_), .B2(new_n690_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(KEYINPUT48), .Z(new_n692_));
  NAND3_X1  g491(.A1(new_n680_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1333gat));
  INV_X1    g493(.A(G71gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n686_), .B2(new_n402_), .ZN(new_n696_));
  XOR2_X1   g495(.A(new_n696_), .B(KEYINPUT49), .Z(new_n697_));
  NAND3_X1  g496(.A1(new_n680_), .A2(new_n695_), .A3(new_n402_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(G1334gat));
  INV_X1    g498(.A(G78gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n686_), .B2(new_n328_), .ZN(new_n701_));
  XOR2_X1   g500(.A(new_n701_), .B(KEYINPUT50), .Z(new_n702_));
  NOR2_X1   g501(.A1(new_n327_), .A2(G78gat), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n703_), .B(KEYINPUT110), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n680_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n702_), .A2(new_n705_), .ZN(G1335gat));
  AND2_X1   g505(.A1(new_n679_), .A2(new_n645_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(new_n439_), .A3(new_n359_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n640_), .A2(new_n636_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(new_n678_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT111), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n709_), .A2(KEYINPUT111), .A3(new_n678_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n712_), .A2(new_n359_), .A3(new_n713_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n708_), .B1(new_n714_), .B2(new_n439_), .ZN(G1336gat));
  NAND3_X1  g514(.A1(new_n707_), .A2(new_n437_), .A3(new_n284_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n712_), .A2(new_n690_), .A3(new_n713_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n716_), .B1(new_n717_), .B2(new_n437_), .ZN(G1337gat));
  NAND4_X1  g517(.A1(new_n640_), .A2(new_n402_), .A3(new_n636_), .A4(new_n678_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n402_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n720_));
  AOI22_X1  g519(.A1(new_n719_), .A2(G99gat), .B1(new_n707_), .B2(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n723_), .B(new_n724_), .ZN(G1338gat));
  NAND3_X1  g524(.A1(new_n707_), .A2(new_n415_), .A3(new_n328_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n640_), .A2(new_n328_), .A3(new_n636_), .A4(new_n678_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n727_), .A2(G106gat), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n727_), .B2(G106gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n726_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g531(.A(new_n531_), .B1(new_n580_), .B2(new_n584_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT114), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n491_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n560_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n491_), .B2(new_n733_), .ZN(new_n737_));
  OAI21_X1  g536(.A(KEYINPUT54), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n737_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT54), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n560_), .A4(new_n735_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n738_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n555_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n527_), .B1(new_n515_), .B2(new_n518_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n515_), .B2(new_n514_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n745_), .A2(new_n530_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n490_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n531_), .A2(new_n489_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n467_), .A2(new_n471_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n479_), .A2(new_n468_), .A3(new_n455_), .ZN(new_n751_));
  AOI22_X1  g550(.A1(new_n750_), .A2(KEYINPUT55), .B1(new_n751_), .B2(new_n473_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n472_), .A2(new_n753_), .A3(new_n480_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(KEYINPUT56), .B1(new_n755_), .B2(new_n486_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT56), .ZN(new_n757_));
  AOI211_X1 g556(.A(new_n757_), .B(new_n488_), .C1(new_n752_), .C2(new_n754_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n749_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n748_), .B1(new_n759_), .B2(KEYINPUT115), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT115), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n749_), .B(new_n761_), .C1(new_n756_), .C2(new_n758_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n743_), .B1(new_n760_), .B2(new_n762_), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n472_), .A2(new_n753_), .A3(new_n480_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n477_), .A2(new_n479_), .A3(KEYINPUT55), .A4(new_n455_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n751_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n470_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n486_), .B1(new_n764_), .B2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(KEYINPUT117), .A3(new_n757_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n488_), .B1(new_n752_), .B2(new_n754_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(KEYINPUT56), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(KEYINPUT56), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n769_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  AND2_X1   g573(.A1(new_n746_), .A2(new_n489_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT58), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n560_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n774_), .A2(KEYINPUT58), .A3(new_n775_), .ZN(new_n779_));
  AOI22_X1  g578(.A1(KEYINPUT57), .A2(new_n763_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n759_), .A2(KEYINPUT115), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n762_), .A3(new_n747_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n555_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n783_), .A2(KEYINPUT116), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT116), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n786_), .B1(new_n763_), .B2(KEYINPUT57), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n780_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n742_), .B1(new_n788_), .B2(new_n598_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n329_), .A2(new_n359_), .A3(new_n402_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n790_), .A2(KEYINPUT118), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n794_), .B1(new_n789_), .B2(new_n791_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(G113gat), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n797_), .A3(new_n531_), .ZN(new_n798_));
  XOR2_X1   g597(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n799_));
  NOR2_X1   g598(.A1(new_n791_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n738_), .A2(new_n741_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n783_), .A2(new_n784_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n585_), .B1(new_n780_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT120), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n801_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n778_), .A2(new_n779_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n782_), .A2(KEYINPUT57), .A3(new_n555_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n763_), .A2(KEYINPUT57), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n804_), .B(new_n586_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n800_), .B1(new_n805_), .B2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT59), .B1(new_n789_), .B2(new_n791_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  AND2_X1   g613(.A1(new_n814_), .A2(new_n531_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n798_), .B1(new_n815_), .B2(new_n797_), .ZN(G1340gat));
  NAND3_X1  g615(.A1(new_n812_), .A2(new_n492_), .A3(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(G120gat), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n491_), .A2(KEYINPUT60), .ZN(new_n819_));
  MUX2_X1   g618(.A(new_n819_), .B(KEYINPUT60), .S(G120gat), .Z(new_n820_));
  NAND3_X1  g619(.A1(new_n793_), .A2(new_n795_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n818_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT121), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n818_), .A2(new_n824_), .A3(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n825_), .ZN(G1341gat));
  INV_X1    g625(.A(G127gat), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n796_), .A2(new_n827_), .A3(new_n585_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n598_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n814_), .A2(new_n829_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n828_), .B1(new_n830_), .B2(new_n827_), .ZN(G1342gat));
  AOI21_X1  g630(.A(G134gat), .B1(new_n796_), .B2(new_n743_), .ZN(new_n832_));
  XOR2_X1   g631(.A(KEYINPUT122), .B(G134gat), .Z(new_n833_));
  NAND2_X1  g632(.A1(new_n561_), .A2(new_n833_), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT123), .Z(new_n835_));
  AOI21_X1  g634(.A(new_n832_), .B1(new_n814_), .B2(new_n835_), .ZN(G1343gat));
  NOR2_X1   g635(.A1(new_n789_), .A2(new_n402_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n690_), .A2(new_n358_), .A3(new_n327_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n839_), .A2(new_n532_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(new_n288_), .ZN(G1344gat));
  NOR2_X1   g640(.A1(new_n839_), .A2(new_n491_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(new_n289_), .ZN(G1345gat));
  NOR2_X1   g642(.A1(new_n839_), .A2(new_n586_), .ZN(new_n844_));
  XOR2_X1   g643(.A(KEYINPUT61), .B(G155gat), .Z(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1346gat));
  INV_X1    g645(.A(G162gat), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n837_), .A2(new_n847_), .A3(new_n743_), .A4(new_n838_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n839_), .A2(new_n560_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n847_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  OAI211_X1 g651(.A(KEYINPUT124), .B(new_n848_), .C1(new_n849_), .C2(new_n847_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1347gat));
  OAI21_X1  g653(.A(new_n586_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT120), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n856_), .A2(new_n801_), .A3(new_n810_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT22), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n690_), .A2(new_n371_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n859_), .A2(new_n328_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n857_), .A2(new_n858_), .A3(new_n531_), .A4(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT62), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n862_), .A2(G169gat), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n857_), .A2(new_n860_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n864_), .A2(KEYINPUT62), .A3(new_n532_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n225_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n863_), .B1(new_n866_), .B2(new_n862_), .ZN(G1348gat));
  INV_X1    g666(.A(new_n864_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G176gat), .B1(new_n868_), .B2(new_n492_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n789_), .A2(new_n328_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n859_), .A2(new_n226_), .A3(new_n491_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n869_), .B1(new_n870_), .B2(new_n871_), .ZN(G1349gat));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n868_), .A2(new_n873_), .A3(new_n829_), .A4(new_n253_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n870_), .A2(new_n585_), .A3(new_n371_), .A4(new_n690_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n214_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n829_), .A2(new_n253_), .ZN(new_n877_));
  OAI21_X1  g676(.A(KEYINPUT125), .B1(new_n864_), .B2(new_n877_), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n874_), .A2(new_n876_), .A3(new_n878_), .ZN(G1350gat));
  OAI21_X1  g678(.A(G190gat), .B1(new_n864_), .B2(new_n560_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n555_), .A2(new_n252_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n864_), .B2(new_n881_), .ZN(G1351gat));
  NOR2_X1   g681(.A1(new_n359_), .A2(new_n327_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n690_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n837_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT126), .ZN(new_n887_));
  NOR4_X1   g686(.A1(new_n789_), .A2(KEYINPUT126), .A3(new_n402_), .A4(new_n884_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(G197gat), .B1(new_n890_), .B2(new_n531_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n837_), .B2(new_n885_), .ZN(new_n893_));
  OAI211_X1 g692(.A(G197gat), .B(new_n531_), .C1(new_n893_), .C2(new_n888_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n891_), .A2(new_n895_), .ZN(G1352gat));
  OAI21_X1  g695(.A(new_n492_), .B1(new_n893_), .B2(new_n888_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(KEYINPUT127), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n598_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n900_), .B1(new_n890_), .B2(new_n901_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n901_), .B(new_n900_), .C1(new_n893_), .C2(new_n888_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n902_), .A2(new_n904_), .ZN(G1354gat));
  INV_X1    g704(.A(G218gat), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n890_), .A2(new_n906_), .A3(new_n743_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n560_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n906_), .B2(new_n908_), .ZN(G1355gat));
endmodule


