//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n772_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n908_, new_n909_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT75), .B(G8gat), .Z(new_n203_));
  INV_X1    g002(.A(G1gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n202_), .B1(new_n205_), .B2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n209_), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n202_), .B(new_n208_), .C1(new_n205_), .C2(new_n206_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G231gat), .A2(G233gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G57gat), .B(G64gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT11), .ZN(new_n216_));
  XOR2_X1   g015(.A(G71gat), .B(G78gat), .Z(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n217_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n215_), .A2(KEYINPUT11), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n214_), .B(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n224_), .A2(KEYINPUT76), .ZN(new_n225_));
  XOR2_X1   g024(.A(G127gat), .B(G155gat), .Z(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT16), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G183gat), .B(G211gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(KEYINPUT76), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n225_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT77), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n224_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n224_), .A2(new_n234_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n229_), .B(KEYINPUT17), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT36), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G232gat), .A2(G233gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT34), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G85gat), .A2(G92gat), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT66), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G85gat), .A2(G92gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n247_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT66), .B1(new_n249_), .B2(new_n244_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT7), .ZN(new_n252_));
  INV_X1    g051(.A(G99gat), .ZN(new_n253_));
  INV_X1    g052(.A(G106gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT65), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT65), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n257_), .A2(new_n252_), .A3(new_n253_), .A4(new_n254_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT64), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT64), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n261_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n256_), .A2(new_n258_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G99gat), .A2(G106gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT67), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n266_), .A2(KEYINPUT6), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT6), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n268_), .A2(KEYINPUT67), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n265_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(KEYINPUT67), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n266_), .A2(KEYINPUT6), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(new_n264_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n251_), .B1(new_n263_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT8), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n256_), .A2(new_n258_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n264_), .B(KEYINPUT6), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n260_), .A2(new_n262_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n248_), .A2(new_n250_), .A3(new_n276_), .ZN(new_n281_));
  OAI22_X1  g080(.A1(new_n275_), .A2(new_n276_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G29gat), .B(G36gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G43gat), .B(G50gat), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G43gat), .B(G50gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n283_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n245_), .A2(KEYINPUT9), .A3(new_n247_), .ZN(new_n290_));
  AND2_X1   g089(.A1(new_n278_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(KEYINPUT10), .B(G99gat), .Z(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OAI221_X1 g092(.A(new_n291_), .B1(KEYINPUT9), .B2(new_n247_), .C1(G106gat), .C2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n282_), .A2(new_n289_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AND2_X1   g095(.A1(new_n286_), .A2(new_n288_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT15), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT15), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n289_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n301_), .B1(new_n294_), .B2(new_n282_), .ZN(new_n302_));
  OAI211_X1 g101(.A(KEYINPUT35), .B(new_n243_), .C1(new_n296_), .C2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n282_), .A2(new_n294_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n243_), .A2(KEYINPUT35), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n243_), .A2(KEYINPUT35), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .A4(new_n295_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n303_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G190gat), .B(G218gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT73), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G134gat), .B(G162gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  OAI21_X1  g112(.A(new_n241_), .B1(new_n309_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n303_), .A2(new_n308_), .A3(KEYINPUT74), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n313_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n315_), .A2(new_n241_), .A3(new_n313_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n322_));
  OAI21_X1  g121(.A(G228gat), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G211gat), .B(G218gat), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT88), .B(G197gat), .ZN(new_n327_));
  INV_X1    g126(.A(G204gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT21), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n330_), .B1(G197gat), .B2(G204gat), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n326_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(G197gat), .A2(G204gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n330_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(G197gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(KEYINPUT88), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT88), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(G197gat), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n328_), .B1(new_n339_), .B2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT89), .B1(new_n342_), .B2(new_n333_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT89), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n344_), .B(new_n334_), .C1(new_n327_), .C2(new_n328_), .ZN(new_n345_));
  INV_X1    g144(.A(G211gat), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n346_), .A2(G218gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(G218gat), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT21), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n343_), .A2(new_n345_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT90), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n349_), .B1(new_n335_), .B2(KEYINPUT89), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(KEYINPUT90), .A3(new_n345_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n337_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n358_), .A2(KEYINPUT84), .A3(G155gat), .A4(G162gat), .ZN(new_n359_));
  INV_X1    g158(.A(G141gat), .ZN(new_n360_));
  INV_X1    g159(.A(G148gat), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n359_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT1), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n358_), .A2(G155gat), .A3(G162gat), .ZN(new_n367_));
  OR2_X1    g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT84), .ZN(new_n369_));
  NAND4_X1  g168(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .A4(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n364_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT85), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT85), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n364_), .A2(new_n370_), .A3(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n363_), .A2(KEYINPUT86), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT2), .ZN(new_n377_));
  OR3_X1    g176(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n362_), .A2(KEYINPUT3), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n377_), .A2(new_n378_), .A3(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n376_), .A2(KEYINPUT2), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n365_), .B(new_n368_), .C1(new_n380_), .C2(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n357_), .B1(new_n375_), .B2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n324_), .B1(new_n356_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n332_), .A2(new_n336_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT90), .B1(new_n354_), .B2(new_n345_), .ZN(new_n386_));
  AND4_X1   g185(.A1(KEYINPUT90), .A2(new_n343_), .A3(new_n345_), .A4(new_n350_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n385_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n374_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n373_), .B1(new_n364_), .B2(new_n370_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n382_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT29), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n388_), .A2(new_n392_), .A3(new_n323_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n384_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT92), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n394_), .A2(new_n395_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n396_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n384_), .A2(new_n393_), .A3(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT28), .B1(new_n391_), .B2(KEYINPUT29), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT28), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n375_), .A2(new_n401_), .A3(new_n357_), .A4(new_n382_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G22gat), .B(G50gat), .ZN(new_n403_));
  AND3_X1   g202(.A1(new_n400_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n403_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n397_), .A2(new_n399_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n395_), .B1(new_n394_), .B2(new_n396_), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT93), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n406_), .A2(new_n399_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n408_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT93), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n410_), .A2(new_n411_), .A3(new_n412_), .A4(new_n397_), .ZN(new_n413_));
  OR3_X1    g212(.A1(new_n394_), .A2(KEYINPUT91), .A3(new_n396_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n406_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n394_), .A2(new_n396_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(KEYINPUT91), .A3(new_n399_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n409_), .A2(new_n413_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420_));
  XOR2_X1   g219(.A(G127gat), .B(G134gat), .Z(new_n421_));
  XOR2_X1   g220(.A(G113gat), .B(G120gat), .Z(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n391_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n375_), .A2(new_n382_), .A3(new_n423_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(KEYINPUT4), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n391_), .A2(new_n428_), .A3(new_n424_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n420_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n425_), .A2(new_n426_), .B1(G225gat), .B2(G233gat), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G1gat), .B(G29gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(G85gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT0), .B(G57gat), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n434_), .B(new_n435_), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n432_), .A2(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n430_), .A2(new_n436_), .A3(new_n431_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G169gat), .A2(G176gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT80), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT80), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(G169gat), .A3(G176gat), .ZN(new_n445_));
  INV_X1    g244(.A(G169gat), .ZN(new_n446_));
  INV_X1    g245(.A(G176gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n443_), .A2(new_n445_), .A3(new_n448_), .A4(KEYINPUT24), .ZN(new_n449_));
  OR2_X1    g248(.A1(new_n448_), .A2(KEYINPUT24), .ZN(new_n450_));
  INV_X1    g249(.A(G183gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT25), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT25), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G183gat), .ZN(new_n454_));
  INV_X1    g253(.A(G190gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT26), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT26), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(G190gat), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n452_), .A2(new_n454_), .A3(new_n456_), .A4(new_n458_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n449_), .A2(new_n450_), .A3(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT23), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(G183gat), .A3(G190gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT81), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n463_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT23), .B1(new_n451_), .B2(new_n455_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n464_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n443_), .A2(new_n445_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT82), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n446_), .A2(KEYINPUT22), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n446_), .A2(KEYINPUT22), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n446_), .A2(KEYINPUT22), .ZN(new_n473_));
  AOI21_X1  g272(.A(G176gat), .B1(new_n473_), .B2(KEYINPUT82), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n468_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n466_), .A2(KEYINPUT83), .A3(new_n462_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n451_), .A2(new_n455_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT83), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n478_), .A2(new_n461_), .A3(G183gat), .A4(G190gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n476_), .A2(new_n477_), .A3(new_n479_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n460_), .A2(new_n467_), .B1(new_n475_), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G71gat), .B(G99gat), .ZN(new_n482_));
  INV_X1    g281(.A(G43gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n481_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(new_n424_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G227gat), .A2(G233gat), .ZN(new_n487_));
  INV_X1    g286(.A(G15gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT30), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT31), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n486_), .B(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n441_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT102), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT101), .ZN(new_n495_));
  XOR2_X1   g294(.A(G8gat), .B(G36gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G64gat), .B(G92gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(KEYINPUT19), .A2(G226gat), .A3(G233gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT19), .B1(G226gat), .B2(G233gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n505_), .B(KEYINPUT94), .Z(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n450_), .A2(new_n459_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n448_), .A2(KEYINPUT24), .A3(new_n442_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n476_), .A2(new_n479_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n467_), .A2(new_n477_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n470_), .A2(new_n471_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n468_), .B1(new_n514_), .B2(new_n447_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n510_), .A2(new_n512_), .B1(new_n513_), .B2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT96), .B1(new_n356_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT96), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n513_), .A2(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n508_), .A2(new_n509_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n519_), .B1(new_n520_), .B2(new_n511_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n388_), .A2(new_n518_), .A3(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n385_), .B(new_n481_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT20), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT95), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n524_), .A2(new_n527_), .A3(KEYINPUT20), .ZN(new_n528_));
  AND4_X1   g327(.A1(new_n507_), .A2(new_n523_), .A3(new_n526_), .A4(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n505_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n388_), .A2(new_n521_), .ZN(new_n531_));
  XOR2_X1   g330(.A(KEYINPUT100), .B(KEYINPUT20), .Z(new_n532_));
  NOR2_X1   g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT97), .B1(new_n356_), .B2(new_n481_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT97), .ZN(new_n535_));
  INV_X1    g334(.A(new_n481_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n388_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n534_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n530_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n501_), .B1(new_n529_), .B2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n523_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n506_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n531_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n538_), .A2(KEYINPUT20), .A3(new_n530_), .A4(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n500_), .A3(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n540_), .A2(new_n545_), .A3(KEYINPUT27), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n524_), .A2(new_n527_), .A3(KEYINPUT20), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n527_), .B1(new_n524_), .B2(KEYINPUT20), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n507_), .B1(new_n549_), .B2(new_n523_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n530_), .A2(KEYINPUT20), .ZN(new_n551_));
  AOI211_X1 g350(.A(new_n551_), .B(new_n531_), .C1(new_n534_), .C2(new_n537_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n501_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n545_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT27), .ZN(new_n555_));
  AOI22_X1  g354(.A1(new_n495_), .A2(new_n546_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n540_), .A2(new_n545_), .A3(KEYINPUT101), .A4(KEYINPUT27), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n494_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n546_), .A2(new_n495_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n545_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n500_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n555_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  AND4_X1   g361(.A1(new_n494_), .A2(new_n559_), .A3(new_n557_), .A4(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n419_), .B(new_n493_), .C1(new_n558_), .C2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT33), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n565_), .B1(new_n432_), .B2(new_n437_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n425_), .A2(new_n426_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT99), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n420_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n569_), .B1(new_n568_), .B2(new_n567_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n427_), .A2(new_n420_), .A3(new_n429_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n437_), .A3(new_n571_), .ZN(new_n572_));
  OAI211_X1 g371(.A(KEYINPUT33), .B(new_n436_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n566_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n560_), .A2(new_n574_), .A3(new_n561_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n500_), .A2(KEYINPUT32), .ZN(new_n576_));
  AND3_X1   g375(.A1(new_n542_), .A2(new_n544_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n533_), .A2(new_n538_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n505_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n523_), .A2(new_n526_), .A3(new_n507_), .A4(new_n528_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n576_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n577_), .A2(new_n440_), .A3(new_n581_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n419_), .B1(new_n575_), .B2(new_n582_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n559_), .A2(new_n562_), .A3(new_n557_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n409_), .A2(new_n413_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n416_), .A2(new_n418_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n440_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n583_), .B1(new_n584_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(new_n492_), .ZN(new_n590_));
  AOI211_X1 g389(.A(new_n240_), .B(new_n319_), .C1(new_n564_), .C2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G230gat), .A2(G233gat), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n282_), .A2(new_n294_), .A3(new_n222_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(KEYINPUT68), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT68), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n282_), .A2(new_n596_), .A3(new_n294_), .A4(new_n222_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n222_), .B1(new_n282_), .B2(new_n294_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n593_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n594_), .A2(new_n592_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT69), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT12), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n304_), .B2(new_n223_), .ZN(new_n604_));
  XOR2_X1   g403(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n605_));
  AOI211_X1 g404(.A(new_n222_), .B(new_n605_), .C1(new_n282_), .C2(new_n294_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n601_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n600_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(G120gat), .B(G148gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(G176gat), .B(G204gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT71), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n608_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n600_), .A2(new_n607_), .A3(new_n613_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT13), .ZN(new_n618_));
  OAI211_X1 g417(.A(new_n616_), .B(new_n617_), .C1(KEYINPUT72), .C2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n616_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n617_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n619_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT79), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G229gat), .A2(G233gat), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n210_), .A2(new_n297_), .A3(new_n211_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n297_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n627_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n212_), .A2(new_n289_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n298_), .A2(new_n210_), .A3(new_n211_), .A4(new_n300_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n626_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n630_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G113gat), .B(G141gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G169gat), .B(G197gat), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n635_), .B(new_n636_), .Z(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n625_), .B1(new_n634_), .B2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n630_), .A2(new_n633_), .A3(KEYINPUT79), .A4(new_n637_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n634_), .A2(new_n638_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n624_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT103), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n591_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n440_), .ZN(new_n648_));
  OR2_X1    g447(.A1(new_n319_), .A2(KEYINPUT37), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n319_), .A2(KEYINPUT37), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n624_), .A2(new_n649_), .A3(new_n239_), .A4(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT78), .Z(new_n652_));
  INV_X1    g451(.A(new_n643_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n564_), .B2(new_n590_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n655_), .A2(new_n204_), .A3(new_n441_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT38), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n657_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n648_), .A2(new_n658_), .A3(new_n659_), .ZN(G1324gat));
  NOR2_X1   g459(.A1(new_n558_), .A2(new_n563_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n655_), .A2(new_n203_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n661_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G8gat), .B1(new_n647_), .B2(new_n663_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n664_), .A2(KEYINPUT39), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(KEYINPUT39), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n662_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI211_X1 g468(.A(KEYINPUT40), .B(new_n662_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1325gat));
  OAI21_X1  g470(.A(G15gat), .B1(new_n647_), .B2(new_n492_), .ZN(new_n672_));
  XOR2_X1   g471(.A(KEYINPUT104), .B(KEYINPUT41), .Z(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT105), .ZN(new_n674_));
  OR2_X1    g473(.A1(new_n672_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(new_n674_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n492_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n655_), .A2(new_n488_), .A3(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n675_), .A2(new_n676_), .A3(new_n678_), .ZN(G1326gat));
  INV_X1    g478(.A(G22gat), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n680_), .B1(new_n646_), .B2(new_n587_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(KEYINPUT106), .B(KEYINPUT42), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n655_), .A2(new_n680_), .A3(new_n587_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1327gat));
  AND2_X1   g484(.A1(new_n645_), .A2(new_n240_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n564_), .A2(new_n590_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n649_), .A2(new_n650_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n687_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n689_), .ZN(new_n691_));
  AOI211_X1 g490(.A(KEYINPUT43), .B(new_n691_), .C1(new_n564_), .C2(new_n590_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n686_), .B1(new_n690_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  OAI211_X1 g494(.A(KEYINPUT44), .B(new_n686_), .C1(new_n690_), .C2(new_n692_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G29gat), .B1(new_n697_), .B2(new_n440_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n240_), .A2(new_n319_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n624_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n654_), .A2(new_n701_), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n440_), .A2(G29gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n698_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(G1328gat));
  NAND3_X1  g505(.A1(new_n695_), .A2(new_n661_), .A3(new_n696_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(KEYINPUT108), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n695_), .A2(new_n709_), .A3(new_n661_), .A4(new_n696_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n708_), .A2(G36gat), .A3(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n702_), .ZN(new_n712_));
  OR2_X1    g511(.A1(new_n661_), .A2(KEYINPUT109), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n661_), .A2(KEYINPUT109), .ZN(new_n714_));
  AOI21_X1  g513(.A(G36gat), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT110), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n712_), .A2(new_n718_), .A3(new_n715_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n717_), .A2(KEYINPUT45), .A3(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT45), .B1(new_n717_), .B2(new_n719_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n711_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT46), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n711_), .A2(KEYINPUT46), .A3(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1329gat));
  OAI21_X1  g526(.A(G43gat), .B1(new_n697_), .B2(new_n492_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n677_), .A2(new_n483_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n728_), .B1(new_n702_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT47), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n730_), .B(new_n731_), .ZN(G1330gat));
  INV_X1    g531(.A(G50gat), .ZN(new_n733_));
  NOR3_X1   g532(.A1(new_n697_), .A2(new_n733_), .A3(new_n419_), .ZN(new_n734_));
  AOI21_X1  g533(.A(G50gat), .B1(new_n712_), .B2(new_n587_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1331gat));
  AOI21_X1  g535(.A(new_n643_), .B1(new_n564_), .B2(new_n590_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n649_), .A2(new_n239_), .A3(new_n650_), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(new_n700_), .A3(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(G57gat), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(new_n441_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n591_), .A2(new_n653_), .A3(new_n700_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n742_), .A2(new_n441_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n741_), .B1(new_n743_), .B2(new_n740_), .ZN(G1332gat));
  INV_X1    g543(.A(G64gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n713_), .A2(new_n714_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n742_), .B2(new_n746_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n747_), .B(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n739_), .A2(new_n745_), .A3(new_n746_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1333gat));
  INV_X1    g550(.A(G71gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n742_), .B2(new_n677_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n739_), .A2(new_n752_), .A3(new_n677_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(G1334gat));
  INV_X1    g556(.A(G78gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n742_), .B2(new_n587_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT50), .Z(new_n760_));
  NAND3_X1  g559(.A1(new_n739_), .A2(new_n758_), .A3(new_n587_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1335gat));
  OR2_X1    g561(.A1(new_n690_), .A2(new_n692_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n624_), .A2(new_n239_), .A3(new_n643_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(G85gat), .B1(new_n766_), .B2(new_n440_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n699_), .A2(new_n624_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n737_), .A2(new_n768_), .ZN(new_n769_));
  OR3_X1    g568(.A1(new_n769_), .A2(G85gat), .A3(new_n440_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(new_n770_), .ZN(G1336gat));
  INV_X1    g570(.A(new_n746_), .ZN(new_n772_));
  OAI21_X1  g571(.A(G92gat), .B1(new_n766_), .B2(new_n772_), .ZN(new_n773_));
  OR3_X1    g572(.A1(new_n769_), .A2(G92gat), .A3(new_n663_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(G1337gat));
  NOR3_X1   g574(.A1(new_n769_), .A2(new_n492_), .A3(new_n293_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n765_), .A2(new_n677_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(G99gat), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT51), .Z(G1338gat));
  NAND4_X1  g578(.A1(new_n737_), .A2(new_n254_), .A3(new_n587_), .A4(new_n768_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n587_), .B(new_n764_), .C1(new_n690_), .C2(new_n692_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(G106gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT114), .B1(new_n782_), .B2(KEYINPUT52), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT114), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT52), .ZN(new_n785_));
  AOI211_X1 g584(.A(new_n784_), .B(new_n785_), .C1(new_n781_), .C2(G106gat), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n783_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n782_), .B2(KEYINPUT52), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n781_), .A2(KEYINPUT113), .A3(new_n785_), .A4(G106gat), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n780_), .B1(new_n787_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(KEYINPUT53), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(new_n780_), .C1(new_n787_), .C2(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n793_), .A2(new_n795_), .ZN(G1339gat));
  INV_X1    g595(.A(KEYINPUT116), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n651_), .A2(new_n643_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n797_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n738_), .A2(new_n799_), .A3(new_n653_), .A4(new_n624_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n798_), .A2(KEYINPUT115), .A3(new_n799_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT116), .B(KEYINPUT54), .C1(new_n651_), .C2(new_n643_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n800_), .A2(new_n803_), .A3(new_n804_), .A4(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n631_), .A2(new_n632_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n626_), .B1(new_n808_), .B2(KEYINPUT118), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(KEYINPUT118), .B2(new_n808_), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n628_), .A2(new_n629_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n637_), .B1(new_n811_), .B2(new_n626_), .ZN(new_n812_));
  AOI22_X1  g611(.A1(new_n639_), .A2(new_n640_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n814_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n604_), .A2(new_n606_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n593_), .B1(new_n816_), .B2(new_n598_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n607_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n601_), .B(KEYINPUT55), .C1(new_n604_), .C2(new_n606_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n615_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT56), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT117), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n615_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n643_), .A2(new_n617_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT56), .B1(new_n821_), .B2(new_n615_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(KEYINPUT117), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n815_), .B1(new_n827_), .B2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n319_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n813_), .A2(new_n617_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n650_), .A2(new_n649_), .B1(new_n834_), .B2(KEYINPUT58), .ZN(new_n835_));
  OR2_X1    g634(.A1(new_n834_), .A2(KEYINPUT58), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n832_), .A2(KEYINPUT57), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n815_), .ZN(new_n838_));
  AND3_X1   g637(.A1(new_n821_), .A2(KEYINPUT56), .A3(new_n615_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n839_), .A2(new_n829_), .A3(KEYINPUT117), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n822_), .A2(KEYINPUT117), .A3(new_n823_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n828_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n838_), .B1(new_n840_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n319_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT119), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(KEYINPUT119), .B(new_n847_), .C1(new_n831_), .C2(new_n319_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n837_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n239_), .B1(new_n851_), .B2(KEYINPUT120), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n837_), .B(new_n853_), .C1(new_n848_), .C2(new_n850_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n807_), .B1(new_n852_), .B2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n663_), .A2(new_n419_), .A3(new_n441_), .A4(new_n677_), .ZN(new_n856_));
  OAI21_X1  g655(.A(KEYINPUT59), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(KEYINPUT59), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n846_), .A2(new_n847_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n239_), .B1(new_n837_), .B2(new_n859_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n858_), .B1(new_n807_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n857_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n643_), .A2(G113gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT123), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n862_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n851_), .A2(KEYINPUT120), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n866_), .A2(new_n240_), .A3(new_n854_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n856_), .B1(new_n867_), .B2(new_n806_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT121), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(KEYINPUT121), .B1(new_n855_), .B2(new_n856_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n870_), .A2(new_n871_), .A3(new_n643_), .ZN(new_n872_));
  INV_X1    g671(.A(G113gat), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n872_), .A2(KEYINPUT122), .A3(new_n873_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n865_), .B1(new_n876_), .B2(new_n877_), .ZN(G1340gat));
  INV_X1    g677(.A(KEYINPUT124), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n862_), .B2(new_n624_), .ZN(new_n880_));
  NAND4_X1  g679(.A1(new_n857_), .A2(KEYINPUT124), .A3(new_n700_), .A4(new_n861_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(G120gat), .A3(new_n881_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n870_), .A2(new_n871_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n624_), .A2(KEYINPUT60), .ZN(new_n884_));
  MUX2_X1   g683(.A(new_n884_), .B(KEYINPUT60), .S(G120gat), .Z(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n882_), .A2(new_n886_), .ZN(G1341gat));
  INV_X1    g686(.A(G127gat), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n883_), .A2(new_n888_), .A3(new_n239_), .ZN(new_n889_));
  OAI21_X1  g688(.A(G127gat), .B1(new_n862_), .B2(new_n240_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1342gat));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n689_), .B(new_n861_), .C1(new_n868_), .C2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(G134gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n845_), .A2(G134gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n870_), .A2(new_n871_), .A3(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT125), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n894_), .A2(new_n899_), .A3(new_n896_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n900_), .ZN(G1343gat));
  NAND4_X1  g700(.A1(new_n772_), .A2(new_n587_), .A3(new_n441_), .A4(new_n492_), .ZN(new_n902_));
  OR2_X1    g701(.A1(new_n855_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n903_), .A2(new_n653_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(new_n360_), .ZN(G1344gat));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n624_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(new_n361_), .ZN(G1345gat));
  NOR2_X1   g706(.A1(new_n903_), .A2(new_n240_), .ZN(new_n908_));
  XOR2_X1   g707(.A(KEYINPUT61), .B(G155gat), .Z(new_n909_));
  XNOR2_X1  g708(.A(new_n908_), .B(new_n909_), .ZN(G1346gat));
  OAI21_X1  g709(.A(G162gat), .B1(new_n903_), .B2(new_n691_), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n845_), .A2(G162gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n911_), .B1(new_n903_), .B2(new_n912_), .ZN(G1347gat));
  NOR2_X1   g712(.A1(new_n807_), .A2(new_n860_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n746_), .A2(new_n493_), .ZN(new_n915_));
  NOR3_X1   g714(.A1(new_n914_), .A2(new_n587_), .A3(new_n915_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n446_), .B1(new_n916_), .B2(new_n643_), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n917_), .A2(KEYINPUT62), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(KEYINPUT62), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n916_), .A2(new_n643_), .A3(new_n514_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n918_), .A2(new_n919_), .A3(new_n920_), .ZN(G1348gat));
  AOI21_X1  g720(.A(G176gat), .B1(new_n916_), .B2(new_n700_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n855_), .A2(new_n587_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n915_), .A2(new_n447_), .A3(new_n624_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1349gat));
  NAND4_X1  g724(.A1(new_n923_), .A2(new_n493_), .A3(new_n239_), .A4(new_n746_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n240_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n926_), .A2(new_n451_), .B1(new_n916_), .B2(new_n927_), .ZN(G1350gat));
  NAND4_X1  g727(.A1(new_n916_), .A2(new_n456_), .A3(new_n458_), .A4(new_n319_), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n916_), .A2(new_n689_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n930_), .B2(new_n455_), .ZN(G1351gat));
  NOR4_X1   g730(.A1(new_n855_), .A2(new_n677_), .A3(new_n588_), .A4(new_n772_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n643_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n700_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n935_), .B1(new_n936_), .B2(G204gat), .ZN(new_n937_));
  XNOR2_X1  g736(.A(KEYINPUT126), .B(G204gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n935_), .B2(new_n938_), .ZN(G1353gat));
  NAND2_X1  g738(.A1(new_n932_), .A2(new_n239_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(KEYINPUT63), .B(G211gat), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n940_), .B2(new_n943_), .ZN(G1354gat));
  NAND2_X1  g743(.A1(new_n932_), .A2(new_n319_), .ZN(new_n945_));
  XOR2_X1   g744(.A(KEYINPUT127), .B(G218gat), .Z(new_n946_));
  NOR2_X1   g745(.A1(new_n691_), .A2(new_n946_), .ZN(new_n947_));
  AOI22_X1  g746(.A1(new_n945_), .A2(new_n946_), .B1(new_n932_), .B2(new_n947_), .ZN(G1355gat));
endmodule


