//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n571_, new_n572_, new_n573_, new_n574_, new_n575_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n804_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n860_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(new_n202_), .B(KEYINPUT95), .Z(new_n203_));
  INV_X1    g002(.A(KEYINPUT4), .ZN(new_n204_));
  NOR3_X1   g003(.A1(KEYINPUT84), .A2(G141gat), .A3(G148gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  OAI22_X1  g007(.A1(new_n205_), .A2(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n209_), .B1(new_n206_), .B2(new_n205_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n208_), .B(KEYINPUT82), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n210_), .B1(KEYINPUT2), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n213_), .B(KEYINPUT83), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n212_), .B(new_n214_), .C1(G155gat), .C2(G162gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(new_n214_), .B2(KEYINPUT1), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(KEYINPUT1), .B2(new_n214_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n211_), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n218_), .B(new_n219_), .C1(G141gat), .C2(G148gat), .ZN(new_n220_));
  XOR2_X1   g019(.A(G127gat), .B(G134gat), .Z(new_n221_));
  XOR2_X1   g020(.A(G113gat), .B(G120gat), .Z(new_n222_));
  OR2_X1    g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n222_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n215_), .A2(new_n220_), .A3(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT94), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n215_), .A2(new_n220_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT85), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT85), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n215_), .A2(new_n230_), .A3(new_n220_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(KEYINPUT81), .ZN(new_n232_));
  XOR2_X1   g031(.A(new_n232_), .B(new_n223_), .Z(new_n233_));
  NAND3_X1  g032(.A1(new_n229_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n204_), .B1(new_n227_), .B2(new_n234_), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n234_), .A2(new_n204_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n203_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n227_), .A2(new_n202_), .A3(new_n234_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G1gat), .B(G29gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(G85gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT0), .B(G57gat), .ZN(new_n241_));
  XOR2_X1   g040(.A(new_n240_), .B(new_n241_), .Z(new_n242_));
  NAND3_X1  g041(.A1(new_n237_), .A2(new_n238_), .A3(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT96), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT33), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n237_), .A2(KEYINPUT96), .A3(new_n238_), .A4(new_n242_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT97), .ZN(new_n249_));
  XOR2_X1   g048(.A(G8gat), .B(G36gat), .Z(new_n250_));
  XNOR2_X1  g049(.A(G64gat), .B(G92gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G211gat), .B(G218gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(G197gat), .B(G204gat), .Z(new_n256_));
  OAI21_X1  g055(.A(new_n255_), .B1(new_n256_), .B2(KEYINPUT87), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n257_), .B1(new_n256_), .B2(new_n255_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT21), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT21), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT23), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n264_), .B1(G183gat), .B2(G190gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n266_));
  OR3_X1    g065(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(G169gat), .ZN(new_n269_));
  INV_X1    g068(.A(G176gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(KEYINPUT24), .B1(new_n269_), .B2(new_n270_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n271_), .B1(new_n273_), .B2(KEYINPUT89), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(KEYINPUT89), .B2(new_n273_), .ZN(new_n275_));
  XOR2_X1   g074(.A(KEYINPUT25), .B(G183gat), .Z(new_n276_));
  XOR2_X1   g075(.A(KEYINPUT26), .B(G190gat), .Z(new_n277_));
  OAI221_X1 g076(.A(new_n264_), .B1(KEYINPUT24), .B2(new_n271_), .C1(new_n276_), .C2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n268_), .B1(new_n275_), .B2(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n262_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT20), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G226gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT19), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n273_), .A2(new_n271_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT79), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n268_), .B1(new_n287_), .B2(new_n278_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n262_), .A2(KEYINPUT90), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT90), .B1(new_n262_), .B2(new_n288_), .ZN(new_n290_));
  OAI211_X1 g089(.A(new_n282_), .B(new_n285_), .C1(new_n289_), .C2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n281_), .B1(new_n262_), .B2(new_n279_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n292_), .B1(new_n262_), .B2(new_n288_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n284_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n254_), .B1(new_n291_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT93), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  AOI211_X1 g096(.A(KEYINPUT93), .B(new_n254_), .C1(new_n291_), .C2(new_n294_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n237_), .A2(KEYINPUT33), .A3(new_n238_), .A4(new_n242_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n291_), .A2(new_n254_), .A3(new_n294_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT92), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n202_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n242_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n227_), .A2(new_n234_), .A3(new_n203_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  AND4_X1   g106(.A1(new_n300_), .A2(new_n301_), .A3(new_n303_), .A4(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT97), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n245_), .A2(new_n309_), .A3(new_n246_), .A4(new_n247_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n249_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n262_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n312_), .B1(G228gat), .B2(G233gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n229_), .A2(new_n231_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT29), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n313_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n228_), .A2(KEYINPUT29), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(new_n262_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(G228gat), .A3(G233gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G78gat), .B(G106gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT88), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n314_), .A2(new_n315_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  XOR2_X1   g127(.A(G22gat), .B(G50gat), .Z(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n314_), .A2(new_n315_), .A3(new_n326_), .ZN(new_n331_));
  AND3_X1   g130(.A1(new_n328_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n330_), .B1(new_n328_), .B2(new_n331_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n324_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n320_), .B(new_n321_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n321_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n320_), .B(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n338_), .B(new_n324_), .C1(new_n333_), .C2(new_n332_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n293_), .A2(new_n284_), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n282_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n341_), .B1(new_n342_), .B2(new_n284_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n254_), .A2(KEYINPUT32), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n345_), .A2(KEYINPUT98), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n291_), .A2(new_n294_), .A3(new_n344_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n347_), .A2(KEYINPUT98), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n237_), .A2(new_n238_), .A3(new_n242_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n242_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n350_));
  OAI221_X1 g149(.A(new_n346_), .B1(new_n345_), .B2(new_n348_), .C1(new_n349_), .C2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n311_), .A2(new_n340_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G227gat), .A2(G233gat), .ZN(new_n353_));
  INV_X1    g152(.A(G71gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G99gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n288_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(new_n233_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G15gat), .B(G43gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(KEYINPUT80), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT30), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT31), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n358_), .B(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT27), .ZN(new_n364_));
  INV_X1    g163(.A(new_n303_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n364_), .B1(new_n365_), .B2(new_n299_), .ZN(new_n366_));
  OAI211_X1 g165(.A(KEYINPUT27), .B(new_n302_), .C1(new_n343_), .C2(new_n254_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n349_), .A2(new_n350_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n366_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n336_), .A2(new_n339_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n363_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n367_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n368_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n363_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n352_), .A2(new_n371_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(G85gat), .A2(G92gat), .ZN(new_n378_));
  AND2_X1   g177(.A1(G85gat), .A2(G92gat), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n378_), .B1(new_n379_), .B2(KEYINPUT9), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT65), .B1(new_n379_), .B2(KEYINPUT9), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT65), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT9), .ZN(new_n383_));
  INV_X1    g182(.A(G85gat), .ZN(new_n384_));
  INV_X1    g183(.A(G92gat), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n382_), .B(new_n383_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n380_), .A2(new_n381_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G99gat), .A2(G106gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT6), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n390_), .A2(G99gat), .A3(G106gat), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT64), .ZN(new_n394_));
  AND2_X1   g193(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n395_));
  NOR2_X1   g194(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(G106gat), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n394_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NOR4_X1   g198(.A1(new_n395_), .A2(new_n396_), .A3(KEYINPUT64), .A4(G106gat), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n387_), .B(new_n393_), .C1(new_n399_), .C2(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n379_), .A2(new_n378_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT7), .ZN(new_n403_));
  INV_X1    g202(.A(G99gat), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(new_n404_), .A3(new_n398_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n402_), .B1(new_n392_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT8), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT8), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n410_), .B(new_n402_), .C1(new_n392_), .C2(new_n407_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(KEYINPUT66), .A2(new_n401_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT10), .B(G99gat), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT64), .B1(new_n413_), .B2(G106gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n397_), .A2(new_n394_), .A3(new_n398_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n392_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT66), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n417_), .A3(new_n387_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G29gat), .B(G36gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G43gat), .B(G50gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n412_), .A2(new_n418_), .A3(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G232gat), .A2(G233gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT34), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n401_), .A2(KEYINPUT66), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n409_), .A2(new_n411_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(new_n418_), .ZN(new_n427_));
  XOR2_X1   g226(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n428_));
  XNOR2_X1  g227(.A(new_n421_), .B(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  AND2_X1   g229(.A1(new_n430_), .A2(KEYINPUT73), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(KEYINPUT73), .ZN(new_n432_));
  OAI221_X1 g231(.A(new_n422_), .B1(KEYINPUT35), .B2(new_n424_), .C1(new_n431_), .C2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n424_), .A2(KEYINPUT35), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(G190gat), .B(G218gat), .Z(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT74), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G134gat), .B(G162gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  NOR2_X1   g238(.A1(new_n439_), .A2(KEYINPUT36), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n435_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n439_), .B(KEYINPUT36), .Z(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n435_), .A2(new_n443_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n377_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G15gat), .B(G22gat), .ZN(new_n447_));
  INV_X1    g246(.A(G1gat), .ZN(new_n448_));
  INV_X1    g247(.A(G8gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT14), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G1gat), .B(G8gat), .ZN(new_n452_));
  XOR2_X1   g251(.A(new_n451_), .B(new_n452_), .Z(new_n453_));
  NAND2_X1  g252(.A1(G231gat), .A2(G233gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n453_), .B(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT67), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G57gat), .B(G64gat), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n456_), .B1(new_n457_), .B2(KEYINPUT11), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(new_n457_), .A2(KEYINPUT11), .ZN(new_n460_));
  XOR2_X1   g259(.A(G71gat), .B(G78gat), .Z(new_n461_));
  NAND3_X1  g260(.A1(new_n457_), .A2(new_n456_), .A3(KEYINPUT11), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n459_), .A2(new_n460_), .A3(new_n461_), .A4(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n461_), .B1(KEYINPUT11), .B2(new_n457_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n462_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n464_), .B1(new_n465_), .B2(new_n458_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n455_), .B(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT17), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G127gat), .B(G155gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT16), .ZN(new_n472_));
  XOR2_X1   g271(.A(G183gat), .B(G211gat), .Z(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n469_), .A2(new_n470_), .A3(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(KEYINPUT17), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n475_), .B1(new_n469_), .B2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n453_), .B(new_n421_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G229gat), .A2(G233gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n453_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n429_), .A2(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n480_), .B1(new_n453_), .B2(new_n421_), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n478_), .A2(new_n480_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G113gat), .B(G141gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT78), .ZN(new_n486_));
  XOR2_X1   g285(.A(G169gat), .B(G197gat), .Z(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n484_), .A2(new_n488_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n427_), .A2(KEYINPUT12), .A3(new_n468_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n467_), .B1(new_n412_), .B2(new_n418_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n493_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n467_), .A2(new_n426_), .A3(new_n425_), .A4(new_n418_), .ZN(new_n498_));
  INV_X1    g297(.A(G230gat), .ZN(new_n499_));
  INV_X1    g298(.A(G233gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(KEYINPUT69), .B1(new_n497_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n498_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n501_), .B1(new_n505_), .B2(new_n494_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n503_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n427_), .A2(new_n468_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(new_n495_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT69), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n507_), .A2(new_n509_), .A3(new_n510_), .A4(new_n493_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n504_), .A2(new_n506_), .A3(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G120gat), .B(G148gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT5), .ZN(new_n514_));
  XOR2_X1   g313(.A(G176gat), .B(G204gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n512_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n512_), .A2(new_n516_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(KEYINPUT70), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT70), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n512_), .A2(new_n520_), .A3(new_n516_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n522_), .A2(KEYINPUT13), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n519_), .A2(KEYINPUT13), .A3(new_n521_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT71), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n523_), .A2(KEYINPUT71), .A3(new_n524_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n492_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n446_), .A2(new_n477_), .A3(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(G1gat), .B1(new_n530_), .B2(new_n368_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT38), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n527_), .A2(new_n528_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT76), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT37), .ZN(new_n535_));
  OAI211_X1 g334(.A(KEYINPUT75), .B(new_n535_), .C1(new_n441_), .C2(new_n444_), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n435_), .A2(new_n443_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n535_), .A2(KEYINPUT75), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n435_), .A2(new_n440_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n535_), .A2(KEYINPUT75), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .A4(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n536_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n477_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n534_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n536_), .A2(new_n541_), .A3(KEYINPUT76), .A4(new_n477_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n533_), .A2(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n547_), .A2(KEYINPUT77), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(KEYINPUT77), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n377_), .A2(new_n492_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n551_), .A2(new_n448_), .A3(new_n374_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n552_), .A2(KEYINPUT99), .A3(new_n532_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT99), .B1(new_n552_), .B2(new_n532_), .ZN(new_n554_));
  OAI221_X1 g353(.A(new_n531_), .B1(new_n532_), .B2(new_n552_), .C1(new_n553_), .C2(new_n554_), .ZN(G1324gat));
  NAND3_X1  g354(.A1(new_n551_), .A2(new_n449_), .A3(new_n372_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n372_), .ZN(new_n557_));
  OAI21_X1  g356(.A(G8gat), .B1(new_n530_), .B2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n558_), .A2(KEYINPUT39), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(KEYINPUT39), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n556_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT40), .Z(G1325gat));
  NAND4_X1  g361(.A1(new_n446_), .A2(new_n477_), .A3(new_n363_), .A4(new_n529_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(G15gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT100), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT100), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n563_), .A2(new_n566_), .A3(G15gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT41), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(G15gat), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n551_), .A2(new_n571_), .A3(new_n363_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n565_), .A2(KEYINPUT41), .A3(new_n567_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT101), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(G1326gat));
  OAI21_X1  g375(.A(G22gat), .B1(new_n530_), .B2(new_n340_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT42), .ZN(new_n578_));
  INV_X1    g377(.A(G22gat), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n551_), .A2(new_n579_), .A3(new_n370_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(G1327gat));
  AND2_X1   g380(.A1(new_n529_), .A2(new_n543_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n542_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n377_), .A2(KEYINPUT43), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT43), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n373_), .A2(new_n376_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n351_), .A2(new_n340_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n300_), .A2(new_n301_), .A3(new_n303_), .A4(new_n307_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n588_), .B1(new_n248_), .B2(KEYINPUT97), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n587_), .B1(new_n589_), .B2(new_n310_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n369_), .A2(new_n370_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n375_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n586_), .B1(new_n590_), .B2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n585_), .B1(new_n593_), .B2(new_n542_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n582_), .B1(new_n584_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT44), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(KEYINPUT43), .B1(new_n377_), .B2(new_n583_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n593_), .A2(new_n585_), .A3(new_n542_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(KEYINPUT44), .A3(new_n582_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT102), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n597_), .A2(new_n601_), .A3(new_n602_), .A4(new_n374_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n603_), .A2(G29gat), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n597_), .A2(new_n601_), .A3(new_n374_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT102), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT103), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  AND4_X1   g406(.A1(KEYINPUT103), .A2(new_n606_), .A3(G29gat), .A4(new_n603_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n445_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n609_), .A2(new_n477_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n550_), .A2(new_n533_), .A3(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n368_), .A2(G29gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT104), .ZN(new_n613_));
  OAI22_X1  g412(.A1(new_n607_), .A2(new_n608_), .B1(new_n611_), .B2(new_n613_), .ZN(G1328gat));
  NOR2_X1   g413(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT105), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT46), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n611_), .A2(G36gat), .A3(new_n557_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT45), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n597_), .A2(new_n601_), .A3(new_n372_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(G36gat), .ZN(new_n623_));
  AOI211_X1 g422(.A(new_n615_), .B(new_n618_), .C1(new_n621_), .C2(new_n623_), .ZN(new_n624_));
  AND4_X1   g423(.A1(new_n616_), .A2(new_n621_), .A3(new_n617_), .A4(new_n623_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1329gat));
  AND2_X1   g425(.A1(new_n597_), .A2(new_n601_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n627_), .A2(G43gat), .A3(new_n363_), .ZN(new_n628_));
  INV_X1    g427(.A(G43gat), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n629_), .B1(new_n611_), .B2(new_n375_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(G1330gat));
  INV_X1    g432(.A(new_n611_), .ZN(new_n634_));
  AOI21_X1  g433(.A(G50gat), .B1(new_n634_), .B2(new_n370_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n370_), .A2(G50gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n627_), .B2(new_n636_), .ZN(G1331gat));
  AND2_X1   g436(.A1(new_n527_), .A2(new_n528_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n638_), .A2(new_n477_), .A3(new_n492_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n446_), .ZN(new_n640_));
  INV_X1    g439(.A(G57gat), .ZN(new_n641_));
  NOR4_X1   g440(.A1(new_n639_), .A2(new_n640_), .A3(new_n641_), .A4(new_n368_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT110), .ZN(new_n643_));
  INV_X1    g442(.A(new_n492_), .ZN(new_n644_));
  OAI21_X1  g443(.A(KEYINPUT108), .B1(new_n377_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT108), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n593_), .A2(new_n646_), .A3(new_n492_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT109), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n546_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(KEYINPUT107), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT107), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n638_), .A2(new_n652_), .A3(new_n546_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n648_), .A2(new_n649_), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n649_), .B1(new_n648_), .B2(new_n654_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n643_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n377_), .A2(KEYINPUT108), .A3(new_n644_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n646_), .B1(new_n593_), .B2(new_n492_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n651_), .A2(new_n653_), .ZN(new_n661_));
  OAI21_X1  g460(.A(KEYINPUT109), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n648_), .A2(new_n649_), .A3(new_n654_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(KEYINPUT110), .A3(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n657_), .A2(new_n664_), .A3(new_n374_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n641_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT111), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n665_), .A2(KEYINPUT111), .A3(new_n641_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n642_), .B1(new_n668_), .B2(new_n669_), .ZN(G1332gat));
  INV_X1    g469(.A(G64gat), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n640_), .A2(new_n639_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(new_n372_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT48), .Z(new_n674_));
  NOR2_X1   g473(.A1(new_n655_), .A2(new_n656_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(new_n671_), .A3(new_n372_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1333gat));
  AOI21_X1  g476(.A(new_n354_), .B1(new_n672_), .B2(new_n363_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT49), .Z(new_n679_));
  NAND3_X1  g478(.A1(new_n675_), .A2(new_n354_), .A3(new_n363_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1334gat));
  INV_X1    g480(.A(G78gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n672_), .B2(new_n370_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT50), .Z(new_n684_));
  NAND3_X1  g483(.A1(new_n675_), .A2(new_n682_), .A3(new_n370_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1335gat));
  AND3_X1   g485(.A1(new_n648_), .A2(new_n638_), .A3(new_n610_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n687_), .A2(new_n384_), .A3(new_n374_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n543_), .A2(new_n492_), .ZN(new_n689_));
  OR3_X1    g488(.A1(new_n533_), .A2(KEYINPUT112), .A3(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT112), .B1(new_n533_), .B2(new_n689_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n600_), .A2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G85gat), .B1(new_n693_), .B2(new_n368_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n688_), .A2(new_n694_), .ZN(G1336gat));
  NAND3_X1  g494(.A1(new_n687_), .A2(new_n385_), .A3(new_n372_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G92gat), .B1(new_n693_), .B2(new_n557_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT113), .ZN(G1337gat));
  NAND3_X1  g498(.A1(new_n687_), .A2(new_n397_), .A3(new_n363_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G99gat), .B1(new_n693_), .B2(new_n375_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g502(.A1(new_n687_), .A2(new_n398_), .A3(new_n370_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT52), .ZN(new_n705_));
  INV_X1    g504(.A(new_n693_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(new_n370_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(new_n707_), .B2(G106gat), .ZN(new_n708_));
  AOI211_X1 g507(.A(KEYINPUT52), .B(new_n398_), .C1(new_n706_), .C2(new_n370_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n704_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT53), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT53), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n712_), .B(new_n704_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1339gat));
  INV_X1    g513(.A(KEYINPUT57), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n517_), .A2(new_n644_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT55), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n504_), .A2(new_n718_), .A3(new_n511_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT114), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n504_), .A2(KEYINPUT114), .A3(new_n718_), .A4(new_n511_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n509_), .A2(new_n498_), .A3(new_n493_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n501_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n507_), .A2(new_n509_), .A3(new_n493_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n718_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n723_), .A2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT115), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n723_), .A2(KEYINPUT115), .A3(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT56), .B1(new_n733_), .B2(new_n516_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT115), .B1(new_n723_), .B2(new_n728_), .ZN(new_n735_));
  AOI211_X1 g534(.A(new_n730_), .B(new_n727_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n736_));
  OAI211_X1 g535(.A(KEYINPUT56), .B(new_n516_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n717_), .B1(new_n734_), .B2(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n479_), .B1(new_n453_), .B2(new_n421_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n482_), .A2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n488_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n490_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n522_), .A2(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n445_), .B1(new_n739_), .B2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n715_), .B1(new_n745_), .B2(KEYINPUT116), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n516_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT56), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n716_), .B1(new_n749_), .B2(new_n737_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n744_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n609_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(new_n753_), .A3(KEYINPUT57), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n746_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n517_), .A2(new_n743_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n749_), .B2(new_n737_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n583_), .B1(new_n757_), .B2(KEYINPUT58), .ZN(new_n758_));
  INV_X1    g557(.A(new_n756_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n759_), .B1(new_n734_), .B2(new_n738_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT58), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n758_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n477_), .B1(new_n755_), .B2(new_n763_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n525_), .A2(new_n583_), .A3(new_n477_), .A4(new_n492_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT54), .Z(new_n766_));
  NOR2_X1   g565(.A1(new_n764_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n373_), .A2(new_n374_), .A3(new_n363_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n768_), .A2(KEYINPUT59), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  OR3_X1    g569(.A1(new_n767_), .A2(KEYINPUT118), .A3(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT118), .B1(new_n767_), .B2(new_n770_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  OAI211_X1 g572(.A(KEYINPUT58), .B(new_n759_), .C1(new_n734_), .C2(new_n738_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n542_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n749_), .A2(new_n737_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT58), .B1(new_n776_), .B2(new_n759_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n773_), .B1(new_n775_), .B2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n758_), .A2(new_n762_), .A3(KEYINPUT117), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n752_), .A2(new_n753_), .A3(KEYINPUT57), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT57), .B1(new_n752_), .B2(new_n753_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n778_), .B(new_n779_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n766_), .B1(new_n782_), .B2(new_n543_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT59), .B1(new_n783_), .B2(new_n768_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n771_), .A2(new_n772_), .A3(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(G113gat), .B1(new_n785_), .B2(new_n492_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n783_), .A2(new_n768_), .ZN(new_n787_));
  INV_X1    g586(.A(G113gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n787_), .A2(new_n788_), .A3(new_n644_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(G1340gat));
  OAI21_X1  g589(.A(G120gat), .B1(new_n785_), .B2(new_n533_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT60), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT119), .B1(new_n792_), .B2(G120gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(G120gat), .B1(new_n638_), .B2(new_n792_), .ZN(new_n794_));
  MUX2_X1   g593(.A(new_n793_), .B(KEYINPUT119), .S(new_n794_), .Z(new_n795_));
  NAND2_X1  g594(.A1(new_n787_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n791_), .A2(new_n796_), .ZN(G1341gat));
  OAI21_X1  g596(.A(G127gat), .B1(new_n785_), .B2(new_n543_), .ZN(new_n798_));
  INV_X1    g597(.A(G127gat), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n787_), .A2(new_n799_), .A3(new_n477_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n798_), .A2(new_n800_), .ZN(G1342gat));
  OAI21_X1  g600(.A(G134gat), .B1(new_n785_), .B2(new_n583_), .ZN(new_n802_));
  INV_X1    g601(.A(G134gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n787_), .A2(new_n803_), .A3(new_n445_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1343gat));
  INV_X1    g604(.A(new_n783_), .ZN(new_n806_));
  NOR4_X1   g605(.A1(new_n372_), .A2(new_n340_), .A3(new_n368_), .A4(new_n363_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n644_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n638_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g612(.A1(new_n808_), .A2(new_n543_), .ZN(new_n814_));
  XOR2_X1   g613(.A(KEYINPUT61), .B(G155gat), .Z(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(G1346gat));
  NAND4_X1  g615(.A1(new_n806_), .A2(G162gat), .A3(new_n542_), .A4(new_n807_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n775_), .A2(new_n773_), .A3(new_n777_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT117), .B1(new_n758_), .B2(new_n762_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n477_), .B1(new_n820_), .B2(new_n755_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n445_), .B(new_n807_), .C1(new_n821_), .C2(new_n766_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823_));
  INV_X1    g622(.A(G162gat), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n817_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT121), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  OAI211_X1 g628(.A(KEYINPUT121), .B(new_n817_), .C1(new_n825_), .C2(new_n826_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(G1347gat));
  XOR2_X1   g630(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n832_));
  OR2_X1    g631(.A1(new_n764_), .A2(new_n766_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n557_), .A2(new_n374_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n363_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND4_X1  g635(.A1(new_n833_), .A2(new_n644_), .A3(new_n340_), .A4(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n832_), .B1(new_n837_), .B2(KEYINPUT22), .ZN(new_n838_));
  OAI21_X1  g637(.A(G169gat), .B1(new_n837_), .B2(new_n832_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n269_), .B2(new_n838_), .ZN(G1348gat));
  NOR2_X1   g640(.A1(new_n533_), .A2(G176gat), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n833_), .A2(new_n340_), .A3(new_n836_), .A4(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n638_), .A2(new_n836_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT123), .B1(new_n783_), .B2(new_n370_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT123), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n846_), .B(new_n340_), .C1(new_n821_), .C2(new_n766_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n844_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n843_), .B1(new_n848_), .B2(new_n270_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT124), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n851_), .B(new_n843_), .C1(new_n848_), .C2(new_n270_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1349gat));
  NAND2_X1  g652(.A1(new_n845_), .A2(new_n847_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n835_), .A2(new_n543_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G183gat), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  AND4_X1   g655(.A1(new_n340_), .A2(new_n833_), .A3(new_n276_), .A4(new_n855_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1350gat));
  NAND3_X1  g657(.A1(new_n833_), .A2(new_n340_), .A3(new_n836_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G190gat), .B1(new_n859_), .B2(new_n583_), .ZN(new_n860_));
  OR2_X1    g659(.A1(new_n609_), .A2(new_n277_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n859_), .B2(new_n861_), .ZN(G1351gat));
  NOR4_X1   g661(.A1(new_n557_), .A2(new_n340_), .A3(new_n374_), .A4(new_n363_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n806_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n644_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g666(.A1(new_n864_), .A2(new_n533_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(KEYINPUT125), .B(G204gat), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1353gat));
  NOR2_X1   g669(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n871_));
  AND2_X1   g670(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n872_));
  NOR4_X1   g671(.A1(new_n864_), .A2(new_n543_), .A3(new_n871_), .A4(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n864_), .B2(new_n543_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT126), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI211_X1 g675(.A(KEYINPUT126), .B(new_n871_), .C1(new_n864_), .C2(new_n543_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n873_), .B1(new_n876_), .B2(new_n877_), .ZN(G1354gat));
  NOR3_X1   g677(.A1(new_n864_), .A2(KEYINPUT127), .A3(new_n609_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(G218gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(KEYINPUT127), .B1(new_n864_), .B2(new_n609_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n542_), .A2(G218gat), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n880_), .A2(new_n881_), .B1(new_n865_), .B2(new_n882_), .ZN(G1355gat));
endmodule


