//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n866_, new_n867_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_;
  AND3_X1   g000(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n202_));
  AOI21_X1  g001(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  INV_X1    g004(.A(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(KEYINPUT24), .A3(new_n208_), .ZN(new_n209_));
  OR3_X1    g008(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n210_));
  AND3_X1   g009(.A1(new_n204_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n213_));
  AND2_X1   g012(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n215_));
  OAI22_X1  g014(.A1(new_n212_), .A2(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT81), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT25), .B(G183gat), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT26), .B(G190gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(new_n220_), .A3(KEYINPUT81), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n211_), .A2(new_n218_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT82), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT22), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n206_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(G169gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OR2_X1    g028(.A1(G183gat), .A2(G190gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n229_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n205_), .B(new_n206_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n226_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n222_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT30), .B(G15gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G71gat), .B(G99gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G227gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G43gat), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G113gat), .B(G120gat), .ZN(new_n243_));
  INV_X1    g042(.A(G134gat), .ZN(new_n244_));
  OR2_X1    g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n244_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT83), .B(G127gat), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT84), .ZN(new_n250_));
  NOR3_X1   g049(.A1(new_n248_), .A2(new_n249_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n245_), .A2(new_n246_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n247_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT84), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n251_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT31), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT85), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n239_), .A2(new_n241_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n242_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n257_), .B(KEYINPUT31), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(KEYINPUT85), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(new_n242_), .B2(new_n263_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n264_), .A2(new_n268_), .ZN(new_n269_));
  NOR2_X1   g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G141gat), .A2(G148gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n273_), .A2(KEYINPUT1), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT86), .ZN(new_n275_));
  NOR2_X1   g074(.A1(G155gat), .A2(G162gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(KEYINPUT1), .B2(new_n273_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n271_), .B(new_n272_), .C1(new_n275_), .C2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n270_), .A2(KEYINPUT88), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT2), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(G141gat), .B2(G148gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n272_), .A2(KEYINPUT2), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n280_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(G141gat), .ZN(new_n285_));
  INV_X1    g084(.A(G148gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(new_n286_), .A3(KEYINPUT87), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT88), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT3), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT3), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n287_), .A2(new_n288_), .A3(new_n291_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n284_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT89), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n273_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n272_), .A2(KEYINPUT2), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n281_), .A2(G141gat), .A3(G148gat), .ZN(new_n297_));
  AOI22_X1  g096(.A1(new_n296_), .A2(new_n297_), .B1(KEYINPUT88), .B2(new_n270_), .ZN(new_n298_));
  AOI211_X1 g097(.A(KEYINPUT88), .B(KEYINPUT3), .C1(new_n270_), .C2(KEYINPUT87), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n291_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n300_));
  OAI211_X1 g099(.A(new_n294_), .B(new_n298_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n277_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n279_), .B1(new_n295_), .B2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n248_), .A2(new_n249_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n298_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT89), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n308_), .A2(new_n277_), .A3(new_n301_), .A4(new_n273_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT90), .ZN(new_n310_));
  AND3_X1   g109(.A1(new_n309_), .A2(new_n310_), .A3(new_n279_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(new_n309_), .B2(new_n279_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OAI211_X1 g112(.A(KEYINPUT4), .B(new_n306_), .C1(new_n313_), .C2(new_n257_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G225gat), .A2(G233gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(new_n315_), .B(KEYINPUT96), .Z(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n303_), .A2(KEYINPUT90), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n309_), .A2(new_n310_), .A3(new_n279_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n257_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT4), .ZN(new_n321_));
  AOI21_X1  g120(.A(KEYINPUT97), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n304_), .A2(KEYINPUT84), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n254_), .A2(new_n255_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n250_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n321_), .B(new_n326_), .C1(new_n311_), .C2(new_n312_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT97), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  OAI211_X1 g128(.A(new_n314_), .B(new_n317_), .C1(new_n322_), .C2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n318_), .A2(new_n319_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n305_), .B1(new_n331_), .B2(new_n326_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n315_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G1gat), .B(G29gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G85gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(KEYINPUT0), .B(G57gat), .ZN(new_n337_));
  XOR2_X1   g136(.A(new_n336_), .B(new_n337_), .Z(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n330_), .A2(new_n333_), .A3(new_n338_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n269_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT92), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT29), .B1(new_n311_), .B2(new_n312_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G228gat), .A2(G233gat), .ZN(new_n346_));
  INV_X1    g145(.A(G197gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n347_), .A2(G204gat), .ZN(new_n348_));
  INV_X1    g147(.A(G204gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n349_), .A2(G197gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT21), .B1(new_n348_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(G197gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n347_), .A2(G204gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT21), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n352_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  XNOR2_X1  g154(.A(G211gat), .B(G218gat), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n351_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n356_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n354_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n345_), .A2(new_n346_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n363_), .B1(new_n309_), .B2(new_n279_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n357_), .A2(new_n360_), .ZN(new_n365_));
  OAI211_X1 g164(.A(G228gat), .B(G233gat), .C1(new_n364_), .C2(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G78gat), .B(G106gat), .Z(new_n367_));
  NOR2_X1   g166(.A1(new_n367_), .A2(KEYINPUT91), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n362_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n362_), .B2(new_n366_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT28), .B1(new_n331_), .B2(KEYINPUT29), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT28), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n313_), .A2(new_n373_), .A3(new_n363_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G22gat), .B(G50gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n372_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n344_), .B1(new_n371_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n362_), .A2(new_n366_), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n382_), .A2(new_n367_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n367_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n380_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n368_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n382_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n362_), .A2(new_n366_), .A3(new_n368_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n372_), .A2(new_n374_), .A3(new_n376_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n376_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n389_), .A2(new_n392_), .A3(KEYINPUT92), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n381_), .A2(new_n385_), .A3(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G8gat), .B(G36gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(G92gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT18), .B(G64gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G226gat), .A2(G233gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AND2_X1   g201(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n206_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n232_), .A2(new_n405_), .A3(new_n208_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n204_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n216_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n406_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n409_), .A2(new_n361_), .A3(KEYINPUT94), .ZN(new_n410_));
  AOI21_X1  g209(.A(KEYINPUT94), .B1(new_n409_), .B2(new_n361_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n413_));
  INV_X1    g212(.A(new_n234_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n216_), .A2(new_n217_), .ZN(new_n415_));
  AOI21_X1  g214(.A(KEYINPUT81), .B1(new_n219_), .B2(new_n220_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n414_), .B1(new_n417_), .B2(new_n211_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n413_), .B1(new_n418_), .B2(new_n365_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n402_), .B1(new_n412_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT20), .B1(new_n409_), .B2(new_n361_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n235_), .A2(new_n361_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n422_), .A2(new_n423_), .A3(new_n402_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n398_), .B1(new_n420_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n409_), .A2(new_n361_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT94), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n365_), .A2(new_n222_), .A3(new_n234_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n409_), .A2(new_n361_), .A3(KEYINPUT94), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(KEYINPUT20), .A4(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n401_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n398_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n422_), .A2(new_n423_), .A3(new_n402_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n425_), .A2(KEYINPUT95), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT95), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n432_), .A2(new_n437_), .A3(new_n433_), .A4(new_n434_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT27), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n421_), .A2(KEYINPUT100), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT100), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n443_), .B(KEYINPUT20), .C1(new_n409_), .C2(new_n361_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n444_), .A3(new_n423_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT101), .B1(new_n446_), .B2(new_n402_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n412_), .A2(new_n419_), .A3(new_n402_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT101), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n445_), .A2(new_n449_), .A3(new_n401_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n447_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT102), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n451_), .A2(new_n452_), .A3(new_n398_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n452_), .B1(new_n451_), .B2(new_n398_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n435_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n453_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n441_), .B1(new_n456_), .B2(KEYINPUT27), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n343_), .A2(new_n394_), .A3(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT98), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(KEYINPUT33), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n341_), .A2(new_n460_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n320_), .A2(new_n305_), .A3(new_n316_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n315_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n463_), .B1(new_n332_), .B2(KEYINPUT4), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n327_), .A2(new_n328_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n331_), .A2(KEYINPUT97), .A3(new_n321_), .A4(new_n326_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n462_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n439_), .B1(new_n468_), .B2(new_n339_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n460_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n330_), .A2(new_n333_), .A3(new_n338_), .A4(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n461_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n433_), .A2(KEYINPUT32), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n473_), .A2(KEYINPUT99), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n432_), .A2(new_n434_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n473_), .A2(KEYINPUT99), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n474_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n473_), .B2(new_n451_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n330_), .A2(new_n333_), .A3(new_n338_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n338_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n478_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n472_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n394_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n381_), .A2(new_n385_), .A3(new_n393_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n479_), .A2(new_n480_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n457_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n483_), .A2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n458_), .B1(new_n487_), .B2(new_n269_), .ZN(new_n488_));
  XOR2_X1   g287(.A(KEYINPUT10), .B(G99gat), .Z(new_n489_));
  INV_X1    g288(.A(G106gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT64), .ZN(new_n492_));
  XOR2_X1   g291(.A(G85gat), .B(G92gat), .Z(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT9), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G99gat), .A2(G106gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT6), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT9), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(G85gat), .A3(G92gat), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n492_), .A2(new_n494_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT65), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT65), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n492_), .A2(new_n502_), .A3(new_n494_), .A4(new_n499_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT66), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n496_), .B1(new_n504_), .B2(KEYINPUT7), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(KEYINPUT7), .ZN(new_n506_));
  NOR2_X1   g305(.A1(G99gat), .A2(G106gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n493_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT8), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT8), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n511_), .B(new_n493_), .C1(new_n505_), .C2(new_n508_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n501_), .A2(new_n503_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT67), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND4_X1  g315(.A1(new_n501_), .A2(KEYINPUT67), .A3(new_n503_), .A4(new_n513_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT69), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT70), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n521_), .A2(new_n522_), .A3(KEYINPUT11), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n522_), .B1(new_n521_), .B2(KEYINPUT11), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n521_), .A2(KEYINPUT11), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT68), .B(G71gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(G78gat), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  OAI22_X1  g329(.A1(new_n523_), .A2(new_n524_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n518_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n516_), .A2(new_n517_), .A3(new_n532_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G230gat), .A2(G233gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT12), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n535_), .A2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n532_), .A2(new_n514_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT12), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n541_), .A2(new_n534_), .A3(new_n537_), .A4(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n539_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT5), .B(G176gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(G204gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G120gat), .B(G148gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(new_n548_), .Z(new_n549_));
  XOR2_X1   g348(.A(new_n549_), .B(KEYINPUT71), .Z(new_n550_));
  NAND2_X1  g349(.A1(new_n545_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT72), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n545_), .A2(new_n549_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n545_), .A2(KEYINPUT72), .A3(new_n550_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n553_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(KEYINPUT13), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT13), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n553_), .A2(new_n554_), .A3(new_n558_), .A4(new_n555_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G43gat), .B(G50gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(G29gat), .B(G36gat), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT15), .Z(new_n567_));
  XNOR2_X1  g366(.A(G15gat), .B(G22gat), .ZN(new_n568_));
  INV_X1    g367(.A(G1gat), .ZN(new_n569_));
  INV_X1    g368(.A(G8gat), .ZN(new_n570_));
  OAI21_X1  g369(.A(KEYINPUT14), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G1gat), .B(G8gat), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n573_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n567_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n566_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(new_n575_), .A3(new_n574_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G229gat), .A2(G233gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT80), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n576_), .A2(new_n566_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n579_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(G229gat), .A3(G233gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G169gat), .B(G197gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n588_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n591_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n488_), .A2(new_n561_), .A3(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n597_));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G183gat), .B(G211gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT17), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n576_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n532_), .B(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT17), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n603_), .B1(new_n607_), .B2(new_n601_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n606_), .A2(KEYINPUT79), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n518_), .A2(new_n578_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n514_), .A2(new_n567_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT35), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT73), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n615_), .B1(new_n613_), .B2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT34), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n614_), .A2(new_n620_), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n619_), .A2(KEYINPUT35), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n612_), .A2(new_n619_), .A3(new_n613_), .A4(new_n617_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(G190gat), .B(G218gat), .Z(new_n625_));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n628_));
  NAND3_X1  g427(.A1(new_n624_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT37), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n627_), .B(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .A4(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n629_), .A2(new_n630_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT77), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n632_), .B(KEYINPUT76), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .A4(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n629_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT37), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n635_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(KEYINPUT77), .A3(KEYINPUT37), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n611_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n596_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n644_), .A2(new_n569_), .A3(new_n342_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT38), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n647_), .B1(new_n560_), .B2(new_n594_), .ZN(new_n648_));
  AOI211_X1 g447(.A(KEYINPUT103), .B(new_n595_), .C1(new_n557_), .C2(new_n559_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n457_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n484_), .B1(new_n481_), .B2(new_n472_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n269_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n458_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n629_), .A2(new_n633_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(new_n611_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n650_), .A2(new_n655_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AOI211_X1 g459(.A(KEYINPUT104), .B(new_n569_), .C1(new_n660_), .C2(new_n342_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT104), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n342_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n663_), .B2(G1gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n646_), .B1(new_n661_), .B2(new_n664_), .ZN(G1324gat));
  INV_X1    g464(.A(new_n457_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n644_), .A2(new_n570_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT39), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n660_), .A2(new_n666_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n669_), .B2(G8gat), .ZN(new_n670_));
  AOI211_X1 g469(.A(KEYINPUT39), .B(new_n570_), .C1(new_n660_), .C2(new_n666_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n667_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT40), .Z(G1325gat));
  OR3_X1    g472(.A1(new_n643_), .A2(G15gat), .A3(new_n269_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n269_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n660_), .A2(new_n675_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n676_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(KEYINPUT41), .B1(new_n676_), .B2(G15gat), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n677_), .B2(new_n678_), .ZN(G1326gat));
  OR3_X1    g478(.A1(new_n643_), .A2(G22gat), .A3(new_n394_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G22gat), .B1(new_n659_), .B2(new_n394_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n681_), .A2(KEYINPUT42), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(KEYINPUT42), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(G1327gat));
  NOR2_X1   g483(.A1(new_n656_), .A2(new_n610_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n596_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G29gat), .B1(new_n687_), .B2(new_n342_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n640_), .A2(new_n641_), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n689_), .B(new_n690_), .C1(new_n488_), .C2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n641_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n639_), .B2(new_n635_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n689_), .A2(new_n690_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n655_), .A2(new_n694_), .A3(new_n695_), .A4(new_n696_), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n692_), .A2(new_n697_), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n698_), .A2(KEYINPUT44), .A3(new_n650_), .A4(new_n611_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n692_), .A2(new_n650_), .A3(new_n697_), .A4(new_n611_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT44), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n699_), .A2(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(new_n342_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n688_), .B1(new_n704_), .B2(G29gat), .ZN(G1328gat));
  NOR3_X1   g504(.A1(new_n686_), .A2(G36gat), .A3(new_n457_), .ZN(new_n706_));
  XOR2_X1   g505(.A(new_n706_), .B(KEYINPUT45), .Z(new_n707_));
  NAND3_X1  g506(.A1(new_n699_), .A2(new_n666_), .A3(new_n702_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(G36gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G36gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(KEYINPUT46), .B(new_n707_), .C1(new_n710_), .C2(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1329gat));
  AOI21_X1  g515(.A(G43gat), .B1(new_n687_), .B2(new_n675_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n675_), .A2(G43gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n703_), .B2(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g519(.A(G50gat), .B1(new_n687_), .B2(new_n484_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n484_), .A2(G50gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n703_), .B2(new_n722_), .ZN(G1331gat));
  NOR2_X1   g522(.A1(new_n560_), .A2(new_n594_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n655_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(new_n658_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G57gat), .B1(new_n727_), .B2(new_n485_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n691_), .A2(new_n610_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n725_), .A2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n342_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n728_), .B1(G57gat), .B2(new_n731_), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT107), .Z(G1332gat));
  OAI21_X1  g532(.A(G64gat), .B1(new_n727_), .B2(new_n457_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT48), .ZN(new_n735_));
  INV_X1    g534(.A(new_n730_), .ZN(new_n736_));
  OR2_X1    g535(.A1(new_n457_), .A2(G64gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n735_), .B1(new_n736_), .B2(new_n737_), .ZN(G1333gat));
  NAND3_X1  g537(.A1(new_n726_), .A2(new_n675_), .A3(new_n658_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(new_n740_), .A3(G71gat), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT49), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n740_), .B1(new_n739_), .B2(G71gat), .ZN(new_n744_));
  OR3_X1    g543(.A1(new_n742_), .A2(new_n743_), .A3(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n743_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n730_), .A2(new_n675_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n745_), .B(new_n746_), .C1(G71gat), .C2(new_n747_), .ZN(G1334gat));
  OAI21_X1  g547(.A(G78gat), .B1(new_n727_), .B2(new_n394_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT50), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n394_), .A2(G78gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n736_), .B2(new_n751_), .ZN(G1335gat));
  INV_X1    g551(.A(G85gat), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n726_), .A2(new_n685_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(new_n485_), .ZN(new_n755_));
  OR2_X1    g554(.A1(new_n755_), .A2(KEYINPUT109), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(KEYINPUT109), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n698_), .A2(new_n611_), .A3(new_n724_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n342_), .A2(G85gat), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n756_), .B(new_n757_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT110), .Z(G1336gat));
  INV_X1    g560(.A(G92gat), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n758_), .A2(new_n762_), .A3(new_n457_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n754_), .ZN(new_n764_));
  AOI21_X1  g563(.A(G92gat), .B1(new_n764_), .B2(new_n666_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n758_), .B2(new_n269_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n489_), .A3(new_n675_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g569(.A(G106gat), .B1(new_n758_), .B2(new_n394_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT52), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n773_), .B(G106gat), .C1(new_n758_), .C2(new_n394_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n764_), .A2(new_n490_), .A3(new_n484_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n775_), .A2(new_n776_), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(G1339gat));
  XOR2_X1   g579(.A(KEYINPUT112), .B(KEYINPUT55), .Z(new_n781_));
  NAND2_X1  g580(.A1(new_n544_), .A2(new_n781_), .ZN(new_n782_));
  AOI22_X1  g581(.A1(new_n518_), .A2(new_n533_), .B1(new_n542_), .B2(KEYINPUT12), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT112), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n783_), .A2(new_n537_), .A3(new_n541_), .A4(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n541_), .A2(new_n534_), .A3(new_n543_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n538_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n782_), .A2(new_n786_), .A3(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n550_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT56), .B1(new_n789_), .B2(new_n550_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n790_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n789_), .A2(KEYINPUT113), .A3(KEYINPUT56), .A4(new_n550_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(new_n594_), .A3(new_n554_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n586_), .A2(new_n581_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n580_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n797_), .B(new_n591_), .C1(new_n798_), .C2(new_n581_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n592_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n556_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n657_), .B1(new_n796_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT57), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n595_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n805_), .A2(new_n554_), .B1(new_n556_), .B2(new_n800_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n804_), .B1(new_n806_), .B2(new_n657_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n789_), .A2(new_n550_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(KEYINPUT114), .A3(new_n790_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT114), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n789_), .A2(new_n812_), .A3(KEYINPUT56), .A4(new_n550_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n813_), .A2(new_n554_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(new_n814_), .A3(new_n800_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(KEYINPUT115), .A2(KEYINPUT58), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n816_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n811_), .A2(new_n814_), .A3(new_n800_), .A4(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n694_), .A3(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n803_), .A2(new_n807_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(new_n611_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n594_), .B1(new_n557_), .B2(new_n559_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n642_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n823_), .B1(new_n642_), .B2(new_n824_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n822_), .A2(new_n828_), .ZN(new_n829_));
  NOR4_X1   g628(.A1(new_n666_), .A2(new_n484_), .A3(new_n485_), .A4(new_n269_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(G113gat), .B1(new_n832_), .B2(new_n594_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n820_), .C1(new_n802_), .C2(KEYINPUT57), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n803_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n834_), .B1(new_n807_), .B2(new_n820_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n611_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n828_), .ZN(new_n839_));
  XOR2_X1   g638(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n830_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n831_), .A2(KEYINPUT59), .ZN(new_n842_));
  AND2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n594_), .A2(G113gat), .ZN(new_n844_));
  XOR2_X1   g643(.A(new_n844_), .B(KEYINPUT118), .Z(new_n845_));
  AOI21_X1  g644(.A(new_n833_), .B1(new_n843_), .B2(new_n845_), .ZN(G1340gat));
  NAND3_X1  g645(.A1(new_n841_), .A2(new_n561_), .A3(new_n842_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(G120gat), .ZN(new_n848_));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n560_), .B2(KEYINPUT60), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n832_), .B(new_n850_), .C1(KEYINPUT60), .C2(new_n849_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(G1341gat));
  AOI21_X1  g651(.A(G127gat), .B1(new_n832_), .B2(new_n610_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n610_), .A2(G127gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT119), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n843_), .B2(new_n855_), .ZN(G1342gat));
  XNOR2_X1  g655(.A(KEYINPUT120), .B(G134gat), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n841_), .A2(new_n842_), .A3(new_n694_), .A4(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n244_), .B1(new_n831_), .B2(new_n656_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1343gat));
  NOR3_X1   g659(.A1(new_n666_), .A2(new_n485_), .A3(new_n675_), .ZN(new_n861_));
  AND3_X1   g660(.A1(new_n829_), .A2(new_n484_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n594_), .ZN(new_n863_));
  XOR2_X1   g662(.A(KEYINPUT121), .B(G141gat), .Z(new_n864_));
  XNOR2_X1  g663(.A(new_n863_), .B(new_n864_), .ZN(G1344gat));
  NAND2_X1  g664(.A1(new_n862_), .A2(new_n561_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT122), .B(G148gat), .Z(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1345gat));
  NAND4_X1  g667(.A1(new_n829_), .A2(new_n484_), .A3(new_n610_), .A4(new_n861_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT123), .ZN(new_n870_));
  XOR2_X1   g669(.A(KEYINPUT61), .B(G155gat), .Z(new_n871_));
  AOI21_X1  g670(.A(new_n827_), .B1(new_n821_), .B2(new_n611_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n872_), .A2(new_n394_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n610_), .A4(new_n861_), .ZN(new_n875_));
  AND3_X1   g674(.A1(new_n870_), .A2(new_n871_), .A3(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n871_), .B1(new_n870_), .B2(new_n875_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1346gat));
  AOI21_X1  g677(.A(G162gat), .B1(new_n862_), .B2(new_n657_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n694_), .A2(G162gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT124), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n862_), .B2(new_n881_), .ZN(G1347gat));
  NAND2_X1  g681(.A1(new_n666_), .A2(new_n343_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n484_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n838_), .B2(new_n828_), .ZN(new_n886_));
  AOI211_X1 g685(.A(KEYINPUT62), .B(new_n205_), .C1(new_n886_), .C2(new_n594_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n839_), .A2(new_n594_), .A3(new_n884_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(G169gat), .ZN(new_n890_));
  INV_X1    g689(.A(new_n886_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n594_), .B1(new_n404_), .B2(new_n403_), .ZN(new_n892_));
  XOR2_X1   g691(.A(new_n892_), .B(KEYINPUT125), .Z(new_n893_));
  OAI22_X1  g692(.A1(new_n887_), .A2(new_n890_), .B1(new_n891_), .B2(new_n893_), .ZN(G1348gat));
  AOI21_X1  g693(.A(G176gat), .B1(new_n886_), .B2(new_n561_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n883_), .ZN(new_n896_));
  NOR4_X1   g695(.A1(new_n872_), .A2(new_n206_), .A3(new_n560_), .A4(new_n484_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(G1349gat));
  NOR3_X1   g697(.A1(new_n891_), .A2(new_n219_), .A3(new_n611_), .ZN(new_n899_));
  INV_X1    g698(.A(G183gat), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n829_), .A2(new_n394_), .A3(new_n610_), .A4(new_n896_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n900_), .B2(new_n901_), .ZN(G1350gat));
  OAI21_X1  g701(.A(G190gat), .B1(new_n891_), .B2(new_n691_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n886_), .A2(new_n220_), .A3(new_n657_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1351gat));
  NOR2_X1   g704(.A1(new_n394_), .A2(new_n342_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n666_), .A2(new_n269_), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n872_), .A2(new_n907_), .A3(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n594_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n561_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n912_), .B(new_n913_), .Z(G1353gat));
  AND2_X1   g713(.A1(new_n909_), .A2(new_n610_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n916_));
  AND2_X1   g715(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n916_), .B2(new_n917_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(new_n915_), .B2(new_n916_), .ZN(G1354gat));
  NOR2_X1   g718(.A1(new_n872_), .A2(new_n908_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n920_), .A2(G218gat), .A3(new_n906_), .A4(new_n694_), .ZN(new_n921_));
  NOR4_X1   g720(.A1(new_n872_), .A2(new_n907_), .A3(new_n656_), .A4(new_n908_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(G218gat), .B2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(KEYINPUT127), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT127), .ZN(new_n925_));
  OAI211_X1 g724(.A(new_n921_), .B(new_n925_), .C1(G218gat), .C2(new_n922_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1355gat));
endmodule


