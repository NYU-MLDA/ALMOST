//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n844_, new_n845_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_;
  XNOR2_X1  g000(.A(G22gat), .B(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT28), .ZN(new_n204_));
  NOR3_X1   g003(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT90), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT91), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G141gat), .ZN(new_n210_));
  INV_X1    g009(.A(G148gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n211_), .ZN(new_n213_));
  AOI22_X1  g012(.A1(new_n212_), .A2(KEYINPUT2), .B1(new_n213_), .B2(KEYINPUT3), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n206_), .A2(new_n209_), .A3(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n215_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(G155gat), .B2(G162gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(G155gat), .A3(G162gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT89), .ZN(new_n222_));
  AOI22_X1  g021(.A1(new_n217_), .A2(new_n220_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n223_), .B1(new_n222_), .B2(new_n221_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT88), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n212_), .B1(new_n213_), .B2(new_n225_), .ZN(new_n226_));
  OAI211_X1 g025(.A(new_n224_), .B(new_n226_), .C1(new_n225_), .C2(new_n213_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n218_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT29), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n204_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n218_), .A2(new_n227_), .ZN(new_n231_));
  NOR3_X1   g030(.A1(new_n231_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n203_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n228_), .A2(new_n204_), .A3(new_n229_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT28), .B1(new_n231_), .B2(KEYINPUT29), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(new_n202_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n233_), .A2(new_n236_), .A3(KEYINPUT96), .ZN(new_n237_));
  XOR2_X1   g036(.A(new_n237_), .B(KEYINPUT97), .Z(new_n238_));
  INV_X1    g037(.A(G106gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT95), .ZN(new_n240_));
  INV_X1    g039(.A(G204gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT92), .B1(new_n241_), .B2(G197gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT92), .ZN(new_n243_));
  INV_X1    g042(.A(G197gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(G204gat), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n242_), .B(new_n245_), .C1(new_n244_), .C2(G204gat), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT93), .ZN(new_n247_));
  OR3_X1    g046(.A1(new_n246_), .A2(new_n247_), .A3(KEYINPUT21), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n247_), .B1(new_n246_), .B2(KEYINPUT21), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n241_), .A2(G197gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n244_), .A2(G204gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(KEYINPUT21), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G211gat), .B(G218gat), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n248_), .A2(new_n249_), .A3(new_n252_), .A4(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n253_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n255_), .A2(KEYINPUT94), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(KEYINPUT94), .ZN(new_n257_));
  NAND4_X1  g056(.A1(new_n256_), .A2(KEYINPUT21), .A3(new_n246_), .A4(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n240_), .B1(new_n254_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G228gat), .A2(G233gat), .ZN(new_n260_));
  OAI21_X1  g059(.A(G78gat), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NOR3_X1   g061(.A1(new_n259_), .A2(G78gat), .A3(new_n260_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n239_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n263_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(new_n261_), .A3(G106gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n254_), .A2(new_n258_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n268_), .B1(KEYINPUT29), .B2(new_n231_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n264_), .A2(new_n266_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n233_), .A2(new_n236_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT96), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  AND2_X1   g072(.A1(new_n270_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n269_), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n262_), .A2(new_n263_), .A3(new_n239_), .ZN(new_n276_));
  AOI21_X1  g075(.A(G106gat), .B1(new_n265_), .B2(new_n261_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n275_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n238_), .A2(new_n274_), .A3(new_n278_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n273_), .A3(new_n270_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n237_), .B(KEYINPUT97), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G226gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT19), .ZN(new_n284_));
  INV_X1    g083(.A(G183gat), .ZN(new_n285_));
  INV_X1    g084(.A(G190gat), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT23), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT82), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT23), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(G183gat), .A3(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT79), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT25), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(G183gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT26), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G190gat), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n292_), .A2(new_n294_), .B1(new_n296_), .B2(KEYINPUT80), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT25), .B(G183gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(G190gat), .ZN(new_n299_));
  OAI221_X1 g098(.A(new_n297_), .B1(new_n292_), .B2(new_n298_), .C1(KEYINPUT80), .C2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G169gat), .ZN(new_n301_));
  INV_X1    g100(.A(G176gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(KEYINPUT24), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n306_), .A2(KEYINPUT81), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n303_), .A2(KEYINPUT24), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n308_), .B1(new_n306_), .B2(KEYINPUT81), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n291_), .A2(new_n300_), .A3(new_n307_), .A4(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n304_), .ZN(new_n311_));
  XOR2_X1   g110(.A(KEYINPUT22), .B(G169gat), .Z(new_n312_));
  INV_X1    g111(.A(KEYINPUT83), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n301_), .A2(KEYINPUT22), .ZN(new_n315_));
  AOI21_X1  g114(.A(G176gat), .B1(new_n315_), .B2(KEYINPUT83), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n311_), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n287_), .A2(new_n290_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n285_), .A2(new_n286_), .ZN(new_n319_));
  AND3_X1   g118(.A1(new_n318_), .A2(KEYINPUT84), .A3(new_n319_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT84), .B1(new_n318_), .B2(new_n319_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n317_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n310_), .A2(new_n322_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT20), .B1(new_n323_), .B2(new_n267_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n299_), .A2(new_n298_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n305_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT98), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n308_), .B1(new_n287_), .B2(new_n290_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n291_), .A2(new_n319_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n312_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n311_), .B1(new_n331_), .B2(new_n302_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  AOI22_X1  g132(.A1(new_n329_), .A2(new_n333_), .B1(new_n254_), .B2(new_n258_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n284_), .B1(new_n324_), .B2(new_n334_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n327_), .A2(new_n328_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n268_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n284_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n323_), .A2(new_n267_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n337_), .A2(KEYINPUT20), .A3(new_n338_), .A4(new_n339_), .ZN(new_n340_));
  XOR2_X1   g139(.A(G8gat), .B(G36gat), .Z(new_n341_));
  XNOR2_X1  g140(.A(G64gat), .B(G92gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(KEYINPUT99), .B(KEYINPUT18), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n335_), .A2(new_n340_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT20), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n347_), .B1(new_n268_), .B2(new_n336_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n338_), .B1(new_n348_), .B2(new_n339_), .ZN(new_n349_));
  NOR3_X1   g148(.A1(new_n324_), .A2(new_n334_), .A3(new_n284_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OAI211_X1 g150(.A(KEYINPUT27), .B(new_n346_), .C1(new_n351_), .C2(new_n345_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT27), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n335_), .A2(new_n340_), .A3(new_n345_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n345_), .B1(new_n335_), .B2(new_n340_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n352_), .A2(new_n356_), .A3(KEYINPUT104), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT104), .B1(new_n352_), .B2(new_n356_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n279_), .B(new_n282_), .C1(new_n357_), .C2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G227gat), .A2(G233gat), .ZN(new_n360_));
  XOR2_X1   g159(.A(new_n360_), .B(KEYINPUT85), .Z(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT30), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n323_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G15gat), .B(G43gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G127gat), .B(G134gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G113gat), .B(G120gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n368_), .A2(KEYINPUT87), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n366_), .B(new_n367_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n369_), .B1(new_n370_), .B2(KEYINPUT87), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT31), .ZN(new_n372_));
  XOR2_X1   g171(.A(G71gat), .B(G99gat), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT86), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n372_), .B(new_n374_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n365_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n365_), .A2(new_n375_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  XOR2_X1   g178(.A(G1gat), .B(G29gat), .Z(new_n380_));
  XNOR2_X1  g179(.A(G57gat), .B(G85gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n382_), .B(new_n383_), .Z(new_n384_));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n231_), .A2(new_n371_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n218_), .A2(new_n227_), .A3(new_n370_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n385_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT4), .B1(new_n231_), .B2(new_n371_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G225gat), .A2(G233gat), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT100), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n392_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n384_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n384_), .ZN(new_n397_));
  AOI211_X1 g196(.A(new_n397_), .B(new_n394_), .C1(new_n390_), .C2(new_n392_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n379_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT105), .B1(new_n359_), .B2(new_n401_), .ZN(new_n402_));
  OR2_X1    g201(.A1(new_n357_), .A2(new_n358_), .ZN(new_n403_));
  AND2_X1   g202(.A1(new_n280_), .A2(new_n281_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n280_), .A2(new_n281_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT105), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n378_), .A2(new_n399_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n403_), .A2(new_n406_), .A3(new_n407_), .A4(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n352_), .A2(new_n356_), .ZN(new_n410_));
  NOR2_X1   g209(.A1(new_n410_), .A2(new_n399_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n411_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n386_), .A2(KEYINPUT102), .A3(new_n387_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n392_), .ZN(new_n414_));
  AOI21_X1  g213(.A(KEYINPUT102), .B1(new_n386_), .B2(new_n387_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n384_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n392_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT103), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n419_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n416_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NOR3_X1   g221(.A1(new_n422_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n396_), .B(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n335_), .A2(new_n340_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n345_), .A2(KEYINPUT32), .ZN(new_n427_));
  MUX2_X1   g226(.A(new_n351_), .B(new_n426_), .S(new_n427_), .Z(new_n428_));
  AOI22_X1  g227(.A1(new_n423_), .A2(new_n425_), .B1(new_n399_), .B2(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n279_), .A2(new_n282_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n412_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n402_), .A2(new_n409_), .B1(new_n431_), .B2(new_n378_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT67), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G99gat), .A2(G106gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT6), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT6), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(G99gat), .A3(G106gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  AND2_X1   g237(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n439_));
  NOR2_X1   g238(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT64), .B1(new_n441_), .B2(new_n239_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT64), .ZN(new_n443_));
  NOR4_X1   g242(.A1(new_n439_), .A2(new_n440_), .A3(new_n443_), .A4(G106gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n438_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(G85gat), .A2(G92gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT9), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G85gat), .A2(G92gat), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(G85gat), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n451_), .A2(KEYINPUT65), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(KEYINPUT65), .ZN(new_n453_));
  NOR2_X1   g252(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n454_));
  AND2_X1   g253(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n455_));
  OAI22_X1  g254(.A1(new_n452_), .A2(new_n453_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n450_), .B1(new_n456_), .B2(new_n448_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n433_), .B1(new_n445_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n448_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n450_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n438_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT10), .B(G99gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n443_), .B1(new_n463_), .B2(G106gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n441_), .A2(KEYINPUT64), .A3(new_n239_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n462_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n461_), .A2(new_n466_), .A3(KEYINPUT67), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT8), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT68), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n438_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT7), .ZN(new_n471_));
  INV_X1    g270(.A(G99gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n239_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n435_), .A2(new_n437_), .A3(KEYINPUT68), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n470_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n449_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n479_), .A2(new_n446_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n468_), .B1(new_n478_), .B2(new_n480_), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n468_), .B(new_n480_), .C1(new_n462_), .C2(new_n475_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n458_), .B(new_n467_), .C1(new_n481_), .C2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G29gat), .B(G36gat), .Z(new_n485_));
  XOR2_X1   g284(.A(G43gat), .B(G50gat), .Z(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT15), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n485_), .B(new_n486_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT15), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n484_), .A2(new_n488_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G232gat), .A2(G233gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT34), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n494_), .A2(KEYINPUT35), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n492_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(KEYINPUT35), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n484_), .A2(new_n487_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n500_));
  OAI211_X1 g299(.A(KEYINPUT35), .B(new_n494_), .C1(new_n492_), .C2(new_n498_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G190gat), .B(G218gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G134gat), .B(G162gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(new_n505_), .B(KEYINPUT36), .Z(new_n506_));
  NAND2_X1  g305(.A1(new_n502_), .A2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n505_), .A2(KEYINPUT36), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n500_), .A2(new_n508_), .A3(new_n501_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n432_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G15gat), .B(G22gat), .ZN(new_n513_));
  INV_X1    g312(.A(G1gat), .ZN(new_n514_));
  INV_X1    g313(.A(G8gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT14), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n513_), .A2(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G1gat), .B(G8gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G231gat), .A2(G233gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G57gat), .B(G64gat), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n522_), .A2(KEYINPUT69), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT11), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(KEYINPUT69), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n523_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n522_), .A2(KEYINPUT69), .ZN(new_n527_));
  INV_X1    g326(.A(G64gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(G57gat), .ZN(new_n529_));
  INV_X1    g328(.A(G57gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(G64gat), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n529_), .A2(new_n531_), .A3(KEYINPUT69), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT11), .B1(new_n527_), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G71gat), .B(G78gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n526_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  OAI211_X1 g335(.A(KEYINPUT11), .B(new_n534_), .C1(new_n527_), .C2(new_n532_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n521_), .B(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G127gat), .B(G155gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT16), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G183gat), .B(G211gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT75), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n544_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n540_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n547_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n544_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n549_), .B1(KEYINPUT17), .B2(new_n550_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n548_), .B1(new_n551_), .B2(new_n540_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT106), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n484_), .A2(new_n539_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n480_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n475_), .B1(new_n438_), .B2(new_n469_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(new_n477_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n482_), .B1(new_n558_), .B2(new_n468_), .ZN(new_n559_));
  NAND4_X1  g358(.A1(new_n538_), .A2(new_n559_), .A3(new_n458_), .A4(new_n467_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G230gat), .A2(G233gat), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G120gat), .B(G148gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT5), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G176gat), .B(G204gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT70), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n560_), .A2(new_n569_), .A3(new_n562_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT12), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n484_), .A2(new_n571_), .A3(new_n539_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n571_), .B1(new_n484_), .B2(new_n539_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n570_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n569_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n564_), .B(new_n568_), .C1(new_n574_), .C2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT72), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n555_), .A2(KEYINPUT12), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n484_), .A2(new_n539_), .A3(new_n571_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n575_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n581_), .A2(new_n582_), .A3(new_n570_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n583_), .A2(KEYINPUT72), .A3(new_n564_), .A4(new_n568_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n578_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n564_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n568_), .B(KEYINPUT71), .Z(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n585_), .A2(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n592_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n488_), .A2(new_n519_), .A3(new_n491_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G229gat), .A2(G233gat), .ZN(new_n597_));
  INV_X1    g396(.A(new_n519_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(new_n489_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n596_), .A2(new_n597_), .A3(new_n599_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n600_), .A2(KEYINPUT77), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n487_), .A2(new_n519_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n597_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n600_), .A2(new_n605_), .A3(KEYINPUT77), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n601_), .A2(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(G113gat), .B(G141gat), .Z(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT78), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G169gat), .B(G197gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n609_), .B(new_n610_), .Z(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n607_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n611_), .B1(new_n601_), .B2(new_n606_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n554_), .B1(new_n595_), .B2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n615_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n594_), .A2(KEYINPUT106), .A3(new_n617_), .ZN(new_n618_));
  NAND4_X1  g417(.A1(new_n512_), .A2(new_n553_), .A3(new_n616_), .A4(new_n618_), .ZN(new_n619_));
  OR2_X1    g418(.A1(new_n619_), .A2(new_n400_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT74), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n507_), .A2(new_n621_), .A3(new_n509_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT37), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n507_), .A2(new_n621_), .A3(KEYINPUT37), .A4(new_n509_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n553_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT76), .ZN(new_n629_));
  NOR4_X1   g428(.A1(new_n629_), .A2(new_n432_), .A3(new_n615_), .A4(new_n595_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(new_n514_), .A3(new_n399_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632_));
  AOI22_X1  g431(.A1(G1gat), .A2(new_n620_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n633_), .B1(new_n632_), .B2(new_n631_), .ZN(G1324gat));
  INV_X1    g433(.A(new_n403_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n630_), .A2(new_n515_), .A3(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G8gat), .B1(new_n619_), .B2(new_n403_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n637_), .A2(KEYINPUT39), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(KEYINPUT39), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n636_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT40), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(KEYINPUT40), .B(new_n636_), .C1(new_n638_), .C2(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1325gat));
  INV_X1    g443(.A(G15gat), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n630_), .A2(new_n645_), .A3(new_n379_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT107), .ZN(new_n647_));
  OAI21_X1  g446(.A(G15gat), .B1(new_n619_), .B2(new_n378_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT41), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(KEYINPUT41), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n647_), .A2(new_n649_), .A3(new_n650_), .ZN(G1326gat));
  OAI21_X1  g450(.A(G22gat), .B1(new_n619_), .B2(new_n406_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT42), .ZN(new_n653_));
  INV_X1    g452(.A(G22gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n630_), .A2(new_n654_), .A3(new_n430_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n653_), .A2(new_n655_), .ZN(G1327gat));
  NAND2_X1  g455(.A1(new_n402_), .A2(new_n409_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n431_), .A2(new_n378_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n510_), .A2(new_n553_), .ZN(new_n660_));
  AND4_X1   g459(.A1(new_n617_), .A2(new_n659_), .A3(new_n594_), .A4(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(G29gat), .B1(new_n661_), .B2(new_n399_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT43), .B1(new_n432_), .B2(new_n627_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n659_), .A2(new_n664_), .A3(new_n626_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n616_), .A2(new_n552_), .A3(new_n618_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT44), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670_));
  AOI211_X1 g469(.A(new_n670_), .B(new_n667_), .C1(new_n663_), .C2(new_n665_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n399_), .A2(G29gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n662_), .B1(new_n672_), .B2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(KEYINPUT46), .ZN(new_n675_));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n672_), .B2(new_n635_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n661_), .A2(new_n676_), .A3(new_n635_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT45), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n678_), .B(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n675_), .B1(new_n677_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n678_), .B(KEYINPUT45), .ZN(new_n682_));
  NOR3_X1   g481(.A1(new_n669_), .A2(new_n671_), .A3(new_n403_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n682_), .B(KEYINPUT46), .C1(new_n683_), .C2(new_n676_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(G1329gat));
  AOI21_X1  g484(.A(G43gat), .B1(new_n661_), .B2(new_n379_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n379_), .A2(G43gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n672_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT47), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(G1330gat));
  AOI21_X1  g489(.A(G50gat), .B1(new_n661_), .B2(new_n430_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n430_), .A2(G50gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n691_), .B1(new_n672_), .B2(new_n692_), .ZN(G1331gat));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n659_), .B2(new_n615_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n432_), .A2(KEYINPUT108), .A3(new_n617_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n698_), .A2(new_n594_), .A3(new_n629_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n699_), .A2(new_n530_), .A3(new_n399_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n617_), .A2(new_n552_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n512_), .A2(new_n595_), .A3(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(new_n399_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n700_), .B1(new_n530_), .B2(new_n703_), .ZN(G1332gat));
  AOI21_X1  g503(.A(new_n528_), .B1(new_n702_), .B2(new_n635_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT48), .Z(new_n706_));
  NAND3_X1  g505(.A1(new_n699_), .A2(new_n528_), .A3(new_n635_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1333gat));
  INV_X1    g507(.A(G71gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n699_), .A2(new_n709_), .A3(new_n379_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n702_), .B2(new_n379_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT109), .B(KEYINPUT49), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n711_), .A2(new_n712_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(G1334gat));
  INV_X1    g514(.A(G78gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n716_), .B1(new_n702_), .B2(new_n430_), .ZN(new_n717_));
  XOR2_X1   g516(.A(new_n717_), .B(KEYINPUT50), .Z(new_n718_));
  NAND3_X1  g517(.A1(new_n699_), .A2(new_n716_), .A3(new_n430_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(G1335gat));
  NAND2_X1  g519(.A1(new_n595_), .A2(new_n660_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n697_), .A2(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n451_), .B1(new_n723_), .B2(new_n400_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n725_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n666_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n617_), .A2(new_n553_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n595_), .A2(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n452_), .A2(new_n453_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n400_), .A2(new_n732_), .ZN(new_n733_));
  AOI22_X1  g532(.A1(new_n726_), .A2(new_n727_), .B1(new_n731_), .B2(new_n733_), .ZN(G1336gat));
  NAND3_X1  g533(.A1(new_n697_), .A2(new_n635_), .A3(new_n722_), .ZN(new_n735_));
  INV_X1    g534(.A(G92gat), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n455_), .A2(new_n454_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n403_), .A2(new_n737_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n735_), .A2(new_n736_), .B1(new_n731_), .B2(new_n738_), .ZN(G1337gat));
  NOR3_X1   g538(.A1(new_n728_), .A2(new_n378_), .A3(new_n730_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n379_), .A2(new_n441_), .ZN(new_n741_));
  OAI22_X1  g540(.A1(new_n740_), .A2(new_n472_), .B1(new_n723_), .B2(new_n741_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n742_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g542(.A1(new_n697_), .A2(new_n239_), .A3(new_n430_), .A4(new_n722_), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n666_), .A2(new_n430_), .A3(new_n595_), .A4(new_n729_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(new_n746_), .A3(G106gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(G106gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n744_), .B(new_n750_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1339gat));
  INV_X1    g553(.A(G113gat), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT55), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n756_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n581_), .A2(new_n582_), .A3(KEYINPUT55), .A4(new_n570_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n560_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n563_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n757_), .A2(new_n758_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n587_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT56), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n761_), .A2(KEYINPUT56), .A3(new_n587_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n614_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n596_), .A2(new_n604_), .A3(new_n599_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n603_), .A2(new_n597_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n769_), .A3(new_n611_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n585_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT114), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n771_), .B1(new_n578_), .B2(new_n584_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n766_), .A2(new_n774_), .A3(KEYINPUT58), .A4(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT115), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n764_), .A2(new_n765_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n781_), .A2(KEYINPUT115), .A3(KEYINPUT58), .A4(new_n774_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n761_), .A2(KEYINPUT56), .A3(new_n587_), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT56), .B1(new_n761_), .B2(new_n587_), .ZN(new_n785_));
  OAI22_X1  g584(.A1(new_n773_), .A2(KEYINPUT114), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n775_), .A2(new_n776_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n780_), .A2(new_n626_), .A3(new_n782_), .A4(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n615_), .B1(new_n578_), .B2(new_n584_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n790_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n589_), .A2(new_n772_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n510_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT57), .ZN(new_n795_));
  OAI21_X1  g594(.A(KEYINPUT116), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n511_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(new_n798_), .A3(KEYINPUT57), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n789_), .A2(new_n796_), .A3(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT113), .B1(new_n797_), .B2(KEYINPUT57), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT113), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n771_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n766_), .B2(new_n790_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n802_), .B(new_n795_), .C1(new_n804_), .C2(new_n511_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n801_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n552_), .B1(new_n800_), .B2(new_n806_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n624_), .A2(new_n625_), .A3(new_n701_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT54), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n808_), .B(new_n809_), .C1(new_n591_), .C2(new_n593_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT112), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n594_), .A2(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT54), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n594_), .A2(new_n814_), .A3(new_n809_), .A4(new_n808_), .ZN(new_n815_));
  AND3_X1   g614(.A1(new_n811_), .A2(new_n813_), .A3(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n807_), .A2(new_n817_), .ZN(new_n818_));
  NOR3_X1   g617(.A1(new_n359_), .A2(new_n378_), .A3(new_n400_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n755_), .B1(new_n820_), .B2(new_n615_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n821_), .A2(KEYINPUT117), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(KEYINPUT117), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(KEYINPUT59), .ZN(new_n824_));
  AND4_X1   g623(.A1(new_n798_), .A2(new_n793_), .A3(KEYINPUT57), .A4(new_n510_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n798_), .B1(new_n797_), .B2(KEYINPUT57), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n794_), .A2(new_n795_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n827_), .A2(new_n789_), .A3(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n552_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n817_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n819_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n824_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n617_), .A2(G113gat), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT118), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n822_), .A2(new_n823_), .B1(new_n835_), .B2(new_n837_), .ZN(G1340gat));
  OAI21_X1  g637(.A(G120gat), .B1(new_n834_), .B2(new_n594_), .ZN(new_n839_));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n594_), .B2(KEYINPUT60), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(KEYINPUT60), .B2(new_n840_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n839_), .B1(new_n820_), .B2(new_n842_), .ZN(G1341gat));
  OAI21_X1  g642(.A(G127gat), .B1(new_n834_), .B2(new_n552_), .ZN(new_n844_));
  OR2_X1    g643(.A1(new_n552_), .A2(G127gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n820_), .B2(new_n845_), .ZN(G1342gat));
  INV_X1    g645(.A(G134gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n820_), .B2(new_n510_), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n848_), .A2(KEYINPUT119), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(KEYINPUT119), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT120), .B(G134gat), .Z(new_n851_));
  NOR2_X1   g650(.A1(new_n627_), .A2(new_n851_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n849_), .A2(new_n850_), .B1(new_n835_), .B2(new_n852_), .ZN(G1343gat));
  AOI21_X1  g652(.A(new_n406_), .B1(new_n807_), .B2(new_n817_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n635_), .A2(new_n379_), .A3(new_n400_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n617_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(KEYINPUT122), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n801_), .A2(new_n805_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n827_), .A3(new_n789_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n816_), .B1(new_n859_), .B2(new_n552_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n855_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n860_), .A2(new_n406_), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT122), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n863_), .A3(new_n617_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n857_), .A2(new_n864_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT121), .B(G141gat), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n857_), .A2(new_n864_), .A3(new_n866_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1344gat));
  NAND2_X1  g669(.A1(new_n862_), .A2(new_n595_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g671(.A1(new_n854_), .A2(new_n553_), .A3(new_n855_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(KEYINPUT123), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n862_), .A2(new_n875_), .A3(new_n553_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n874_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n874_), .B2(new_n876_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1346gat));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n881_));
  INV_X1    g680(.A(G162gat), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n862_), .A2(new_n882_), .A3(new_n511_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n882_), .B1(new_n862_), .B2(new_n626_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n881_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n854_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n887_), .A2(new_n627_), .A3(new_n861_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n883_), .B(KEYINPUT124), .C1(new_n888_), .C2(new_n882_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n889_), .ZN(G1347gat));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n816_), .B1(new_n829_), .B2(new_n552_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n403_), .A2(new_n401_), .A3(new_n430_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n892_), .A2(new_n615_), .A3(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n896_));
  OAI21_X1  g695(.A(G169gat), .B1(new_n895_), .B2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n831_), .A2(new_n893_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n898_), .A2(KEYINPUT125), .A3(new_n615_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n891_), .B1(new_n897_), .B2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n895_), .A2(new_n331_), .ZN(new_n901_));
  OAI21_X1  g700(.A(KEYINPUT125), .B1(new_n898_), .B2(new_n615_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n895_), .A2(new_n896_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n902_), .A2(new_n903_), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n900_), .A2(new_n901_), .A3(new_n904_), .ZN(G1348gat));
  NOR2_X1   g704(.A1(new_n892_), .A2(new_n894_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G176gat), .B1(new_n906_), .B2(new_n595_), .ZN(new_n907_));
  NOR4_X1   g706(.A1(new_n860_), .A2(new_n302_), .A3(new_n594_), .A4(new_n894_), .ZN(new_n908_));
  OR3_X1    g707(.A1(new_n907_), .A2(new_n908_), .A3(KEYINPUT126), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT126), .B1(new_n907_), .B2(new_n908_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1349gat));
  NOR3_X1   g710(.A1(new_n898_), .A2(new_n298_), .A3(new_n552_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n818_), .A2(new_n553_), .A3(new_n893_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n285_), .B2(new_n913_), .ZN(G1350gat));
  OAI21_X1  g713(.A(G190gat), .B1(new_n898_), .B2(new_n627_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n906_), .A2(new_n299_), .A3(new_n511_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1351gat));
  NOR2_X1   g716(.A1(new_n379_), .A2(new_n399_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n635_), .A2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n818_), .A2(new_n430_), .A3(new_n920_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(KEYINPUT127), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT127), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n854_), .A2(new_n923_), .A3(new_n920_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(G197gat), .B1(new_n925_), .B2(new_n617_), .ZN(new_n926_));
  AOI211_X1 g725(.A(new_n244_), .B(new_n615_), .C1(new_n922_), .C2(new_n924_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1352gat));
  AOI21_X1  g727(.A(new_n923_), .B1(new_n854_), .B2(new_n920_), .ZN(new_n929_));
  NOR4_X1   g728(.A1(new_n860_), .A2(KEYINPUT127), .A3(new_n406_), .A4(new_n919_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n595_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(G204gat), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n925_), .A2(new_n241_), .A3(new_n595_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(G1353gat));
  XOR2_X1   g733(.A(KEYINPUT63), .B(G211gat), .Z(new_n935_));
  OAI211_X1 g734(.A(new_n553_), .B(new_n935_), .C1(new_n929_), .C2(new_n930_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n552_), .B1(new_n922_), .B2(new_n924_), .ZN(new_n937_));
  OR2_X1    g736(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n936_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n939_), .ZN(G1354gat));
  INV_X1    g739(.A(G218gat), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n925_), .A2(new_n941_), .A3(new_n511_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n627_), .B1(new_n922_), .B2(new_n924_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n941_), .B2(new_n943_), .ZN(G1355gat));
endmodule


