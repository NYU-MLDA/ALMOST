//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n964_,
    new_n965_, new_n966_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT10), .B(G99gat), .Z(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G106gat), .Z(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G85gat), .B(G92gat), .Z(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G99gat), .A2(G106gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT6), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT9), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(G85gat), .A3(G92gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n205_), .A2(new_n207_), .A3(new_n209_), .A4(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT8), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT6), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(KEYINPUT66), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n208_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219_));
  INV_X1    g018(.A(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT7), .B1(new_n221_), .B2(G99gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n219_), .A2(new_n223_), .A3(new_n224_), .A4(new_n220_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n208_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n216_), .A2(KEYINPUT66), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n214_), .A2(KEYINPUT6), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n218_), .A2(new_n222_), .A3(new_n225_), .A4(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n213_), .B1(new_n230_), .B2(new_n206_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n206_), .A2(new_n213_), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n222_), .A2(new_n225_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n232_), .B1(new_n233_), .B2(new_n209_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n212_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G57gat), .B(G64gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT11), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G71gat), .B(G78gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G57gat), .ZN(new_n240_));
  INV_X1    g039(.A(G64gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT11), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G57gat), .A2(G64gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n237_), .A2(new_n239_), .A3(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n236_), .A2(new_n238_), .A3(KEYINPUT11), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n235_), .A2(KEYINPUT12), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n235_), .A2(KEYINPUT67), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n251_), .B(new_n212_), .C1(new_n231_), .C2(new_n234_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n252_), .A3(new_n248_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT12), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n249_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G230gat), .A2(G233gat), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n250_), .A2(new_n252_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n246_), .A2(new_n247_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n257_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n255_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n253_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n248_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n257_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(KEYINPUT69), .B(G204gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(G120gat), .B(G148gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT5), .B(G176gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT68), .ZN(new_n270_));
  XOR2_X1   g069(.A(new_n270_), .B(KEYINPUT70), .Z(new_n271_));
  AND3_X1   g070(.A1(new_n261_), .A2(new_n264_), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n202_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n261_), .A2(new_n264_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n271_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n261_), .A2(new_n264_), .A3(new_n271_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(KEYINPUT13), .A3(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n274_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT85), .ZN(new_n281_));
  XOR2_X1   g080(.A(G127gat), .B(G134gat), .Z(new_n282_));
  INV_X1    g081(.A(G113gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G127gat), .B(G134gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(G113gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G120gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n284_), .A2(G120gat), .A3(new_n286_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G71gat), .B(G99gat), .ZN(new_n292_));
  AND2_X1   g091(.A1(G227gat), .A2(G233gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n291_), .A2(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G15gat), .B(G43gat), .Z(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n289_), .A2(new_n290_), .A3(new_n294_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n296_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n298_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n301_));
  OR2_X1    g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(G183gat), .A3(G190gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT82), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n303_), .B1(G183gat), .B2(G190gat), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n306_), .A2(KEYINPUT81), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(KEYINPUT81), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n305_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G169gat), .ZN(new_n310_));
  INV_X1    g109(.A(G176gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n312_), .A2(KEYINPUT24), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT80), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n316_), .A2(KEYINPUT24), .A3(new_n312_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT25), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT79), .B1(new_n318_), .B2(G183gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT26), .B(G190gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT25), .B(G183gat), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n319_), .B(new_n320_), .C1(new_n321_), .C2(KEYINPUT79), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n309_), .A2(new_n313_), .A3(new_n317_), .A4(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n306_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(new_n304_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT22), .B(G169gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n311_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n328_), .A2(new_n330_), .A3(new_n316_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n323_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n332_), .B1(new_n323_), .B2(new_n331_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n336_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n335_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n339_), .B2(new_n333_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n302_), .A2(new_n337_), .A3(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n300_), .A2(new_n301_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n337_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n336_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n342_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n281_), .B1(new_n341_), .B2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n342_), .A2(new_n344_), .A3(new_n343_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n302_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n348_), .A3(KEYINPUT85), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(G228gat), .ZN(new_n351_));
  INV_X1    g150(.A(G233gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(G197gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(G204gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT89), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT21), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n355_), .A2(G204gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G211gat), .B(G218gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT90), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n358_), .B1(new_n359_), .B2(new_n356_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n360_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n358_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT90), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n361_), .B(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G155gat), .B(G162gat), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n371_), .A2(KEYINPUT1), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G141gat), .A2(G148gat), .ZN(new_n373_));
  NOR2_X1   g172(.A1(G141gat), .A2(G148gat), .ZN(new_n374_));
  AND2_X1   g173(.A1(G155gat), .A2(G162gat), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n375_), .B2(KEYINPUT1), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n372_), .A2(new_n373_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT86), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n374_), .B1(new_n378_), .B2(KEYINPUT3), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n380_), .B(KEYINPUT86), .C1(G141gat), .C2(G148gat), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n379_), .A2(new_n381_), .B1(new_n378_), .B2(KEYINPUT3), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n373_), .B(KEYINPUT2), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n371_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT29), .B1(new_n377_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT88), .ZN(new_n386_));
  AND3_X1   g185(.A1(new_n370_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n386_), .B1(new_n370_), .B2(new_n385_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n354_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n370_), .A2(new_n385_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT88), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n370_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n353_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G78gat), .B(G106gat), .Z(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT91), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n382_), .A2(new_n383_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n371_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n372_), .A2(new_n373_), .A3(new_n376_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n403_), .A2(KEYINPUT29), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G22gat), .B(G50gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n404_), .B(new_n407_), .Z(new_n408_));
  INV_X1    g207(.A(new_n395_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n389_), .A2(new_n393_), .A3(new_n409_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n398_), .A2(new_n408_), .B1(new_n396_), .B2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n396_), .A2(KEYINPUT91), .A3(new_n410_), .A4(new_n408_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n350_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n409_), .B1(new_n389_), .B2(new_n393_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n408_), .B1(new_n415_), .B2(KEYINPUT91), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n396_), .A2(new_n410_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n347_), .A2(new_n348_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n412_), .A3(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n414_), .A2(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT18), .B(G64gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(G92gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G8gat), .B(G36gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n423_), .B(new_n424_), .Z(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(G226gat), .A2(G233gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(new_n427_), .B(KEYINPUT92), .Z(new_n428_));
  XOR2_X1   g227(.A(new_n428_), .B(KEYINPUT19), .Z(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n323_), .A2(new_n365_), .A3(new_n369_), .A4(new_n331_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT20), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(KEYINPUT93), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT93), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(new_n434_), .A3(KEYINPUT20), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n320_), .A2(new_n321_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n312_), .A2(KEYINPUT24), .A3(new_n314_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n325_), .A2(new_n313_), .A3(new_n437_), .A4(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n330_), .A2(new_n316_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT94), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n330_), .A2(new_n316_), .A3(KEYINPUT94), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n309_), .A2(new_n327_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n440_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n370_), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT95), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n309_), .A2(new_n327_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n443_), .A2(new_n444_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n439_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT95), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n452_), .A2(new_n453_), .A3(new_n370_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n449_), .A2(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n430_), .B1(new_n436_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n447_), .A2(new_n448_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT20), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n323_), .A2(new_n331_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n459_), .B2(new_n370_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n460_), .A3(new_n430_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n426_), .B1(new_n456_), .B2(new_n462_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n433_), .A2(new_n435_), .B1(new_n449_), .B2(new_n454_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n425_), .B(new_n461_), .C1(new_n464_), .C2(new_n430_), .ZN(new_n465_));
  AOI21_X1  g264(.A(KEYINPUT27), .B1(new_n463_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT101), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n465_), .B(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT27), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT99), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n452_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n447_), .A2(KEYINPUT99), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n448_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n430_), .B1(new_n473_), .B2(new_n460_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n436_), .A2(new_n455_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n475_), .B1(new_n429_), .B2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n469_), .B1(new_n477_), .B2(new_n426_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n466_), .B1(new_n468_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n290_), .ZN(new_n480_));
  AOI21_X1  g279(.A(G120gat), .B1(new_n284_), .B2(new_n286_), .ZN(new_n481_));
  OAI22_X1  g280(.A1(new_n377_), .A2(new_n384_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(KEYINPUT96), .B1(new_n482_), .B2(KEYINPUT4), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n401_), .A2(new_n289_), .A3(new_n402_), .A4(new_n290_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n484_), .A3(KEYINPUT4), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT96), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT4), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n403_), .A2(new_n291_), .A3(new_n486_), .A4(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n483_), .A2(new_n485_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G225gat), .A2(G233gat), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n491_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT0), .B(G57gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(G85gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(G1gat), .B(G29gat), .Z(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT100), .B1(new_n495_), .B2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n495_), .A2(new_n500_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n493_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT100), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n504_), .A3(new_n499_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n502_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n421_), .A2(new_n479_), .A3(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n411_), .A2(new_n413_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n425_), .A2(KEYINPUT32), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n476_), .A2(new_n429_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n511_), .B1(new_n512_), .B2(new_n474_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n461_), .B(new_n510_), .C1(new_n464_), .C2(new_n430_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT98), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n476_), .A2(new_n429_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n517_), .A2(KEYINPUT98), .A3(new_n461_), .A4(new_n510_), .ZN(new_n518_));
  AND4_X1   g317(.A1(new_n506_), .A2(new_n513_), .A3(new_n516_), .A4(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n463_), .A2(new_n465_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT33), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT97), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n495_), .A2(new_n500_), .A3(new_n522_), .ZN(new_n523_));
  OAI211_X1 g322(.A(KEYINPUT97), .B(new_n521_), .C1(new_n503_), .C2(new_n499_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n489_), .A2(new_n491_), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n482_), .A2(new_n484_), .A3(new_n491_), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n526_), .A2(new_n500_), .A3(new_n527_), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n520_), .A2(new_n525_), .A3(new_n528_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n509_), .B(new_n350_), .C1(new_n519_), .C2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n508_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G113gat), .B(G141gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(new_n310_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(G197gat), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(KEYINPUT78), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT77), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537_));
  NAND2_X1  g336(.A1(G1gat), .A2(G8gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT14), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(G1gat), .ZN(new_n541_));
  INV_X1    g340(.A(G8gat), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n538_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n544_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n537_), .A2(new_n538_), .A3(new_n543_), .A4(new_n539_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(G29gat), .ZN(new_n548_));
  INV_X1    g347(.A(G36gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(G43gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G29gat), .A2(G36gat), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(G50gat), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n551_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G29gat), .B(G36gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(G43gat), .ZN(new_n559_));
  AOI21_X1  g358(.A(G50gat), .B1(new_n559_), .B2(new_n553_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT15), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n557_), .A2(new_n560_), .A3(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n555_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n559_), .A2(G50gat), .A3(new_n553_), .ZN(new_n564_));
  AOI21_X1  g363(.A(KEYINPUT15), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n547_), .B1(new_n562_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G229gat), .A2(G233gat), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n563_), .A2(new_n545_), .A3(new_n564_), .A4(new_n546_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n563_), .A2(new_n564_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n570_), .A2(new_n547_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n567_), .B1(new_n571_), .B2(new_n568_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n536_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n572_), .A2(KEYINPUT77), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n535_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n535_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n575_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n568_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n561_), .B1(new_n557_), .B2(new_n560_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n563_), .A2(KEYINPUT15), .A3(new_n564_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n579_), .B1(new_n582_), .B2(new_n547_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n572_), .B1(new_n583_), .B2(new_n567_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n577_), .B(new_n578_), .C1(new_n584_), .C2(new_n536_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n576_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n531_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT102), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n531_), .A2(KEYINPUT102), .A3(new_n586_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n280_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n570_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT34), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT35), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(KEYINPUT35), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n235_), .A2(new_n582_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n593_), .A2(new_n596_), .A3(new_n597_), .A4(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n598_), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT35), .B(new_n595_), .C1(new_n592_), .C2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G190gat), .B(G218gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(G134gat), .ZN(new_n604_));
  INV_X1    g403(.A(G162gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n607_), .A2(KEYINPUT36), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(KEYINPUT36), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n602_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n611_), .A2(KEYINPUT71), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n599_), .A2(new_n608_), .A3(new_n601_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(KEYINPUT71), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n612_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n611_), .A2(new_n613_), .ZN(new_n616_));
  OAI21_X1  g415(.A(KEYINPUT72), .B1(new_n616_), .B2(KEYINPUT37), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT72), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT37), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n611_), .A2(new_n618_), .A3(new_n619_), .A4(new_n613_), .ZN(new_n620_));
  AOI22_X1  g419(.A1(new_n615_), .A2(KEYINPUT37), .B1(new_n617_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(G231gat), .A2(G233gat), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n545_), .A2(new_n546_), .A3(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n622_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n259_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n622_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n547_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n545_), .A2(new_n546_), .A3(new_n622_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n627_), .A2(new_n248_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT73), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n625_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n630_), .B1(new_n625_), .B2(new_n629_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G127gat), .B(G155gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G183gat), .B(G211gat), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n635_), .A2(new_n637_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT17), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n631_), .A2(new_n632_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n625_), .A2(new_n629_), .A3(KEYINPUT75), .ZN(new_n643_));
  OR3_X1    g442(.A1(new_n638_), .A2(new_n639_), .A3(KEYINPUT17), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n640_), .ZN(new_n645_));
  AOI21_X1  g444(.A(KEYINPUT75), .B1(new_n625_), .B2(new_n629_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT76), .B1(new_n645_), .B2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n643_), .A2(new_n644_), .A3(new_n640_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT76), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n646_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n642_), .B1(new_n648_), .B2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n621_), .A2(new_n652_), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n591_), .A2(new_n541_), .A3(new_n506_), .A4(new_n653_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(KEYINPUT103), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(KEYINPUT103), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT38), .ZN(new_n657_));
  OR3_X1    g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n616_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(new_n652_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n531_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n586_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n280_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT104), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(new_n506_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G1gat), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n657_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n658_), .A2(new_n667_), .A3(new_n668_), .ZN(G1324gat));
  INV_X1    g468(.A(new_n479_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n591_), .A2(new_n542_), .A3(new_n670_), .A4(new_n653_), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n531_), .A2(new_n663_), .A3(new_n670_), .A4(new_n660_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(G8gat), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT39), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n673_), .A2(new_n674_), .A3(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n673_), .A2(new_n674_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n672_), .A2(KEYINPUT105), .A3(G8gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(KEYINPUT39), .A3(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n671_), .A2(new_n676_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT106), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT106), .ZN(new_n682_));
  NAND4_X1  g481(.A1(new_n671_), .A2(new_n679_), .A3(new_n682_), .A4(new_n676_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n681_), .A2(KEYINPUT40), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT40), .B1(new_n681_), .B2(new_n683_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1325gat));
  INV_X1    g485(.A(G15gat), .ZN(new_n687_));
  INV_X1    g486(.A(new_n350_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n665_), .B2(new_n688_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n689_), .B(KEYINPUT41), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n591_), .A2(new_n653_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n692_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n690_), .A2(new_n693_), .ZN(G1326gat));
  INV_X1    g493(.A(G22gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n509_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n665_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n692_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1327gat));
  INV_X1    g500(.A(new_n280_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n645_), .A2(KEYINPUT76), .A3(new_n647_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n650_), .B1(new_n649_), .B2(new_n646_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n641_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n616_), .A2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT102), .B1(new_n531_), .B2(new_n586_), .ZN(new_n707_));
  AOI211_X1 g506(.A(new_n588_), .B(new_n662_), .C1(new_n508_), .C2(new_n530_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n702_), .B(new_n706_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G29gat), .B1(new_n710_), .B2(new_n506_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n531_), .A2(new_n712_), .A3(new_n621_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n712_), .B1(new_n531_), .B2(new_n621_), .ZN(new_n715_));
  OAI211_X1 g514(.A(new_n663_), .B(new_n652_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n715_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n713_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n720_), .A2(KEYINPUT44), .A3(new_n663_), .A4(new_n652_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n718_), .A2(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n507_), .A2(new_n548_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n711_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  NAND3_X1  g523(.A1(new_n718_), .A2(new_n721_), .A3(new_n670_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(G36gat), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n479_), .B(KEYINPUT107), .Z(new_n727_));
  NAND4_X1  g526(.A1(new_n591_), .A2(new_n549_), .A3(new_n706_), .A4(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT45), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT45), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n710_), .A2(new_n730_), .A3(new_n549_), .A4(new_n727_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n726_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT46), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n726_), .A2(new_n732_), .A3(KEYINPUT46), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1329gat));
  NAND4_X1  g536(.A1(new_n718_), .A2(new_n721_), .A3(G43gat), .A4(new_n419_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT108), .B(G43gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n739_), .B1(new_n709_), .B2(new_n350_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n741_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g541(.A(G50gat), .B1(new_n710_), .B2(new_n696_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n509_), .A2(new_n555_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n722_), .B2(new_n744_), .ZN(G1331gat));
  AOI21_X1  g544(.A(new_n240_), .B1(new_n506_), .B2(KEYINPUT110), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n702_), .A2(new_n586_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n661_), .A2(new_n747_), .ZN(new_n748_));
  AOI211_X1 g547(.A(new_n746_), .B(new_n748_), .C1(KEYINPUT110), .C2(new_n240_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n653_), .A2(KEYINPUT109), .A3(new_n280_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n662_), .A3(new_n531_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT109), .B1(new_n653_), .B2(new_n280_), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n753_), .A2(new_n507_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n749_), .B1(new_n754_), .B2(new_n240_), .ZN(G1332gat));
  INV_X1    g554(.A(new_n727_), .ZN(new_n756_));
  OAI21_X1  g555(.A(G64gat), .B1(new_n748_), .B2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT48), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n727_), .A2(new_n241_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n753_), .B2(new_n759_), .ZN(G1333gat));
  OAI21_X1  g559(.A(G71gat), .B1(new_n748_), .B2(new_n350_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT49), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n350_), .A2(G71gat), .ZN(new_n763_));
  XOR2_X1   g562(.A(new_n763_), .B(KEYINPUT111), .Z(new_n764_));
  OAI21_X1  g563(.A(new_n762_), .B1(new_n753_), .B2(new_n764_), .ZN(G1334gat));
  OAI21_X1  g564(.A(G78gat), .B1(new_n748_), .B2(new_n509_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT50), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n509_), .A2(G78gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n753_), .B2(new_n768_), .ZN(G1335gat));
  NAND3_X1  g568(.A1(new_n531_), .A2(new_n706_), .A3(new_n747_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(G85gat), .B1(new_n771_), .B2(new_n506_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n720_), .A2(new_n652_), .A3(new_n747_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n773_), .A2(new_n507_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n774_), .B2(G85gat), .ZN(G1336gat));
  INV_X1    g574(.A(G92gat), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n773_), .A2(new_n776_), .A3(new_n756_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n770_), .B2(new_n479_), .ZN(new_n778_));
  XOR2_X1   g577(.A(new_n778_), .B(KEYINPUT112), .Z(new_n779_));
  NOR2_X1   g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1337gat));
  OAI21_X1  g579(.A(G99gat), .B1(new_n773_), .B2(new_n350_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n771_), .A2(new_n203_), .A3(new_n419_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g583(.A1(new_n720_), .A2(new_n696_), .A3(new_n652_), .A4(new_n747_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT52), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(G106gat), .A3(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n786_), .A2(KEYINPUT52), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n771_), .A2(new_n204_), .A3(new_n696_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n789_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n785_), .A2(G106gat), .A3(new_n792_), .A4(new_n787_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n790_), .A2(new_n791_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(KEYINPUT53), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n790_), .A2(new_n796_), .A3(new_n791_), .A4(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1339gat));
  INV_X1    g597(.A(KEYINPUT114), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n799_), .B1(new_n652_), .B2(new_n586_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n705_), .A2(KEYINPUT114), .A3(new_n576_), .A4(new_n585_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT115), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n802_), .A2(new_n803_), .A3(new_n279_), .A4(new_n274_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n800_), .A2(new_n801_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT115), .B1(new_n280_), .B2(new_n805_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n615_), .A2(KEYINPUT37), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n617_), .A2(new_n620_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(KEYINPUT116), .A2(KEYINPUT54), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n807_), .A2(new_n810_), .A3(new_n813_), .A4(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n804_), .A2(new_n806_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n811_), .B(new_n812_), .C1(new_n816_), .C2(new_n621_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT57), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n574_), .A2(new_n575_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n583_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n583_), .A2(new_n821_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n822_), .A2(G229gat), .A3(G233gat), .A4(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n571_), .A2(new_n568_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n534_), .B1(new_n825_), .B2(new_n567_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n826_), .B(new_n827_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n534_), .A2(new_n820_), .B1(new_n824_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT120), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n829_), .B(KEYINPUT120), .C1(new_n272_), .C2(new_n273_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n255_), .A2(KEYINPUT55), .A3(new_n260_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n258_), .A2(new_n259_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n256_), .B1(new_n255_), .B2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT55), .B1(new_n255_), .B2(new_n260_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n836_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n269_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n835_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n261_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n253_), .A2(new_n254_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n249_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n837_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n257_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n255_), .A2(KEYINPUT55), .A3(new_n260_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n845_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n843_), .B1(new_n851_), .B2(new_n269_), .ZN(new_n852_));
  AOI22_X1  g651(.A1(new_n842_), .A2(new_n843_), .B1(new_n852_), .B2(new_n835_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n261_), .A2(new_n264_), .A3(new_n841_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n854_), .A2(new_n586_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n834_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n819_), .B1(new_n856_), .B2(new_n659_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT121), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT56), .B1(new_n840_), .B2(new_n841_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n851_), .A2(new_n843_), .A3(new_n269_), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n859_), .A2(new_n854_), .A3(new_n829_), .A4(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n858_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n860_), .A2(new_n854_), .A3(new_n829_), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n864_), .A2(KEYINPUT121), .A3(KEYINPUT58), .A4(new_n859_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n861_), .A2(new_n862_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n863_), .A2(new_n621_), .A3(new_n865_), .A4(new_n866_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n835_), .B(KEYINPUT56), .C1(new_n840_), .C2(new_n841_), .ZN(new_n868_));
  AOI21_X1  g667(.A(KEYINPUT117), .B1(new_n851_), .B2(new_n269_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n868_), .B(new_n855_), .C1(KEYINPUT56), .C2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n834_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n872_), .A2(KEYINPUT57), .A3(new_n616_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n857_), .A2(new_n867_), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n818_), .B1(new_n652_), .B2(new_n874_), .ZN(new_n875_));
  NOR4_X1   g674(.A1(new_n875_), .A2(new_n507_), .A3(new_n420_), .A4(new_n670_), .ZN(new_n876_));
  AOI21_X1  g675(.A(G113gat), .B1(new_n876_), .B2(new_n586_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT59), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n878_), .B1(new_n875_), .B2(KEYINPUT122), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n874_), .A2(new_n652_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n818_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT122), .ZN(new_n884_));
  AOI21_X1  g683(.A(KEYINPUT59), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n420_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n883_), .A2(new_n506_), .A3(new_n886_), .A4(new_n479_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n662_), .B1(new_n880_), .B2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n877_), .B1(new_n889_), .B2(G113gat), .ZN(G1340gat));
  OAI21_X1  g689(.A(new_n288_), .B1(new_n702_), .B2(KEYINPUT60), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n876_), .B(new_n891_), .C1(KEYINPUT60), .C2(new_n288_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n702_), .B1(new_n880_), .B2(new_n888_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n288_), .ZN(G1341gat));
  AOI21_X1  g693(.A(G127gat), .B1(new_n876_), .B2(new_n705_), .ZN(new_n895_));
  INV_X1    g694(.A(G127gat), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n896_), .B1(new_n880_), .B2(new_n888_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n897_), .B2(new_n705_), .ZN(G1342gat));
  AOI21_X1  g697(.A(G134gat), .B1(new_n876_), .B2(new_n659_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n880_), .A2(new_n888_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n621_), .A2(G134gat), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT123), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n899_), .B1(new_n900_), .B2(new_n902_), .ZN(G1343gat));
  NOR2_X1   g702(.A1(new_n875_), .A2(new_n507_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n414_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n904_), .A2(new_n586_), .A3(new_n905_), .A4(new_n756_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g706(.A1(new_n904_), .A2(new_n280_), .A3(new_n905_), .A4(new_n756_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g708(.A1(new_n904_), .A2(new_n905_), .A3(new_n756_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n910_), .A2(new_n652_), .ZN(new_n911_));
  XOR2_X1   g710(.A(KEYINPUT61), .B(G155gat), .Z(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1346gat));
  NOR3_X1   g712(.A1(new_n910_), .A2(new_n605_), .A3(new_n810_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n910_), .A2(new_n616_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n605_), .B2(new_n915_), .ZN(G1347gat));
  NAND2_X1  g715(.A1(new_n727_), .A2(new_n507_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n883_), .A2(new_n509_), .A3(new_n688_), .A4(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(G169gat), .B1(new_n919_), .B2(new_n662_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(KEYINPUT62), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n922_), .B(G169gat), .C1(new_n919_), .C2(new_n662_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n875_), .A2(new_n696_), .A3(new_n917_), .ZN(new_n925_));
  AOI21_X1  g724(.A(KEYINPUT124), .B1(new_n925_), .B2(new_n688_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n917_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n927_));
  AND4_X1   g726(.A1(KEYINPUT124), .A2(new_n927_), .A3(new_n509_), .A4(new_n688_), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n586_), .B(new_n329_), .C1(new_n926_), .C2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n924_), .A2(new_n929_), .ZN(G1348gat));
  OAI211_X1 g729(.A(new_n311_), .B(new_n280_), .C1(new_n926_), .C2(new_n928_), .ZN(new_n931_));
  OAI21_X1  g730(.A(G176gat), .B1(new_n919_), .B2(new_n702_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1349gat));
  NOR2_X1   g732(.A1(new_n919_), .A2(new_n652_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(G183gat), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n919_), .A2(new_n936_), .ZN(new_n937_));
  NAND4_X1  g736(.A1(new_n927_), .A2(KEYINPUT124), .A3(new_n509_), .A4(new_n688_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n321_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n935_), .B1(new_n705_), .B2(new_n939_), .ZN(G1350gat));
  OAI21_X1  g739(.A(new_n320_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n810_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n942_));
  INV_X1    g741(.A(G190gat), .ZN(new_n943_));
  OAI22_X1  g742(.A1(new_n941_), .A2(new_n616_), .B1(new_n942_), .B2(new_n943_), .ZN(G1351gat));
  NOR3_X1   g743(.A1(new_n875_), .A2(new_n414_), .A3(new_n917_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n945_), .A2(new_n586_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n280_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g748(.A(new_n652_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n950_), .A2(KEYINPUT125), .ZN(new_n951_));
  OR2_X1    g750(.A1(new_n950_), .A2(KEYINPUT125), .ZN(new_n952_));
  NAND4_X1  g751(.A1(new_n927_), .A2(new_n905_), .A3(new_n951_), .A4(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(KEYINPUT126), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955_));
  NAND4_X1  g754(.A1(new_n945_), .A2(new_n955_), .A3(new_n951_), .A4(new_n952_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n954_), .A2(new_n956_), .ZN(new_n957_));
  INV_X1    g756(.A(KEYINPUT63), .ZN(new_n958_));
  INV_X1    g757(.A(G211gat), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n957_), .A2(new_n960_), .ZN(new_n961_));
  NAND4_X1  g760(.A1(new_n954_), .A2(new_n956_), .A3(new_n958_), .A4(new_n959_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n961_), .A2(new_n962_), .ZN(G1354gat));
  NAND2_X1  g762(.A1(new_n945_), .A2(new_n659_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(KEYINPUT127), .B(G218gat), .ZN(new_n965_));
  NOR4_X1   g764(.A1(new_n875_), .A2(new_n414_), .A3(new_n917_), .A4(new_n965_), .ZN(new_n966_));
  AOI22_X1  g765(.A1(new_n964_), .A2(new_n965_), .B1(new_n966_), .B2(new_n621_), .ZN(G1355gat));
endmodule


