//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n955_, new_n956_, new_n958_, new_n959_, new_n960_,
    new_n961_, new_n963_, new_n964_, new_n966_, new_n967_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT22), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G169gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT22), .ZN(new_n213_));
  INV_X1    g012(.A(G176gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n211_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G169gat), .A2(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT99), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n220_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT23), .ZN(new_n223_));
  NOR2_X1   g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n221_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT99), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n215_), .A2(new_n227_), .A3(new_n216_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n218_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G183gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n230_), .A2(KEYINPUT25), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(G183gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT26), .B(G190gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n220_), .A2(KEYINPUT23), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT23), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT83), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT83), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT23), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n237_), .B1(new_n242_), .B2(new_n220_), .ZN(new_n243_));
  OR3_X1    g042(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n212_), .A2(new_n214_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(KEYINPUT24), .A3(new_n216_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n236_), .A2(new_n243_), .A3(new_n244_), .A4(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G204gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(G197gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(KEYINPUT93), .B(G204gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(new_n250_), .B2(G197gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT21), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT21), .ZN(new_n253_));
  INV_X1    g052(.A(G197gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n248_), .A2(KEYINPUT93), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT93), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(G204gat), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n254_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(G197gat), .A2(G204gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n253_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G211gat), .B(G218gat), .ZN(new_n261_));
  AND3_X1   g060(.A1(new_n252_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n253_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(KEYINPUT94), .B1(new_n258_), .B2(new_n259_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT94), .ZN(new_n266_));
  INV_X1    g065(.A(new_n259_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n266_), .B(new_n267_), .C1(new_n250_), .C2(new_n254_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n264_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n229_), .B(new_n247_), .C1(new_n262_), .C2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT84), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n271_), .B1(new_n212_), .B2(KEYINPUT22), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n214_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT85), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(G176gat), .B1(new_n211_), .B2(new_n271_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT85), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT22), .B(G169gat), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n276_), .B(new_n277_), .C1(new_n271_), .C2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n275_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n238_), .B1(G183gat), .B2(G190gat), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(new_n219_), .B2(new_n222_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n216_), .B1(new_n282_), .B2(new_n224_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n280_), .A2(new_n283_), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n221_), .A2(new_n223_), .A3(new_n244_), .A4(new_n246_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT82), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT81), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n287_), .A2(KEYINPUT26), .A3(G190gat), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT26), .B1(new_n287_), .B2(G190gat), .ZN(new_n289_));
  OAI22_X1  g088(.A1(new_n288_), .A2(new_n289_), .B1(KEYINPUT80), .B2(new_n231_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT80), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n232_), .A2(G183gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n230_), .A2(KEYINPUT25), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n286_), .B1(new_n290_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT26), .ZN(new_n296_));
  INV_X1    g095(.A(G190gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n296_), .B1(new_n297_), .B2(KEYINPUT81), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n287_), .A2(KEYINPUT26), .A3(G190gat), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n298_), .A2(new_n299_), .B1(new_n292_), .B2(new_n291_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT80), .B1(new_n231_), .B2(new_n233_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n300_), .A2(new_n301_), .A3(KEYINPUT82), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n285_), .B1(new_n295_), .B2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n284_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n265_), .A2(new_n268_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n263_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n252_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n270_), .B1(new_n304_), .B2(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n209_), .B1(new_n309_), .B2(KEYINPUT20), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n229_), .A2(new_n247_), .ZN(new_n311_));
  OAI211_X1 g110(.A(KEYINPUT20), .B(new_n209_), .C1(new_n308_), .C2(new_n311_), .ZN(new_n312_));
  OAI22_X1  g111(.A1(new_n284_), .A2(new_n303_), .B1(new_n262_), .B2(new_n269_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT100), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  AND4_X1   g114(.A1(new_n221_), .A2(new_n223_), .A3(new_n244_), .A4(new_n246_), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n300_), .A2(new_n301_), .A3(KEYINPUT82), .ZN(new_n317_));
  AOI21_X1  g116(.A(KEYINPUT82), .B1(new_n300_), .B2(new_n301_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n243_), .A2(new_n225_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n320_), .A2(new_n216_), .A3(new_n275_), .A4(new_n279_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(new_n308_), .A3(KEYINPUT100), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n312_), .B1(new_n315_), .B2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n206_), .B1(new_n310_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n209_), .A2(KEYINPUT20), .ZN(new_n326_));
  INV_X1    g125(.A(new_n308_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n311_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n326_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n322_), .A2(new_n308_), .A3(KEYINPUT100), .ZN(new_n330_));
  AOI21_X1  g129(.A(KEYINPUT100), .B1(new_n322_), .B2(new_n308_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT20), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n327_), .A2(new_n322_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n334_), .B2(new_n270_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n332_), .B(new_n205_), .C1(new_n209_), .C2(new_n335_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n325_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT102), .B(KEYINPUT27), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT96), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n308_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n306_), .A2(new_n307_), .A3(KEYINPUT96), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n333_), .B1(new_n343_), .B2(new_n328_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n315_), .A2(new_n323_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n209_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n335_), .A2(new_n209_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n206_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n348_), .A2(KEYINPUT27), .A3(new_n336_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G1gat), .B(G29gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT0), .ZN(new_n351_));
  INV_X1    g150(.A(G57gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(G85gat), .ZN(new_n354_));
  INV_X1    g153(.A(G155gat), .ZN(new_n355_));
  INV_X1    g154(.A(G162gat), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT1), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(G155gat), .A3(G162gat), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n356_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(G141gat), .ZN(new_n362_));
  INV_X1    g161(.A(G148gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G141gat), .A2(G148gat), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(KEYINPUT88), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT88), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n361_), .A2(new_n369_), .A3(new_n366_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n364_), .A2(KEYINPUT3), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n365_), .A2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n372_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT89), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n378_), .A2(G141gat), .A3(G148gat), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT89), .B1(new_n362_), .B2(new_n363_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n377_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT90), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n362_), .A2(new_n363_), .A3(KEYINPUT89), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n378_), .B1(G141gat), .B2(G148gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(KEYINPUT90), .A3(new_n377_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n376_), .B1(new_n383_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n360_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n355_), .A2(new_n356_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n371_), .B1(new_n388_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT91), .ZN(new_n394_));
  XOR2_X1   g193(.A(G127gat), .B(G134gat), .Z(new_n395_));
  XNOR2_X1  g194(.A(G113gat), .B(G120gat), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n395_), .A2(new_n396_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n376_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT90), .B1(new_n386_), .B2(new_n377_), .ZN(new_n402_));
  AOI211_X1 g201(.A(new_n382_), .B(KEYINPUT3), .C1(new_n384_), .C2(new_n385_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n401_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n391_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT91), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n371_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n394_), .A2(new_n400_), .A3(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n400_), .A2(KEYINPUT101), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT101), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n399_), .A2(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n371_), .B(new_n405_), .C1(new_n410_), .C2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n408_), .A2(new_n409_), .A3(new_n413_), .ZN(new_n414_));
  AND3_X1   g213(.A1(new_n408_), .A2(KEYINPUT4), .A3(new_n413_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n394_), .A2(new_n416_), .A3(new_n400_), .A4(new_n407_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n409_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n354_), .B(new_n414_), .C1(new_n415_), .C2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n408_), .A2(new_n413_), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n418_), .B(new_n417_), .C1(new_n422_), .C2(new_n416_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n354_), .B1(new_n423_), .B2(new_n414_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n421_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n339_), .A2(new_n349_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n428_));
  XOR2_X1   g227(.A(G22gat), .B(G50gat), .Z(new_n429_));
  NAND2_X1  g228(.A1(new_n394_), .A2(new_n407_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT29), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n429_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n429_), .ZN(new_n433_));
  AOI211_X1 g232(.A(KEYINPUT29), .B(new_n433_), .C1(new_n394_), .C2(new_n407_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n428_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n405_), .A2(new_n406_), .A3(new_n371_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n406_), .B1(new_n405_), .B2(new_n371_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n431_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(new_n433_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n430_), .A2(new_n431_), .A3(new_n429_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n428_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n435_), .A2(KEYINPUT97), .A3(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G78gat), .B(G106gat), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n435_), .A2(new_n442_), .A3(KEYINPUT97), .A4(new_n444_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT97), .B1(new_n435_), .B2(new_n442_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n327_), .B1(G228gat), .B2(G233gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n450_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT95), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n431_), .B1(new_n405_), .B2(new_n371_), .ZN(new_n453_));
  OAI211_X1 g252(.A(G228gat), .B(G233gat), .C1(new_n343_), .C2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT95), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n450_), .B(new_n455_), .C1(new_n430_), .C2(new_n431_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n452_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n449_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n448_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT30), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(new_n284_), .B2(new_n303_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G15gat), .B(G43gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT86), .ZN(new_n463_));
  XOR2_X1   g262(.A(G71gat), .B(G99gat), .Z(new_n464_));
  NAND2_X1  g263(.A1(G227gat), .A2(G233gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n463_), .B(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n319_), .A2(new_n321_), .A3(KEYINPUT30), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n461_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n461_), .B2(new_n468_), .ZN(new_n470_));
  OAI21_X1  g269(.A(KEYINPUT31), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n467_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n468_), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT30), .B1(new_n319_), .B2(new_n321_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n472_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT31), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n461_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  AND3_X1   g277(.A1(new_n471_), .A2(new_n399_), .A3(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n399_), .B1(new_n471_), .B2(new_n478_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT87), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NOR3_X1   g282(.A1(new_n469_), .A2(new_n470_), .A3(KEYINPUT31), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n476_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n400_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n471_), .A2(new_n478_), .A3(new_n399_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n482_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n483_), .A2(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n446_), .B(new_n447_), .C1(new_n449_), .C2(new_n457_), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n459_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n486_), .A2(new_n487_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n493_), .B1(new_n459_), .B2(new_n491_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n427_), .B1(new_n492_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n459_), .A2(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n498_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n332_), .B(new_n497_), .C1(new_n209_), .C2(new_n335_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n499_), .B(new_n500_), .C1(new_n421_), .C2(new_n424_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT33), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n420_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n422_), .A2(new_n418_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n408_), .A2(KEYINPUT4), .A3(new_n409_), .A4(new_n413_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n417_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n354_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n423_), .A2(KEYINPUT33), .A3(new_n354_), .A4(new_n414_), .ZN(new_n509_));
  NAND4_X1  g308(.A1(new_n503_), .A2(new_n337_), .A3(new_n508_), .A4(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n501_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n496_), .A2(new_n490_), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n495_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G230gat), .A2(G233gat), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT68), .B(G71gat), .ZN(new_n516_));
  INV_X1    g315(.A(G78gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G57gat), .B(G64gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT11), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n516_), .B(G78gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(KEYINPUT11), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT10), .B(G99gat), .Z(new_n526_));
  INV_X1    g325(.A(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT64), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G99gat), .A2(G106gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT6), .ZN(new_n531_));
  INV_X1    g330(.A(G85gat), .ZN(new_n532_));
  INV_X1    g331(.A(G92gat), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT65), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  AOI22_X1  g333(.A1(new_n534_), .A2(KEYINPUT9), .B1(new_n532_), .B2(new_n533_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n535_), .B1(KEYINPUT9), .B2(new_n534_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n529_), .A2(new_n531_), .A3(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G85gat), .B(G92gat), .ZN(new_n538_));
  NOR3_X1   g337(.A1(KEYINPUT66), .A2(G99gat), .A3(G106gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT7), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n540_), .B2(new_n531_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n541_), .A2(KEYINPUT8), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n537_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n538_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT8), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n540_), .B(KEYINPUT67), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n545_), .B1(new_n546_), .B2(new_n531_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n525_), .B1(new_n543_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT69), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n543_), .A2(new_n547_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n525_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n554_), .B1(new_n549_), .B2(KEYINPUT69), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n515_), .B1(new_n551_), .B2(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n543_), .A2(new_n547_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n525_), .B(KEYINPUT70), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(KEYINPUT12), .A3(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT12), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n548_), .A2(new_n560_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n559_), .A2(new_n561_), .A3(new_n514_), .A4(new_n554_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n556_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G120gat), .B(G148gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT5), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G176gat), .B(G204gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT71), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n563_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n567_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n556_), .A2(new_n562_), .A3(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT13), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G113gat), .B(G141gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G169gat), .B(G197gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G229gat), .A2(G233gat), .ZN(new_n579_));
  XOR2_X1   g378(.A(KEYINPUT74), .B(KEYINPUT15), .Z(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT14), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT77), .B(G1gat), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n582_), .B1(new_n583_), .B2(G8gat), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT78), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G15gat), .B(G22gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G1gat), .B(G8gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G29gat), .B(G36gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G43gat), .B(G50gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n589_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n588_), .B(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n593_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n581_), .B1(new_n595_), .B2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n593_), .A2(new_n580_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n579_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n595_), .A2(new_n598_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n579_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AOI211_X1 g403(.A(KEYINPUT79), .B(new_n578_), .C1(new_n601_), .C2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT79), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n601_), .A2(new_n604_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n607_), .B2(new_n577_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n601_), .A2(new_n578_), .A3(new_n604_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n605_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n574_), .A2(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n513_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G232gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT35), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT73), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n557_), .A2(new_n594_), .A3(new_n580_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n616_), .A2(KEYINPUT35), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n580_), .B1(new_n543_), .B2(new_n547_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n620_), .B1(new_n621_), .B2(new_n593_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n618_), .B1(new_n619_), .B2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(new_n622_), .A3(new_n618_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT75), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT75), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n619_), .A2(new_n622_), .A3(new_n626_), .A4(new_n618_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n623_), .B1(new_n625_), .B2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(G190gat), .B(G218gat), .Z(new_n629_));
  XNOR2_X1  g428(.A(G134gat), .B(G162gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n629_), .B(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n632_), .A2(KEYINPUT36), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n628_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT76), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT37), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n631_), .B(KEYINPUT36), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  OAI221_X1 g437(.A(new_n634_), .B1(new_n635_), .B2(new_n636_), .C1(new_n628_), .C2(new_n638_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n635_), .B1(new_n628_), .B2(new_n638_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n628_), .A2(new_n638_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n633_), .ZN(new_n642_));
  AOI211_X1 g441(.A(new_n623_), .B(new_n642_), .C1(new_n625_), .C2(new_n627_), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n640_), .B(KEYINPUT37), .C1(new_n641_), .C2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n639_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(G231gat), .A2(G233gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n590_), .B(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(new_n558_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT17), .ZN(new_n651_));
  XOR2_X1   g450(.A(G127gat), .B(G155gat), .Z(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT16), .ZN(new_n653_));
  XNOR2_X1  g452(.A(G183gat), .B(G211gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n650_), .A2(new_n651_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT70), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n525_), .B(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n656_), .B1(new_n658_), .B2(new_n648_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n649_), .A2(new_n553_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n648_), .A2(new_n525_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n655_), .B(KEYINPUT17), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n659_), .A2(new_n663_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n646_), .A2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n613_), .A2(new_n665_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n666_), .A2(new_n425_), .A3(new_n583_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT38), .Z(new_n668_));
  NOR2_X1   g467(.A1(new_n641_), .A2(new_n643_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT103), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n513_), .A2(KEYINPUT104), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(KEYINPUT104), .B1(new_n513_), .B2(new_n670_), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n574_), .A2(new_n611_), .A3(new_n664_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G1gat), .B1(new_n675_), .B2(new_n425_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n668_), .A2(new_n676_), .ZN(G1324gat));
  NAND2_X1  g476(.A1(new_n339_), .A2(new_n349_), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n678_), .B(new_n674_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(G8gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT105), .B1(new_n680_), .B2(KEYINPUT39), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT39), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n679_), .A2(new_n682_), .A3(new_n683_), .A4(G8gat), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n680_), .A2(KEYINPUT39), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n681_), .A2(new_n684_), .A3(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n678_), .ZN(new_n687_));
  OR3_X1    g486(.A1(new_n666_), .A2(G8gat), .A3(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n686_), .A2(KEYINPUT40), .A3(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(G1325gat));
  OAI21_X1  g492(.A(G15gat), .B1(new_n675_), .B2(new_n490_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n694_), .A2(KEYINPUT41), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(KEYINPUT41), .ZN(new_n696_));
  OR3_X1    g495(.A1(new_n666_), .A2(G15gat), .A3(new_n490_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n695_), .A2(new_n696_), .A3(new_n697_), .ZN(G1326gat));
  OR3_X1    g497(.A1(new_n666_), .A2(G22gat), .A3(new_n496_), .ZN(new_n699_));
  OAI21_X1  g498(.A(G22gat), .B1(new_n675_), .B2(new_n496_), .ZN(new_n700_));
  XOR2_X1   g499(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n701_));
  AND2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n700_), .A2(new_n701_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(G1327gat));
  INV_X1    g503(.A(new_n664_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n669_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n613_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n425_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G29gat), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT43), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n645_), .B1(new_n495_), .B2(new_n512_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n712_), .B1(new_n713_), .B2(KEYINPUT107), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT107), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n479_), .A2(new_n480_), .A3(KEYINPUT87), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n716_), .A2(new_n488_), .ZN(new_n717_));
  AOI221_X4 g516(.A(new_n717_), .B1(new_n501_), .B2(new_n510_), .C1(new_n459_), .C2(new_n491_), .ZN(new_n718_));
  AOI211_X1 g517(.A(new_n449_), .B(new_n457_), .C1(new_n446_), .C2(new_n447_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n448_), .A2(new_n458_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n481_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n459_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n718_), .B1(new_n723_), .B2(new_n427_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n715_), .B(KEYINPUT43), .C1(new_n724_), .C2(new_n645_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n714_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n612_), .A2(new_n664_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n726_), .A2(KEYINPUT44), .A3(new_n728_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n729_), .A2(G29gat), .A3(new_n710_), .ZN(new_n730_));
  NOR3_X1   g529(.A1(new_n713_), .A2(KEYINPUT107), .A3(new_n712_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n426_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n646_), .B1(new_n732_), .B2(new_n718_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT43), .B1(new_n733_), .B2(new_n715_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n728_), .B1(new_n731_), .B2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n711_), .B1(new_n730_), .B2(new_n737_), .ZN(G1328gat));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n739_), .B1(KEYINPUT110), .B2(KEYINPUT46), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(KEYINPUT110), .B2(KEYINPUT46), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n678_), .B(KEYINPUT108), .ZN(new_n742_));
  INV_X1    g541(.A(new_n742_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n708_), .A2(G36gat), .A3(new_n743_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT45), .Z(new_n745_));
  NAND2_X1  g544(.A1(new_n729_), .A2(new_n678_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT44), .B1(new_n726_), .B2(new_n728_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G36gat), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n741_), .B1(new_n745_), .B2(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n745_), .A2(new_n748_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT46), .B1(KEYINPUT109), .B2(KEYINPUT110), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n750_), .B2(new_n751_), .ZN(G1329gat));
  INV_X1    g551(.A(G43gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n753_), .B1(new_n708_), .B2(new_n490_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n755_));
  AOI211_X1 g554(.A(new_n736_), .B(new_n727_), .C1(new_n714_), .C2(new_n725_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n747_), .A2(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n493_), .A2(new_n753_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n755_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  AND4_X1   g558(.A1(new_n755_), .A2(new_n737_), .A3(new_n729_), .A4(new_n758_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n754_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  XOR2_X1   g560(.A(KEYINPUT112), .B(KEYINPUT47), .Z(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n762_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n754_), .B(new_n764_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1330gat));
  NOR3_X1   g565(.A1(new_n747_), .A2(new_n756_), .A3(new_n496_), .ZN(new_n767_));
  INV_X1    g566(.A(G50gat), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n496_), .A2(G50gat), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT113), .ZN(new_n770_));
  OAI22_X1  g569(.A1(new_n767_), .A2(new_n768_), .B1(new_n708_), .B2(new_n770_), .ZN(G1331gat));
  INV_X1    g570(.A(new_n574_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(new_n610_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n673_), .A2(new_n705_), .A3(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G57gat), .B1(new_n774_), .B2(new_n425_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n724_), .A2(new_n610_), .A3(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n665_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n710_), .A2(new_n352_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n775_), .B1(new_n777_), .B2(new_n778_), .ZN(G1332gat));
  OR3_X1    g578(.A1(new_n777_), .A2(G64gat), .A3(new_n743_), .ZN(new_n780_));
  OAI21_X1  g579(.A(G64gat), .B1(new_n774_), .B2(new_n743_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n781_), .A2(KEYINPUT48), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n781_), .A2(KEYINPUT48), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n780_), .B1(new_n782_), .B2(new_n783_), .ZN(G1333gat));
  OAI21_X1  g583(.A(G71gat), .B1(new_n774_), .B2(new_n490_), .ZN(new_n785_));
  XOR2_X1   g584(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n786_), .ZN(new_n788_));
  OAI211_X1 g587(.A(G71gat), .B(new_n788_), .C1(new_n774_), .C2(new_n490_), .ZN(new_n789_));
  OR3_X1    g588(.A1(new_n777_), .A2(G71gat), .A3(new_n490_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT115), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n787_), .A2(new_n793_), .A3(new_n789_), .A4(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1334gat));
  OAI21_X1  g594(.A(G78gat), .B1(new_n774_), .B2(new_n496_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n796_), .A2(KEYINPUT50), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(KEYINPUT50), .ZN(new_n798_));
  INV_X1    g597(.A(new_n496_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n517_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT116), .ZN(new_n801_));
  OAI22_X1  g600(.A1(new_n797_), .A2(new_n798_), .B1(new_n777_), .B2(new_n801_), .ZN(G1335gat));
  NAND2_X1  g601(.A1(new_n776_), .A2(new_n707_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n532_), .B1(new_n803_), .B2(new_n425_), .ZN(new_n804_));
  XOR2_X1   g603(.A(new_n804_), .B(KEYINPUT117), .Z(new_n805_));
  NAND3_X1  g604(.A1(new_n726_), .A2(new_n664_), .A3(new_n773_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n806_), .A2(new_n532_), .A3(new_n425_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1336gat));
  OAI21_X1  g607(.A(G92gat), .B1(new_n806_), .B2(new_n743_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n803_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n810_), .A2(new_n533_), .A3(new_n678_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(G1337gat));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(KEYINPUT51), .ZN(new_n814_));
  OAI21_X1  g613(.A(G99gat), .B1(new_n806_), .B2(new_n490_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n810_), .A2(new_n481_), .A3(new_n526_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n814_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n813_), .A2(KEYINPUT51), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n817_), .B(new_n818_), .Z(G1338gat));
  NAND3_X1  g618(.A1(new_n810_), .A2(new_n527_), .A3(new_n799_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n726_), .A2(new_n799_), .A3(new_n664_), .A4(new_n773_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n821_), .A2(new_n822_), .A3(G106gat), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n822_), .B1(new_n821_), .B2(G106gat), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n820_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n825_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g625(.A1(new_n494_), .A2(new_n710_), .A3(new_n687_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT121), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n562_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n558_), .A2(KEYINPUT12), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n554_), .B1(new_n832_), .B2(new_n552_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n561_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n515_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n543_), .A2(new_n547_), .A3(new_n525_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n658_), .A2(new_n560_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(new_n837_), .B2(new_n557_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n838_), .A2(KEYINPUT55), .A3(new_n514_), .A4(new_n561_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n831_), .A2(new_n835_), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT56), .B1(new_n840_), .B2(new_n568_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n840_), .A2(KEYINPUT56), .A3(new_n568_), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n610_), .B(new_n571_), .C1(new_n841_), .C2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n603_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n578_), .B1(new_n602_), .B2(new_n579_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n609_), .A2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n572_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n669_), .B1(new_n843_), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n829_), .B1(new_n849_), .B2(KEYINPUT57), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n607_), .A2(new_n577_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n851_), .A2(KEYINPUT79), .A3(new_n609_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n605_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n853_), .A3(new_n571_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n842_), .A2(new_n841_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n848_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n706_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT57), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(KEYINPUT119), .A3(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n850_), .A2(new_n859_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n847_), .A2(new_n571_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n840_), .A2(KEYINPUT56), .A3(new_n568_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT120), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n841_), .B2(new_n863_), .ZN(new_n864_));
  AOI211_X1 g663(.A(KEYINPUT120), .B(KEYINPUT56), .C1(new_n840_), .C2(new_n568_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n861_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(KEYINPUT58), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n861_), .B(new_n868_), .C1(new_n864_), .C2(new_n865_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n870_), .A2(new_n646_), .B1(new_n849_), .B2(KEYINPUT57), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n705_), .B1(new_n860_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n574_), .A2(new_n610_), .ZN(new_n874_));
  AND3_X1   g673(.A1(new_n665_), .A2(new_n873_), .A3(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n873_), .B1(new_n665_), .B2(new_n874_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n828_), .B1(new_n872_), .B2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT59), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n857_), .A2(new_n858_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n705_), .B1(new_n871_), .B2(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n880_), .B(new_n828_), .C1(new_n882_), .C2(new_n877_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n879_), .A2(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G113gat), .B1(new_n884_), .B2(new_n611_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n611_), .A2(G113gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n878_), .B2(new_n886_), .ZN(G1340gat));
  INV_X1    g686(.A(new_n828_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n870_), .A2(new_n646_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n849_), .A2(KEYINPUT57), .ZN(new_n890_));
  AOI21_X1  g689(.A(KEYINPUT119), .B1(new_n857_), .B2(new_n858_), .ZN(new_n891_));
  AOI211_X1 g690(.A(new_n829_), .B(KEYINPUT57), .C1(new_n856_), .C2(new_n706_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n889_), .B(new_n890_), .C1(new_n891_), .C2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n664_), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n875_), .A2(new_n876_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n888_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n883_), .B(new_n574_), .C1(new_n896_), .C2(new_n880_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(KEYINPUT122), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT122), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n879_), .A2(new_n899_), .A3(new_n574_), .A4(new_n883_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n898_), .A2(new_n900_), .A3(G120gat), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n772_), .A2(KEYINPUT60), .A3(G120gat), .ZN(new_n902_));
  AND2_X1   g701(.A1(KEYINPUT60), .A2(G120gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n896_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n904_), .ZN(G1341gat));
  OAI21_X1  g704(.A(G127gat), .B1(new_n884_), .B2(new_n664_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n664_), .A2(G127gat), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n878_), .B2(new_n907_), .ZN(G1342gat));
  OAI21_X1  g707(.A(G134gat), .B1(new_n884_), .B2(new_n645_), .ZN(new_n909_));
  OR2_X1    g708(.A1(new_n670_), .A2(G134gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n878_), .B2(new_n910_), .ZN(G1343gat));
  NOR2_X1   g710(.A1(new_n742_), .A2(new_n425_), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n492_), .B(new_n912_), .C1(new_n872_), .C2(new_n877_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n611_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n362_), .ZN(G1344gat));
  NOR2_X1   g714(.A1(new_n913_), .A2(new_n772_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(new_n363_), .ZN(G1345gat));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(new_n913_), .B2(new_n664_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n722_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n920_));
  NAND4_X1  g719(.A1(new_n920_), .A2(KEYINPUT123), .A3(new_n705_), .A4(new_n912_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT61), .B(G155gat), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n919_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n922_), .B1(new_n919_), .B2(new_n921_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(G1346gat));
  OAI21_X1  g724(.A(G162gat), .B1(new_n913_), .B2(new_n645_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n670_), .A2(G162gat), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n926_), .B1(new_n913_), .B2(new_n928_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n926_), .B(KEYINPUT124), .C1(new_n913_), .C2(new_n928_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1347gat));
  NOR2_X1   g732(.A1(new_n882_), .A2(new_n877_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n742_), .A2(new_n425_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n717_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n937_), .A2(new_n799_), .ZN(new_n938_));
  INV_X1    g737(.A(new_n938_), .ZN(new_n939_));
  NOR2_X1   g738(.A1(new_n934_), .A2(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(new_n610_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(G169gat), .ZN(new_n942_));
  XNOR2_X1  g741(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n942_), .A2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n943_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n941_), .A2(G169gat), .A3(new_n945_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n278_), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n944_), .B(new_n946_), .C1(new_n947_), .C2(new_n941_), .ZN(G1348gat));
  AOI21_X1  g747(.A(G176gat), .B1(new_n940_), .B2(new_n574_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n799_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n937_), .A2(new_n214_), .A3(new_n772_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n949_), .B1(new_n950_), .B2(new_n951_), .ZN(G1349gat));
  NOR2_X1   g751(.A1(new_n664_), .A2(new_n234_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n937_), .A2(new_n664_), .ZN(new_n954_));
  OAI211_X1 g753(.A(new_n496_), .B(new_n954_), .C1(new_n872_), .C2(new_n877_), .ZN(new_n955_));
  AOI22_X1  g754(.A1(new_n940_), .A2(new_n953_), .B1(new_n955_), .B2(new_n230_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(KEYINPUT126), .ZN(G1350gat));
  INV_X1    g756(.A(new_n235_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n670_), .A2(new_n958_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n940_), .A2(new_n959_), .ZN(new_n960_));
  NOR3_X1   g759(.A1(new_n934_), .A2(new_n645_), .A3(new_n939_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n960_), .B1(new_n961_), .B2(new_n297_), .ZN(G1351gat));
  OAI211_X1 g761(.A(new_n492_), .B(new_n936_), .C1(new_n872_), .C2(new_n877_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n963_), .A2(new_n611_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n964_), .B(new_n254_), .ZN(G1352gat));
  NOR2_X1   g764(.A1(new_n963_), .A2(new_n772_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n966_), .A2(new_n250_), .ZN(new_n967_));
  OAI21_X1  g766(.A(new_n967_), .B1(new_n248_), .B2(new_n966_), .ZN(G1353gat));
  NOR2_X1   g767(.A1(new_n963_), .A2(new_n664_), .ZN(new_n969_));
  INV_X1    g768(.A(KEYINPUT127), .ZN(new_n970_));
  XOR2_X1   g769(.A(KEYINPUT63), .B(G211gat), .Z(new_n971_));
  NAND3_X1  g770(.A1(new_n969_), .A2(new_n970_), .A3(new_n971_), .ZN(new_n972_));
  OR2_X1    g771(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n972_), .B1(new_n969_), .B2(new_n973_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n970_), .B1(new_n969_), .B2(new_n971_), .ZN(new_n975_));
  NOR2_X1   g774(.A1(new_n974_), .A2(new_n975_), .ZN(G1354gat));
  OAI21_X1  g775(.A(G218gat), .B1(new_n963_), .B2(new_n645_), .ZN(new_n977_));
  OR2_X1    g776(.A1(new_n670_), .A2(G218gat), .ZN(new_n978_));
  OAI21_X1  g777(.A(new_n977_), .B1(new_n963_), .B2(new_n978_), .ZN(G1355gat));
endmodule


