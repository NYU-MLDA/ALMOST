//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n925_, new_n926_, new_n927_, new_n929_, new_n930_, new_n931_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202_));
  NOR2_X1   g001(.A1(G141gat), .A2(G148gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G141gat), .A2(G148gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n207_), .B1(new_n209_), .B2(KEYINPUT1), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n206_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n207_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n212_), .A2(new_n209_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT3), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n203_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT2), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n205_), .A2(KEYINPUT86), .A3(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n215_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n216_), .B1(new_n205_), .B2(KEYINPUT86), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n213_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT87), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OAI211_X1 g022(.A(KEYINPUT87), .B(new_n213_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n211_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT29), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G197gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT89), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT89), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G197gat), .ZN(new_n231_));
  INV_X1    g030(.A(G204gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n229_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT21), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n234_), .B1(G197gat), .B2(G204gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT90), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT90), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n233_), .A2(new_n238_), .A3(new_n235_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G211gat), .B(G218gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n228_), .A2(new_n232_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT89), .B(G197gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(new_n232_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n242_), .B1(new_n245_), .B2(new_n234_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n240_), .A2(new_n246_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n245_), .A2(new_n234_), .A3(new_n241_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT92), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n248_), .B1(new_n240_), .B2(new_n246_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT92), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n227_), .B1(new_n251_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G233gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT88), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n257_), .A2(G228gat), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(G228gat), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n256_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT93), .B1(new_n255_), .B2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G78gat), .B(G106gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT91), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n250_), .A2(new_n262_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n266_), .B1(new_n267_), .B2(new_n227_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n252_), .A2(new_n261_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n269_), .B(KEYINPUT91), .C1(new_n226_), .C2(new_n225_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT93), .ZN(new_n272_));
  AOI211_X1 g071(.A(KEYINPUT92), .B(new_n248_), .C1(new_n240_), .C2(new_n246_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n253_), .B1(new_n247_), .B2(new_n249_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n272_), .B(new_n261_), .C1(new_n275_), .C2(new_n227_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n263_), .A2(new_n265_), .A3(new_n271_), .A4(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT94), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n225_), .A2(new_n226_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G22gat), .B(G50gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT28), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n279_), .B(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n202_), .B1(new_n278_), .B2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n282_), .ZN(new_n284_));
  AOI211_X1 g083(.A(KEYINPUT95), .B(new_n284_), .C1(new_n277_), .C2(KEYINPUT94), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n263_), .A2(new_n271_), .A3(new_n276_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(new_n264_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n277_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n283_), .A2(new_n285_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT23), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n294_));
  INV_X1    g093(.A(G183gat), .ZN(new_n295_));
  INV_X1    g094(.A(G190gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n294_), .A3(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n298_), .A2(KEYINPUT83), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G169gat), .A2(G176gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(KEYINPUT83), .ZN(new_n301_));
  INV_X1    g100(.A(G176gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT22), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT82), .B1(new_n303_), .B2(G169gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT22), .B(G169gat), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n302_), .B(new_n304_), .C1(new_n305_), .C2(KEYINPUT82), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .A4(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT81), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT81), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n310_), .B1(G169gat), .B2(G176gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n309_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT24), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n309_), .A2(KEYINPUT24), .A3(new_n311_), .A4(new_n300_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n293_), .A2(new_n294_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT25), .B(G183gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT26), .B(G190gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n314_), .A2(new_n315_), .A3(new_n317_), .A4(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n307_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT30), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT84), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G71gat), .B(G99gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(G43gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G227gat), .A2(G233gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n329_), .B(G15gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n328_), .B(new_n330_), .ZN(new_n331_));
  OR2_X1    g130(.A1(new_n326_), .A2(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(new_n324_), .A2(new_n325_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n326_), .A2(new_n331_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G127gat), .B(G134gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G113gat), .B(G120gat), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n336_), .A2(new_n337_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT31), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n335_), .A2(KEYINPUT85), .A3(new_n342_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n335_), .A2(KEYINPUT85), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n341_), .B1(new_n335_), .B2(KEYINPUT85), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n343_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G1gat), .B(G29gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(G85gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT0), .B(G57gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  NAND2_X1  g149(.A1(G225gat), .A2(G233gat), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n223_), .A2(new_n224_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n340_), .B1(new_n352_), .B2(new_n211_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n340_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n225_), .A2(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n353_), .A2(KEYINPUT4), .A3(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n225_), .A2(new_n354_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n351_), .B1(new_n356_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n351_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n350_), .B1(new_n360_), .B2(new_n362_), .ZN(new_n363_));
  AOI211_X1 g162(.A(new_n211_), .B(new_n340_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n364_));
  NOR3_X1   g163(.A1(new_n357_), .A2(new_n364_), .A3(new_n358_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n353_), .A2(KEYINPUT4), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n361_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n350_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n362_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n368_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n363_), .A2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n346_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G226gat), .A2(G233gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT19), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT20), .B1(new_n250_), .B2(new_n322_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(KEYINPUT26), .B(G190gat), .Z(new_n377_));
  INV_X1    g176(.A(KEYINPUT96), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n319_), .A2(KEYINPUT96), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n318_), .A3(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n315_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT97), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n381_), .A2(KEYINPUT97), .A3(new_n315_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT98), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n386_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT24), .B1(new_n309_), .B2(new_n311_), .ZN(new_n388_));
  NOR3_X1   g187(.A1(new_n388_), .A2(new_n316_), .A3(KEYINPUT98), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n387_), .A2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n384_), .A2(new_n385_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n305_), .A2(new_n302_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n300_), .ZN(new_n393_));
  OR2_X1    g192(.A1(new_n393_), .A2(KEYINPUT99), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(KEYINPUT99), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n298_), .A3(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n374_), .B(new_n376_), .C1(new_n397_), .C2(new_n252_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n391_), .A2(new_n252_), .A3(new_n396_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT20), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n400_), .B1(new_n250_), .B2(new_n322_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n374_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G8gat), .B(G36gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT18), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(new_n406_), .B(new_n407_), .Z(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n398_), .A2(new_n404_), .A3(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n252_), .B1(new_n391_), .B2(new_n396_), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n411_), .A2(new_n403_), .A3(new_n375_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n374_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n408_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n410_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT27), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT104), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT104), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n415_), .A2(new_n419_), .A3(new_n416_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n252_), .B1(new_n307_), .B2(new_n321_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n400_), .B1(new_n397_), .B2(new_n275_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT103), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n421_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n251_), .A2(new_n254_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n391_), .A2(new_n396_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT20), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT103), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n403_), .B1(new_n424_), .B2(new_n428_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(new_n411_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n409_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n398_), .A2(new_n404_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n416_), .B1(new_n432_), .B2(new_n408_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n418_), .A2(new_n420_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n288_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n435_));
  AND4_X1   g234(.A1(new_n290_), .A2(new_n372_), .A3(new_n434_), .A4(new_n435_), .ZN(new_n436_));
  NOR3_X1   g235(.A1(new_n357_), .A2(new_n364_), .A3(new_n351_), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT101), .B1(new_n437_), .B2(new_n350_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n356_), .A2(new_n351_), .A3(new_n359_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n353_), .A2(new_n361_), .A3(new_n355_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT101), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(new_n441_), .A3(new_n368_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n439_), .A3(new_n442_), .ZN(new_n443_));
  AND3_X1   g242(.A1(new_n414_), .A2(new_n410_), .A3(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n368_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT33), .B1(new_n445_), .B2(KEYINPUT100), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT100), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT33), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n363_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n444_), .A2(new_n446_), .A3(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT102), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n408_), .A2(KEYINPUT32), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n363_), .A2(new_n370_), .B1(new_n432_), .B2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n429_), .A2(new_n430_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n454_), .B1(new_n455_), .B2(new_n453_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n444_), .A2(new_n446_), .A3(KEYINPUT102), .A4(new_n449_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n452_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(new_n290_), .A3(new_n435_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n371_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n278_), .A2(new_n282_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT95), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n278_), .A2(new_n202_), .A3(new_n282_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n462_), .A2(new_n463_), .B1(new_n277_), .B2(new_n287_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n434_), .B(new_n460_), .C1(new_n464_), .C2(new_n289_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n459_), .A2(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n436_), .B1(new_n466_), .B2(new_n346_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT79), .ZN(new_n468_));
  XOR2_X1   g267(.A(G29gat), .B(G36gat), .Z(new_n469_));
  XOR2_X1   g268(.A(G43gat), .B(G50gat), .Z(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT74), .B(G15gat), .ZN(new_n473_));
  INV_X1    g272(.A(G22gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G1gat), .ZN(new_n476_));
  INV_X1    g275(.A(G8gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT14), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G1gat), .B(G8gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n479_), .A2(new_n480_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n472_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n479_), .A2(new_n480_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n481_), .A3(new_n471_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G229gat), .A2(G233gat), .ZN(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n471_), .B(KEYINPUT15), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n491_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n492_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G113gat), .B(G141gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G169gat), .B(G197gat), .ZN(new_n495_));
  XOR2_X1   g294(.A(new_n494_), .B(new_n495_), .Z(new_n496_));
  AND3_X1   g295(.A1(new_n490_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n490_), .B2(new_n493_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n468_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n490_), .A2(new_n493_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n496_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n490_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(KEYINPUT79), .A3(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n500_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT80), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n467_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G71gat), .B(G78gat), .ZN(new_n511_));
  INV_X1    g310(.A(G64gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(G57gat), .ZN(new_n513_));
  INV_X1    g312(.A(G57gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(G64gat), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n511_), .A2(KEYINPUT11), .A3(new_n513_), .A4(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n513_), .A2(new_n515_), .A3(KEYINPUT11), .ZN(new_n517_));
  INV_X1    g316(.A(G78gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(G71gat), .ZN(new_n519_));
  INV_X1    g318(.A(G71gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(G78gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n517_), .A2(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT11), .B1(new_n513_), .B2(new_n515_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n516_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  OAI211_X1 g325(.A(G231gat), .B(G233gat), .C1(new_n482_), .C2(new_n483_), .ZN(new_n527_));
  INV_X1    g326(.A(G231gat), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n485_), .B(new_n481_), .C1(new_n528_), .C2(new_n256_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n526_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n527_), .A2(new_n529_), .A3(new_n526_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n531_), .A2(KEYINPUT66), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT66), .ZN(new_n534_));
  INV_X1    g333(.A(new_n532_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n534_), .B1(new_n535_), .B2(new_n530_), .ZN(new_n536_));
  XOR2_X1   g335(.A(G127gat), .B(G155gat), .Z(new_n537_));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT17), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n542_), .B(KEYINPUT76), .Z(new_n543_));
  NAND3_X1  g342(.A1(new_n533_), .A2(new_n536_), .A3(new_n543_), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n541_), .A2(KEYINPUT17), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n531_), .A2(new_n532_), .A3(new_n542_), .A4(new_n545_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n544_), .A2(KEYINPUT77), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT77), .B1(new_n544_), .B2(new_n546_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT78), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n544_), .A2(new_n546_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT77), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT78), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n544_), .A2(KEYINPUT77), .A3(new_n546_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n549_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n556_), .ZN(new_n557_));
  XOR2_X1   g356(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT68), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G120gat), .B(G148gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G176gat), .B(G204gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n561_), .B(new_n562_), .Z(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT65), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT7), .ZN(new_n566_));
  NOR2_X1   g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n566_), .B1(new_n567_), .B2(KEYINPUT64), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT64), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n569_), .A2(G99gat), .A3(G106gat), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n565_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n567_), .A2(KEYINPUT64), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n569_), .B1(G99gat), .B2(G106gat), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n572_), .A2(new_n573_), .A3(KEYINPUT65), .A4(new_n566_), .ZN(new_n574_));
  INV_X1    g373(.A(G99gat), .ZN(new_n575_));
  INV_X1    g374(.A(G106gat), .ZN(new_n576_));
  OAI21_X1  g375(.A(KEYINPUT6), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT6), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(G99gat), .A3(G106gat), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n576_), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n577_), .A2(new_n579_), .B1(new_n580_), .B2(KEYINPUT7), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n571_), .A2(new_n574_), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(G85gat), .ZN(new_n583_));
  INV_X1    g382(.A(G92gat), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G85gat), .A2(G92gat), .ZN(new_n586_));
  AND2_X1   g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AND3_X1   g386(.A1(new_n582_), .A2(KEYINPUT8), .A3(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT8), .B1(new_n582_), .B2(new_n587_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n577_), .A2(new_n579_), .ZN(new_n590_));
  OR2_X1    g389(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n591_));
  NAND2_X1  g390(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n576_), .A3(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n585_), .A2(KEYINPUT9), .A3(new_n586_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n586_), .A2(KEYINPUT9), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n590_), .A2(new_n593_), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR4_X1   g396(.A1(new_n588_), .A2(new_n589_), .A3(new_n526_), .A4(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n525_), .A2(KEYINPUT66), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n516_), .B(new_n534_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(KEYINPUT12), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n582_), .A2(new_n587_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT8), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n597_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n582_), .A2(KEYINPUT8), .A3(new_n587_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n601_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n598_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n603_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(new_n605_), .A3(new_n596_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n526_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT12), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G230gat), .A2(G233gat), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n607_), .A2(new_n612_), .A3(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n604_), .A2(new_n525_), .A3(new_n605_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n610_), .A2(new_n615_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n564_), .B(new_n614_), .C1(new_n613_), .C2(new_n616_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n588_), .A2(new_n589_), .A3(new_n597_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n615_), .B1(new_n618_), .B2(new_n601_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT12), .B1(new_n609_), .B2(new_n526_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n613_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n619_), .A2(new_n620_), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n613_), .B1(new_n610_), .B2(new_n615_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n563_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n617_), .A2(new_n624_), .A3(KEYINPUT69), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT69), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n626_), .B(new_n563_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT13), .ZN(new_n629_));
  XOR2_X1   g428(.A(G190gat), .B(G218gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT70), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT36), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT72), .Z(new_n635_));
  NAND2_X1  g434(.A1(new_n618_), .A2(new_n471_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n609_), .A2(new_n491_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT71), .ZN(new_n638_));
  NAND2_X1  g437(.A1(G232gat), .A2(G233gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT34), .ZN(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT35), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n638_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n636_), .A2(new_n637_), .A3(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n641_), .A2(new_n642_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n645_), .ZN(new_n647_));
  NAND4_X1  g446(.A1(new_n636_), .A2(new_n637_), .A3(new_n647_), .A4(new_n643_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n635_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT36), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n646_), .A2(new_n651_), .A3(new_n648_), .A4(new_n633_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n650_), .A2(KEYINPUT37), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT73), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n650_), .A2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n635_), .A2(KEYINPUT73), .A3(new_n649_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(new_n652_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT37), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n654_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n557_), .A2(new_n629_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n510_), .A2(new_n662_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n663_), .A2(G1gat), .A3(new_n460_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT38), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(KEYINPUT38), .ZN(new_n666_));
  INV_X1    g465(.A(new_n658_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n467_), .A2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n547_), .A2(new_n548_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n507_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n629_), .A2(new_n670_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n668_), .A2(new_n669_), .A3(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G1gat), .B1(new_n672_), .B2(new_n460_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n665_), .A2(new_n666_), .A3(new_n673_), .ZN(G1324gat));
  OAI21_X1  g473(.A(G8gat), .B1(new_n672_), .B2(new_n434_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT39), .ZN(new_n676_));
  INV_X1    g475(.A(new_n663_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n434_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n477_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n676_), .A2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n680_), .B(new_n681_), .ZN(G1325gat));
  OAI21_X1  g481(.A(G15gat), .B1(new_n672_), .B2(new_n346_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT106), .B(KEYINPUT41), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n684_), .ZN(new_n686_));
  OR3_X1    g485(.A1(new_n663_), .A2(G15gat), .A3(new_n346_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n685_), .A2(new_n686_), .A3(new_n687_), .ZN(G1326gat));
  NOR2_X1   g487(.A1(new_n464_), .A2(new_n289_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G22gat), .B1(new_n672_), .B2(new_n689_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT42), .ZN(new_n691_));
  INV_X1    g490(.A(new_n689_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n677_), .A2(new_n474_), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1327gat));
  NOR3_X1   g493(.A1(new_n556_), .A2(new_n629_), .A3(new_n658_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n510_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(G29gat), .B1(new_n697_), .B2(new_n371_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n699_), .A2(KEYINPUT107), .ZN(new_n700_));
  INV_X1    g499(.A(new_n346_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n701_), .B1(new_n459_), .B2(new_n465_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n661_), .B(new_n700_), .C1(new_n702_), .C2(new_n436_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(new_n557_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n705_), .B1(new_n467_), .B2(new_n660_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n704_), .A2(new_n671_), .A3(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n704_), .A2(KEYINPUT44), .A3(new_n671_), .A4(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n371_), .A2(G29gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n698_), .B1(new_n712_), .B2(new_n713_), .ZN(G1328gat));
  OAI21_X1  g513(.A(G36gat), .B1(new_n711_), .B2(new_n434_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n696_), .A2(G36gat), .A3(new_n434_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT45), .Z(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n715_), .A2(new_n717_), .A3(KEYINPUT46), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1329gat));
  NAND2_X1  g521(.A1(new_n701_), .A2(G43gat), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n696_), .A2(new_n346_), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n711_), .A2(new_n723_), .B1(G43gat), .B2(new_n724_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g525(.A(G50gat), .B1(new_n697_), .B2(new_n692_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n692_), .A2(G50gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n712_), .B2(new_n728_), .ZN(G1331gat));
  NAND4_X1  g528(.A1(new_n668_), .A2(new_n509_), .A3(new_n629_), .A4(new_n556_), .ZN(new_n730_));
  OAI21_X1  g529(.A(G57gat), .B1(new_n730_), .B2(new_n460_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n629_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n467_), .A2(new_n507_), .A3(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n556_), .A3(new_n660_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n371_), .A2(new_n514_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(G1332gat));
  OAI21_X1  g535(.A(G64gat), .B1(new_n730_), .B2(new_n434_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT48), .ZN(new_n738_));
  INV_X1    g537(.A(new_n734_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(new_n512_), .A3(new_n678_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT108), .Z(G1333gat));
  OAI21_X1  g541(.A(G71gat), .B1(new_n730_), .B2(new_n346_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT49), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n739_), .A2(new_n520_), .A3(new_n701_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1334gat));
  OAI21_X1  g545(.A(G78gat), .B1(new_n730_), .B2(new_n689_), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n747_), .B(KEYINPUT50), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n739_), .A2(new_n518_), .A3(new_n692_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1335gat));
  NOR2_X1   g549(.A1(new_n556_), .A2(new_n658_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n733_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n583_), .A3(new_n371_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n732_), .A2(new_n507_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n706_), .A2(new_n557_), .A3(new_n703_), .A4(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND4_X1  g557(.A1(new_n704_), .A2(KEYINPUT109), .A3(new_n706_), .A4(new_n755_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(KEYINPUT110), .ZN(new_n760_));
  AOI21_X1  g559(.A(KEYINPUT110), .B1(new_n758_), .B2(new_n759_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n460_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n754_), .B1(new_n762_), .B2(new_n583_), .ZN(G1336gat));
  NAND3_X1  g562(.A1(new_n753_), .A2(new_n584_), .A3(new_n678_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n760_), .A2(new_n761_), .A3(new_n434_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n765_), .B2(new_n584_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT111), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n768_), .B(new_n764_), .C1(new_n765_), .C2(new_n584_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1337gat));
  AND4_X1   g569(.A1(new_n701_), .A2(new_n753_), .A3(new_n591_), .A4(new_n592_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n758_), .A2(new_n759_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(new_n701_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n771_), .B1(new_n773_), .B2(G99gat), .ZN(new_n774_));
  XOR2_X1   g573(.A(new_n774_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g574(.A1(new_n753_), .A2(new_n576_), .A3(new_n692_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n756_), .A2(new_n689_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n576_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT112), .B1(new_n756_), .B2(new_n689_), .ZN(new_n780_));
  XOR2_X1   g579(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n781_));
  AND3_X1   g580(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n776_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n776_), .B(new_n785_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1339gat));
  NAND4_X1  g588(.A1(new_n556_), .A2(new_n732_), .A3(new_n509_), .A4(new_n660_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT54), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n499_), .A2(new_n505_), .A3(new_n617_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n613_), .B1(new_n607_), .B2(new_n612_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n614_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  NOR4_X1   g594(.A1(new_n619_), .A2(new_n620_), .A3(new_n794_), .A4(new_n621_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n563_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  AOI211_X1 g599(.A(new_n800_), .B(new_n564_), .C1(new_n795_), .C2(new_n797_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n792_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n492_), .A2(new_n486_), .A3(new_n489_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n496_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n497_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n625_), .A2(new_n805_), .A3(KEYINPUT115), .A4(new_n627_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n625_), .A2(new_n805_), .A3(new_n627_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT115), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n802_), .A2(new_n806_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n810_), .A2(new_n811_), .A3(new_n658_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n810_), .B2(new_n658_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n805_), .A2(new_n617_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n799_), .B2(KEYINPUT116), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n621_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n622_), .B1(KEYINPUT55), .B2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n563_), .B1(new_n818_), .B2(new_n796_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n800_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n563_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n816_), .A2(new_n823_), .A3(KEYINPUT58), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n816_), .A2(new_n823_), .A3(KEYINPUT118), .A4(KEYINPUT58), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT58), .B1(new_n816_), .B2(new_n823_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT117), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n660_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n828_), .A2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n830_), .B1(new_n829_), .B2(new_n660_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n814_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT119), .B(new_n791_), .C1(new_n834_), .C2(new_n669_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n816_), .A2(new_n823_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT58), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(KEYINPUT117), .A3(new_n661_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n840_), .A2(new_n833_), .A3(new_n827_), .A4(new_n826_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n813_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n810_), .A2(new_n811_), .A3(new_n658_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n669_), .B1(new_n841_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n790_), .B(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n836_), .B1(new_n845_), .B2(new_n847_), .ZN(new_n848_));
  NOR4_X1   g647(.A1(new_n692_), .A2(new_n460_), .A3(new_n678_), .A4(new_n346_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n835_), .A2(new_n848_), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(G113gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n507_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n509_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n791_), .B1(new_n834_), .B2(new_n556_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n856_));
  AND2_X1   g655(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n855_), .B(new_n849_), .C1(new_n856_), .C2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859_));
  AND3_X1   g658(.A1(new_n850_), .A2(new_n859_), .A3(KEYINPUT59), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n850_), .B2(KEYINPUT59), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n854_), .B(new_n858_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n853_), .B1(new_n863_), .B2(new_n852_), .ZN(G1340gat));
  INV_X1    g663(.A(G120gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n732_), .B2(KEYINPUT60), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n851_), .B(new_n866_), .C1(KEYINPUT60), .C2(new_n865_), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n629_), .B(new_n858_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n867_), .B1(new_n869_), .B2(new_n865_), .ZN(G1341gat));
  INV_X1    g669(.A(G127gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n851_), .A2(new_n871_), .A3(new_n556_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n669_), .B(new_n858_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n872_), .B1(new_n874_), .B2(new_n871_), .ZN(G1342gat));
  INV_X1    g674(.A(G134gat), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n660_), .A2(new_n876_), .ZN(new_n877_));
  OAI211_X1 g676(.A(new_n858_), .B(new_n877_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n876_), .B1(new_n850_), .B2(new_n658_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n878_), .A2(KEYINPUT122), .A3(new_n879_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(G1343gat));
  AND3_X1   g683(.A1(new_n835_), .A2(new_n848_), .A3(new_n346_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n689_), .A2(new_n678_), .A3(new_n460_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n507_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n887_), .A2(new_n890_), .A3(new_n629_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n885_), .A2(new_n886_), .ZN(new_n892_));
  OAI21_X1  g691(.A(KEYINPUT124), .B1(new_n892_), .B2(new_n732_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT123), .B(G148gat), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n891_), .A2(new_n893_), .A3(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1345gat));
  NAND2_X1  g696(.A1(new_n887_), .A2(new_n556_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(KEYINPUT61), .B(G155gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1346gat));
  OR3_X1    g699(.A1(new_n892_), .A2(G162gat), .A3(new_n658_), .ZN(new_n901_));
  OAI21_X1  g700(.A(G162gat), .B1(new_n892_), .B2(new_n660_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1347gat));
  NAND2_X1  g702(.A1(new_n678_), .A2(new_n372_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n692_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n855_), .A2(new_n905_), .ZN(new_n906_));
  OAI21_X1  g705(.A(G169gat), .B1(new_n906_), .B2(new_n670_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n907_), .A2(KEYINPUT62), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(KEYINPUT62), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n507_), .A2(new_n305_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT125), .ZN(new_n911_));
  OAI22_X1  g710(.A1(new_n908_), .A2(new_n909_), .B1(new_n906_), .B2(new_n911_), .ZN(G1348gat));
  AND2_X1   g711(.A1(new_n835_), .A2(new_n848_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n904_), .A2(new_n732_), .A3(new_n302_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n913_), .A2(new_n689_), .A3(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n302_), .B1(new_n906_), .B2(new_n732_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n917_), .B(KEYINPUT126), .Z(G1349gat));
  NOR2_X1   g717(.A1(new_n557_), .A2(new_n904_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n913_), .A2(new_n689_), .A3(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n906_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n669_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n318_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n920_), .A2(new_n295_), .B1(new_n921_), .B2(new_n923_), .ZN(G1350gat));
  NAND4_X1  g723(.A1(new_n921_), .A2(new_n379_), .A3(new_n380_), .A4(new_n667_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n921_), .A2(new_n661_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n925_), .B1(new_n927_), .B2(new_n296_), .ZN(G1351gat));
  NOR3_X1   g727(.A1(new_n689_), .A2(new_n371_), .A3(new_n434_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n885_), .A2(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(new_n670_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(new_n228_), .ZN(G1352gat));
  NOR2_X1   g731(.A1(new_n930_), .A2(new_n732_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(new_n232_), .ZN(G1353gat));
  INV_X1    g733(.A(KEYINPUT63), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n922_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(KEYINPUT127), .B1(new_n930_), .B2(new_n937_), .ZN(new_n938_));
  INV_X1    g737(.A(G211gat), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n940_));
  NAND4_X1  g739(.A1(new_n885_), .A2(new_n940_), .A3(new_n929_), .A4(new_n936_), .ZN(new_n941_));
  AND4_X1   g740(.A1(new_n935_), .A2(new_n938_), .A3(new_n939_), .A4(new_n941_), .ZN(new_n942_));
  AOI22_X1  g741(.A1(new_n938_), .A2(new_n941_), .B1(new_n935_), .B2(new_n939_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n942_), .A2(new_n943_), .ZN(G1354gat));
  OAI21_X1  g743(.A(G218gat), .B1(new_n930_), .B2(new_n660_), .ZN(new_n945_));
  OR2_X1    g744(.A1(new_n658_), .A2(G218gat), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n930_), .B2(new_n946_), .ZN(G1355gat));
endmodule


