//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n857_, new_n858_,
    new_n859_, new_n860_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT82), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G141gat), .A2(G148gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT81), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT80), .ZN(new_n215_));
  AOI22_X1  g014(.A1(new_n211_), .A2(new_n213_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT81), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT82), .B1(new_n217_), .B2(KEYINPUT2), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(new_n212_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT3), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n220_), .A2(new_n221_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n220_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(KEYINPUT80), .A3(KEYINPUT3), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n216_), .A2(new_n219_), .A3(new_n222_), .A4(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT83), .ZN(new_n226_));
  NOR2_X1   g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n226_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n229_), .ZN(new_n231_));
  NOR3_X1   g030(.A1(new_n231_), .A2(new_n227_), .A3(KEYINPUT83), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n225_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n223_), .A2(new_n212_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT1), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n227_), .B1(new_n231_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n229_), .A2(KEYINPUT1), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n235_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n234_), .A2(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G127gat), .B(G134gat), .Z(new_n242_));
  XOR2_X1   g041(.A(G113gat), .B(G120gat), .Z(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n241_), .A2(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n239_), .B1(new_n225_), .B2(new_n233_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n244_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(KEYINPUT94), .A3(new_n248_), .ZN(new_n249_));
  OR3_X1    g048(.A1(new_n247_), .A2(KEYINPUT94), .A3(new_n244_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n208_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(KEYINPUT95), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(KEYINPUT95), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n249_), .A2(new_n250_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT4), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n246_), .A2(KEYINPUT4), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n256_), .A2(new_n208_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n206_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n258_), .A2(new_n252_), .A3(new_n205_), .A4(new_n253_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G169gat), .ZN(new_n263_));
  INV_X1    g062(.A(G176gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  MUX2_X1   g066(.A(new_n265_), .B(new_n267_), .S(KEYINPUT24), .Z(new_n268_));
  INV_X1    g067(.A(G190gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT26), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT26), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(G190gat), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G183gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT25), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT75), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT25), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(G183gat), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n275_), .A2(new_n278_), .ZN(new_n279_));
  OAI211_X1 g078(.A(new_n273_), .B(new_n276_), .C1(new_n279_), .C2(KEYINPUT75), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n283_));
  NAND2_X1  g082(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n281_), .A2(KEYINPUT23), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n268_), .B(new_n280_), .C1(new_n285_), .C2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G183gat), .A2(G190gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n283_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n290_), .A2(KEYINPUT79), .B1(KEYINPUT23), .B2(new_n281_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT79), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n283_), .A2(new_n282_), .A3(new_n292_), .A4(new_n284_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n289_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT78), .B(G169gat), .ZN(new_n295_));
  AOI21_X1  g094(.A(G176gat), .B1(KEYINPUT77), .B2(KEYINPUT22), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n288_), .B1(new_n294_), .B2(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G71gat), .B(G99gat), .ZN(new_n300_));
  INV_X1    g099(.A(G43gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n299_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(new_n244_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G227gat), .A2(G233gat), .ZN(new_n305_));
  INV_X1    g104(.A(G15gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT30), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT31), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n304_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n304_), .A2(new_n309_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n262_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT101), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT100), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT98), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT89), .B(KEYINPUT19), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G226gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  XOR2_X1   g119(.A(G211gat), .B(G218gat), .Z(new_n321_));
  INV_X1    g120(.A(G204gat), .ZN(new_n322_));
  OR3_X1    g121(.A1(new_n322_), .A2(KEYINPUT86), .A3(G197gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT86), .B1(new_n322_), .B2(G197gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT85), .B(G197gat), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n323_), .B(new_n324_), .C1(new_n325_), .C2(G204gat), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n321_), .B1(new_n326_), .B2(KEYINPUT21), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT21), .ZN(new_n328_));
  INV_X1    g127(.A(G197gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT85), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT85), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(G197gat), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n322_), .B1(new_n330_), .B2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(G197gat), .A2(G204gat), .ZN(new_n334_));
  OAI211_X1 g133(.A(KEYINPUT87), .B(new_n328_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n334_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n337_), .B1(new_n325_), .B2(new_n322_), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT87), .B1(new_n338_), .B2(new_n328_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n327_), .B1(new_n336_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n330_), .A2(new_n332_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n334_), .B1(new_n341_), .B2(G204gat), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n342_), .A2(KEYINPUT21), .A3(new_n321_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n340_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n290_), .A2(KEYINPUT79), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n281_), .A2(KEYINPUT23), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n293_), .A3(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(KEYINPUT90), .A2(KEYINPUT24), .ZN(new_n348_));
  NOR2_X1   g147(.A1(KEYINPUT90), .A2(KEYINPUT24), .ZN(new_n349_));
  OR2_X1    g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(new_n265_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n275_), .A2(new_n278_), .A3(new_n270_), .A4(new_n272_), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n265_), .B(new_n266_), .C1(new_n348_), .C2(new_n349_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT91), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n355_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n347_), .B(new_n352_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n359_));
  NOR2_X1   g158(.A1(KEYINPUT76), .A2(KEYINPUT23), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n281_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n289_), .B1(new_n361_), .B2(new_n286_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT92), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT22), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n365_), .A2(G169gat), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n263_), .A2(KEYINPUT22), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n364_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n263_), .A2(KEYINPUT22), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n365_), .A2(G169gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n369_), .A2(new_n370_), .A3(KEYINPUT92), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n363_), .B(new_n266_), .C1(new_n372_), .C2(G176gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n358_), .A2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT20), .B1(new_n344_), .B2(new_n374_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n294_), .A2(new_n298_), .ZN(new_n376_));
  AOI22_X1  g175(.A1(new_n376_), .A2(new_n288_), .B1(new_n340_), .B2(new_n343_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n320_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT20), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(new_n344_), .B2(new_n374_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n343_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT87), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n342_), .B2(KEYINPUT21), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(new_n335_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n381_), .B1(new_n384_), .B2(new_n327_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(new_n376_), .A3(new_n288_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n380_), .A2(new_n319_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n378_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT18), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G64gat), .B(G92gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n316_), .B1(new_n388_), .B2(new_n393_), .ZN(new_n394_));
  AOI211_X1 g193(.A(KEYINPUT98), .B(new_n392_), .C1(new_n378_), .C2(new_n387_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT27), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(G176gat), .B1(new_n368_), .B2(new_n371_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n266_), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n397_), .A2(new_n398_), .A3(new_n362_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n353_), .A2(new_n354_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n400_), .A2(KEYINPUT91), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n353_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n351_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n399_), .B1(new_n403_), .B2(new_n347_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT20), .B1(new_n404_), .B2(new_n385_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n344_), .A2(new_n299_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n320_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n379_), .B1(new_n404_), .B2(new_n385_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n344_), .A2(new_n299_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n319_), .A3(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n407_), .A2(new_n392_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT99), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n407_), .A2(new_n410_), .A3(KEYINPUT99), .A4(new_n392_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n315_), .B1(new_n396_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n388_), .A2(new_n393_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n417_), .A2(KEYINPUT98), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n388_), .A2(new_n316_), .A3(new_n393_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n413_), .A2(new_n414_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n420_), .A2(KEYINPUT100), .A3(KEYINPUT27), .A4(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n416_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT29), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n247_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n385_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n426_), .B1(new_n385_), .B2(new_n425_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n247_), .A2(new_n424_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G22gat), .B(G50gat), .Z(new_n431_));
  NOR2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n430_), .A2(new_n431_), .ZN(new_n433_));
  OAI22_X1  g232(.A1(new_n427_), .A2(new_n429_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n427_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n433_), .A2(new_n432_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n436_), .A3(new_n428_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n434_), .A2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G228gat), .A2(G233gat), .ZN(new_n439_));
  INV_X1    g238(.A(G78gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n434_), .A2(new_n437_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT88), .B(G106gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n442_), .A2(new_n446_), .A3(new_n444_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n407_), .A2(new_n410_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n393_), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT27), .B1(new_n452_), .B2(new_n411_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AND4_X1   g253(.A1(new_n314_), .A2(new_n423_), .A3(new_n450_), .A4(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n453_), .B1(new_n416_), .B2(new_n422_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n314_), .B1(new_n456_), .B2(new_n450_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n313_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n262_), .B1(new_n449_), .B2(new_n448_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n423_), .A2(new_n459_), .A3(new_n454_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n448_), .A2(new_n449_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n256_), .A2(new_n207_), .A3(new_n257_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n255_), .B(KEYINPUT97), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n205_), .B1(new_n463_), .B2(new_n208_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n452_), .A2(new_n411_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT93), .ZN(new_n466_));
  AOI22_X1  g265(.A1(new_n462_), .A2(new_n464_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n452_), .A2(KEYINPUT93), .A3(new_n411_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n254_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT96), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n470_), .A2(KEYINPUT33), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n469_), .A2(new_n205_), .A3(new_n258_), .A4(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n261_), .A2(new_n471_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n467_), .A2(new_n468_), .A3(new_n473_), .A4(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n392_), .A2(KEYINPUT32), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n451_), .A2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n476_), .B2(new_n388_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n262_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n461_), .B1(new_n475_), .B2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n312_), .B1(new_n460_), .B2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n458_), .A2(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT10), .B(G99gat), .Z(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT64), .ZN(new_n484_));
  INV_X1    g283(.A(G106gat), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n487_), .B(KEYINPUT6), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT9), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n489_), .A2(KEYINPUT65), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(G85gat), .A3(G92gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n489_), .A2(KEYINPUT65), .ZN(new_n492_));
  OR2_X1    g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G85gat), .B(G92gat), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n488_), .B(new_n491_), .C1(new_n493_), .C2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n486_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT66), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n494_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT8), .ZN(new_n499_));
  NOR2_X1   g298(.A1(G99gat), .A2(G106gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT7), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n488_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n498_), .A2(new_n499_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT67), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n498_), .A2(KEYINPUT67), .A3(new_n499_), .A4(new_n502_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n488_), .A2(KEYINPUT68), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n488_), .A2(KEYINPUT68), .ZN(new_n509_));
  INV_X1    g308(.A(new_n501_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n498_), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT8), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n496_), .B1(new_n507_), .B2(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G29gat), .B(G36gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(new_n515_), .B(KEYINPUT71), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G43gat), .B(G50gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT72), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT72), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n514_), .A2(new_n521_), .A3(new_n518_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT69), .B1(new_n507_), .B2(new_n513_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n507_), .A2(new_n513_), .A3(KEYINPUT69), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n496_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n518_), .B(KEYINPUT15), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n520_), .B(new_n522_), .C1(new_n526_), .C2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT35), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G190gat), .B(G218gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G134gat), .B(G162gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n529_), .A2(new_n530_), .B1(KEYINPUT36), .B2(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G232gat), .A2(G233gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n535_), .B(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n529_), .B2(KEYINPUT73), .ZN(new_n539_));
  AND2_X1   g338(.A1(new_n520_), .A2(new_n522_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n496_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n525_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n541_), .B1(new_n542_), .B2(new_n523_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n527_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT73), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n540_), .A2(new_n544_), .A3(new_n545_), .A4(new_n537_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n534_), .A2(new_n539_), .A3(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n533_), .A2(KEYINPUT36), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n548_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n534_), .A2(new_n539_), .A3(new_n546_), .A4(new_n550_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n549_), .A2(KEYINPUT37), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT37), .B1(new_n549_), .B2(new_n551_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G15gat), .B(G22gat), .ZN(new_n555_));
  INV_X1    g354(.A(G1gat), .ZN(new_n556_));
  INV_X1    g355(.A(G8gat), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT14), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n555_), .A2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G1gat), .B(G8gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n559_), .B(new_n560_), .Z(new_n561_));
  NAND2_X1  g360(.A1(G231gat), .A2(G233gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G57gat), .B(G64gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT11), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G71gat), .B(G78gat), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n564_), .A2(KEYINPUT11), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n570_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n563_), .B(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT17), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G127gat), .B(G155gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT16), .ZN(new_n575_));
  XOR2_X1   g374(.A(G183gat), .B(G211gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n572_), .B1(new_n573_), .B2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(KEYINPUT17), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n578_), .B1(new_n572_), .B2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT74), .Z(new_n581_));
  NOR2_X1   g380(.A1(new_n554_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n561_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n527_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n518_), .A2(new_n561_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G229gat), .A2(G233gat), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n518_), .B(new_n561_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n586_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G113gat), .B(G141gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(G169gat), .B(G197gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n591_), .B(new_n594_), .Z(new_n595_));
  INV_X1    g394(.A(KEYINPUT13), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n507_), .A2(new_n513_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n541_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n571_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT12), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n599_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n600_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n543_), .A2(KEYINPUT12), .A3(new_n599_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(G230gat), .ZN(new_n606_));
  INV_X1    g405(.A(G233gat), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n602_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n608_), .B1(new_n611_), .B2(new_n600_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT5), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G176gat), .B(G204gat), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n615_), .B(new_n616_), .Z(new_n617_));
  NAND2_X1  g416(.A1(new_n613_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n617_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n610_), .A2(new_n612_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n618_), .B1(KEYINPUT70), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n620_), .A2(KEYINPUT70), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n619_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n596_), .B1(new_n621_), .B2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n622_), .A2(new_n623_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n618_), .A2(KEYINPUT70), .A3(new_n620_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n627_), .A3(KEYINPUT13), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n625_), .A2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n482_), .A2(new_n582_), .A3(new_n595_), .A4(new_n629_), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n630_), .B(KEYINPUT102), .Z(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT103), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n556_), .A3(new_n262_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n312_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n473_), .A2(new_n474_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n464_), .A2(new_n462_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n465_), .A2(new_n466_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n468_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n479_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(new_n450_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n456_), .A2(new_n459_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n636_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n423_), .A2(new_n450_), .A3(new_n454_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT101), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n456_), .A2(new_n314_), .A3(new_n450_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n644_), .B1(new_n648_), .B2(new_n313_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n549_), .A2(new_n551_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT105), .ZN(new_n653_));
  INV_X1    g452(.A(new_n581_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n629_), .A2(new_n595_), .A3(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n655_), .B(KEYINPUT104), .Z(new_n656_));
  AND3_X1   g455(.A1(new_n653_), .A2(new_n656_), .A3(KEYINPUT106), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT106), .B1(new_n653_), .B2(new_n656_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n262_), .ZN(new_n660_));
  OAI21_X1  g459(.A(G1gat), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n633_), .A2(new_n634_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n635_), .A2(new_n661_), .A3(new_n662_), .ZN(G1324gat));
  INV_X1    g462(.A(new_n456_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n632_), .A2(new_n557_), .A3(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n653_), .A2(new_n656_), .A3(new_n664_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(G8gat), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n667_), .A2(KEYINPUT39), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(KEYINPUT39), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n665_), .B(KEYINPUT40), .C1(new_n668_), .C2(new_n669_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1325gat));
  OAI21_X1  g473(.A(G15gat), .B1(new_n659_), .B2(new_n312_), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n675_), .A2(KEYINPUT41), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(KEYINPUT41), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n631_), .A2(new_n306_), .A3(new_n636_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT107), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n676_), .A2(new_n677_), .A3(new_n679_), .ZN(G1326gat));
  INV_X1    g479(.A(G22gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n631_), .A2(new_n681_), .A3(new_n461_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n461_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(new_n684_), .A3(G22gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n683_), .B2(G22gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(G1327gat));
  INV_X1    g486(.A(new_n595_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n649_), .A2(new_n688_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n650_), .A2(new_n654_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n689_), .A2(new_n629_), .A3(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(G29gat), .B1(new_n692_), .B2(new_n262_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n552_), .A2(new_n553_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n649_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT43), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n482_), .A2(new_n696_), .A3(new_n554_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n695_), .A2(new_n697_), .ZN(new_n698_));
  AND4_X1   g497(.A1(new_n595_), .A2(new_n698_), .A3(new_n629_), .A4(new_n581_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT44), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n700_), .A2(G29gat), .A3(new_n262_), .ZN(new_n701_));
  XOR2_X1   g500(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n702_));
  OR2_X1    g501(.A1(new_n699_), .A2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n693_), .B1(new_n701_), .B2(new_n703_), .ZN(G1328gat));
  NOR3_X1   g503(.A1(new_n691_), .A2(G36gat), .A3(new_n456_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT45), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n703_), .A2(new_n664_), .A3(new_n700_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n707_), .B2(G36gat), .ZN(new_n708_));
  XOR2_X1   g507(.A(KEYINPUT109), .B(KEYINPUT46), .Z(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(G1329gat));
  OAI21_X1  g509(.A(new_n301_), .B1(new_n691_), .B2(new_n312_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT111), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n312_), .A2(new_n301_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n714_), .B1(new_n699_), .B2(KEYINPUT44), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n703_), .A2(KEYINPUT110), .A3(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT110), .B1(new_n703_), .B2(new_n715_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n712_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT47), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT47), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n720_), .B(new_n712_), .C1(new_n716_), .C2(new_n717_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1330gat));
  AOI21_X1  g521(.A(G50gat), .B1(new_n692_), .B2(new_n461_), .ZN(new_n723_));
  AND3_X1   g522(.A1(new_n700_), .A2(G50gat), .A3(new_n461_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n724_), .B2(new_n703_), .ZN(G1331gat));
  INV_X1    g524(.A(new_n629_), .ZN(new_n726_));
  AND4_X1   g525(.A1(new_n688_), .A2(new_n653_), .A3(new_n726_), .A4(new_n654_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n727_), .A2(G57gat), .A3(new_n262_), .ZN(new_n728_));
  NOR3_X1   g527(.A1(new_n649_), .A2(new_n595_), .A3(new_n629_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n582_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n262_), .B1(new_n730_), .B2(KEYINPUT112), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n731_), .B1(KEYINPUT112), .B2(new_n730_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n728_), .B1(G57gat), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT113), .ZN(G1332gat));
  INV_X1    g533(.A(new_n730_), .ZN(new_n735_));
  INV_X1    g534(.A(G64gat), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n664_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n727_), .B2(new_n664_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT114), .B(KEYINPUT48), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n738_), .A2(new_n739_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(G1333gat));
  INV_X1    g541(.A(G71gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n727_), .B2(new_n636_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT49), .Z(new_n745_));
  NAND3_X1  g544(.A1(new_n735_), .A2(new_n743_), .A3(new_n636_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1334gat));
  AOI21_X1  g546(.A(new_n440_), .B1(new_n727_), .B2(new_n461_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT50), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n735_), .A2(new_n440_), .A3(new_n461_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1335gat));
  NAND2_X1  g550(.A1(new_n729_), .A2(new_n690_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(G85gat), .B1(new_n753_), .B2(new_n262_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n629_), .A2(new_n595_), .A3(new_n654_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n698_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n262_), .A2(G85gat), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT115), .Z(new_n758_));
  AOI21_X1  g557(.A(new_n754_), .B1(new_n756_), .B2(new_n758_), .ZN(G1336gat));
  AOI21_X1  g558(.A(G92gat), .B1(new_n753_), .B2(new_n664_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n664_), .A2(G92gat), .ZN(new_n761_));
  XOR2_X1   g560(.A(new_n761_), .B(KEYINPUT116), .Z(new_n762_));
  AOI21_X1  g561(.A(new_n760_), .B1(new_n756_), .B2(new_n762_), .ZN(G1337gat));
  AND2_X1   g562(.A1(new_n756_), .A2(new_n636_), .ZN(new_n764_));
  INV_X1    g563(.A(G99gat), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n636_), .A2(new_n484_), .ZN(new_n766_));
  OAI22_X1  g565(.A1(new_n764_), .A2(new_n765_), .B1(new_n752_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g567(.A1(new_n753_), .A2(new_n485_), .A3(new_n461_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n696_), .B1(new_n482_), .B2(new_n554_), .ZN(new_n771_));
  AOI211_X1 g570(.A(KEYINPUT43), .B(new_n694_), .C1(new_n458_), .C2(new_n481_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n461_), .B(new_n755_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT117), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT117), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n698_), .A2(new_n775_), .A3(new_n461_), .A4(new_n755_), .ZN(new_n776_));
  AND4_X1   g575(.A1(new_n770_), .A2(new_n774_), .A3(G106gat), .A4(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n485_), .B1(new_n773_), .B2(KEYINPUT117), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n770_), .B1(new_n778_), .B2(new_n776_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n769_), .B1(new_n777_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT119), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n782_), .B(new_n769_), .C1(new_n777_), .C2(new_n779_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n781_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n781_), .B2(new_n783_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1339gat));
  INV_X1    g586(.A(KEYINPUT121), .ZN(new_n788_));
  INV_X1    g587(.A(new_n591_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n584_), .A2(new_n585_), .A3(new_n589_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n594_), .B1(new_n588_), .B2(new_n586_), .ZN(new_n791_));
  AOI22_X1  g590(.A1(new_n789_), .A2(new_n594_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT55), .B1(new_n605_), .B2(new_n609_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n610_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n605_), .A2(KEYINPUT55), .A3(new_n609_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n619_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n620_), .B(new_n792_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n798_));
  AND2_X1   g597(.A1(new_n796_), .A2(new_n797_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n788_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n694_), .B1(new_n800_), .B2(KEYINPUT58), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n801_), .B1(KEYINPUT58), .B2(new_n800_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n626_), .A2(new_n627_), .A3(new_n792_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n796_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n595_), .A3(new_n620_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n796_), .A2(new_n804_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n650_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(KEYINPUT57), .A3(new_n650_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n802_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n581_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n582_), .A2(new_n688_), .A3(new_n629_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n816_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n814_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n648_), .A2(new_n262_), .A3(new_n636_), .ZN(new_n821_));
  XOR2_X1   g620(.A(new_n821_), .B(KEYINPUT122), .Z(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n823_), .B(KEYINPUT59), .ZN(new_n824_));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824_), .B2(new_n688_), .ZN(new_n825_));
  OR2_X1    g624(.A1(new_n688_), .A2(G113gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n823_), .B2(new_n826_), .ZN(G1340gat));
  OAI21_X1  g626(.A(G120gat), .B1(new_n824_), .B2(new_n629_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n823_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT60), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(G120gat), .ZN(new_n831_));
  AOI21_X1  g630(.A(G120gat), .B1(new_n726_), .B2(new_n830_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(KEYINPUT123), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n833_), .B1(KEYINPUT123), .B2(new_n832_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n829_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n828_), .A2(new_n835_), .ZN(G1341gat));
  OAI21_X1  g635(.A(G127gat), .B1(new_n824_), .B2(new_n581_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n581_), .A2(G127gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n823_), .B2(new_n838_), .ZN(G1342gat));
  AOI21_X1  g638(.A(G134gat), .B1(new_n829_), .B2(new_n651_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n824_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT124), .B(G134gat), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n694_), .A2(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n840_), .B1(new_n841_), .B2(new_n843_), .ZN(G1343gat));
  AOI22_X1  g643(.A1(new_n813_), .A2(new_n581_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n450_), .A2(new_n636_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n845_), .A2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n664_), .A2(new_n660_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n848_), .A2(KEYINPUT125), .A3(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT125), .B1(new_n848_), .B2(new_n849_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n595_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(G141gat), .ZN(new_n853_));
  INV_X1    g652(.A(G141gat), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n854_), .B(new_n595_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1344gat));
  OAI21_X1  g655(.A(new_n726_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(G148gat), .ZN(new_n858_));
  INV_X1    g657(.A(G148gat), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n859_), .B(new_n726_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(G1345gat));
  OAI21_X1  g660(.A(new_n654_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT61), .B(G155gat), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n863_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n654_), .B(new_n865_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1346gat));
  INV_X1    g666(.A(G162gat), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n868_), .B(new_n651_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n851_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n848_), .A2(KEYINPUT125), .A3(new_n849_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n694_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n869_), .B1(new_n872_), .B2(new_n868_), .ZN(G1347gat));
  INV_X1    g672(.A(KEYINPUT62), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n664_), .A2(new_n450_), .A3(new_n313_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n845_), .A2(new_n688_), .A3(new_n875_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n874_), .B1(new_n876_), .B2(new_n263_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n875_), .B1(new_n814_), .B2(new_n819_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  OAI211_X1 g678(.A(KEYINPUT62), .B(G169gat), .C1(new_n879_), .C2(new_n688_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n372_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n876_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n877_), .A2(new_n880_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT126), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n877_), .A2(new_n880_), .A3(KEYINPUT126), .A4(new_n882_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1348gat));
  NAND2_X1  g686(.A1(new_n878_), .A2(new_n726_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT127), .B(G176gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1349gat));
  NAND2_X1  g689(.A1(new_n878_), .A2(new_n654_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n891_), .A2(new_n279_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n892_), .B1(new_n274_), .B2(new_n891_), .ZN(G1350gat));
  OAI21_X1  g692(.A(G190gat), .B1(new_n879_), .B2(new_n694_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n878_), .A2(new_n273_), .A3(new_n651_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1351gat));
  NOR4_X1   g695(.A1(new_n845_), .A2(new_n262_), .A3(new_n456_), .A4(new_n847_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n595_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g698(.A1(new_n897_), .A2(new_n726_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g700(.A(new_n581_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n897_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n904_));
  XOR2_X1   g703(.A(new_n903_), .B(new_n904_), .Z(G1354gat));
  INV_X1    g704(.A(G218gat), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n897_), .A2(new_n906_), .A3(new_n651_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n897_), .A2(new_n554_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n906_), .ZN(G1355gat));
endmodule


