//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n960_, new_n961_, new_n963_, new_n964_, new_n965_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n973_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n987_, new_n988_,
    new_n989_;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G15gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(G71gat), .ZN(new_n205_));
  INV_X1    g004(.A(G99gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT82), .B(G43gat), .Z(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT83), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n207_), .B(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G183gat), .A2(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT23), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT81), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n211_), .A2(KEYINPUT81), .A3(KEYINPUT23), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G183gat), .A3(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT24), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  AOI22_X1  g019(.A1(new_n216_), .A2(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G183gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT25), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT25), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n224_), .A2(G183gat), .ZN(new_n225_));
  INV_X1    g024(.A(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT26), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT26), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G190gat), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n223_), .A2(new_n225_), .A3(new_n227_), .A4(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n220_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G169gat), .A2(G176gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(KEYINPUT24), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n230_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT80), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n230_), .A2(new_n233_), .A3(KEYINPUT80), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n221_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n212_), .A2(new_n218_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n239_), .B1(G183gat), .B2(G190gat), .ZN(new_n240_));
  NOR2_X1   g039(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(G169gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n240_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n238_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT30), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n245_), .A2(KEYINPUT84), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(KEYINPUT84), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n210_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n248_), .B1(new_n246_), .B2(new_n210_), .ZN(new_n249_));
  INV_X1    g048(.A(G134gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G127gat), .ZN(new_n251_));
  INV_X1    g050(.A(G127gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G134gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G120gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G113gat), .ZN(new_n256_));
  INV_X1    g055(.A(G113gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G120gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n254_), .A2(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n251_), .A2(new_n253_), .A3(new_n256_), .A4(new_n258_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(KEYINPUT85), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n254_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(new_n256_), .A4(new_n258_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n262_), .A2(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n266_), .B(KEYINPUT31), .Z(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n249_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n249_), .A2(new_n268_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(G218gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(G211gat), .ZN(new_n273_));
  INV_X1    g072(.A(G211gat), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(G218gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n273_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT89), .ZN(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT21), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G211gat), .B(G218gat), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n279_), .A2(KEYINPUT89), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G197gat), .ZN(new_n282_));
  OR2_X1    g081(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(KEYINPUT88), .A2(G204gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(G197gat), .A2(G204gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n283_), .A2(new_n282_), .A3(new_n284_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT21), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n289_), .B1(G197gat), .B2(G204gat), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n276_), .B1(new_n288_), .B2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n292_));
  AOI22_X1  g091(.A1(new_n281_), .A2(new_n287_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  NOR2_X1   g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G141gat), .A2(G148gat), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT2), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(KEYINPUT87), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT3), .ZN(new_n300_));
  INV_X1    g099(.A(G141gat), .ZN(new_n301_));
  INV_X1    g100(.A(G148gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n299_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n298_), .B1(new_n297_), .B2(KEYINPUT87), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n296_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  OR2_X1    g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n308_), .B1(KEYINPUT1), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT86), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n309_), .A2(new_n311_), .A3(KEYINPUT1), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n311_), .B1(new_n309_), .B2(KEYINPUT1), .ZN(new_n313_));
  NOR3_X1   g112(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n297_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n307_), .B1(new_n314_), .B2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n293_), .B1(KEYINPUT29), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT28), .B1(new_n319_), .B2(KEYINPUT29), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NOR3_X1   g121(.A1(new_n319_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n320_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n323_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n289_), .B1(new_n279_), .B2(KEYINPUT89), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n287_), .B(new_n326_), .C1(KEYINPUT89), .C2(new_n279_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n292_), .A2(new_n291_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n319_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT29), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n329_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n325_), .A2(new_n332_), .A3(new_n321_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n324_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G228gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(G78gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G106gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G22gat), .B(G50gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(new_n337_), .B(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n334_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n324_), .A2(new_n333_), .A3(new_n339_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n295_), .B1(new_n294_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n309_), .A2(KEYINPUT1), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT86), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n309_), .A2(new_n311_), .A3(KEYINPUT1), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n345_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n317_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n260_), .A2(new_n261_), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n350_), .A2(new_n307_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT94), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n352_), .A2(new_n353_), .B1(new_n266_), .B2(new_n319_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n350_), .A2(new_n307_), .A3(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n355_), .A2(KEYINPUT94), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n354_), .A2(new_n356_), .A3(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G1gat), .B(G29gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(G85gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT0), .B(G57gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n359_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT95), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n354_), .A2(new_n365_), .A3(KEYINPUT4), .A4(new_n356_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n319_), .A2(new_n266_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n350_), .A2(new_n353_), .A3(new_n307_), .A4(new_n351_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n356_), .A2(KEYINPUT4), .A3(new_n367_), .A4(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT95), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n367_), .A2(KEYINPUT4), .ZN(new_n372_));
  AND2_X1   g171(.A1(new_n372_), .A2(new_n357_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT96), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(KEYINPUT96), .A3(new_n373_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n364_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n354_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n372_), .A2(new_n358_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n371_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n363_), .ZN(new_n384_));
  AOI21_X1  g183(.A(KEYINPUT33), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n381_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT33), .ZN(new_n387_));
  NOR4_X1   g186(.A1(new_n386_), .A2(new_n387_), .A3(new_n380_), .A4(new_n363_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n385_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G226gat), .A2(G233gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT19), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT20), .ZN(new_n393_));
  INV_X1    g192(.A(new_n218_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n394_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(G183gat), .A2(G190gat), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n242_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n212_), .A2(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(new_n230_), .A3(new_n233_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT90), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT90), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n398_), .A2(new_n230_), .A3(new_n401_), .A4(new_n233_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n397_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n393_), .B1(new_n403_), .B2(new_n329_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n293_), .A2(new_n238_), .A3(new_n243_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n392_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n392_), .B1(new_n403_), .B2(new_n329_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n238_), .A2(new_n243_), .B1(new_n328_), .B2(new_n327_), .ZN(new_n408_));
  NOR3_X1   g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n393_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT91), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n406_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G8gat), .B(G36gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G64gat), .B(G92gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n243_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n230_), .A2(new_n233_), .A3(KEYINPUT80), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT80), .B1(new_n230_), .B2(new_n233_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n418_), .B1(new_n421_), .B2(new_n221_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT20), .B1(new_n422_), .B2(new_n293_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT91), .B1(new_n423_), .B2(new_n407_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n411_), .A2(new_n417_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n393_), .B1(new_n244_), .B2(new_n329_), .ZN(new_n426_));
  OR2_X1    g225(.A1(new_n403_), .A2(new_n329_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(new_n410_), .A4(new_n392_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n404_), .A2(new_n405_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n391_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n424_), .A2(new_n428_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n416_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n425_), .A2(new_n432_), .A3(KEYINPUT93), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT93), .B1(new_n425_), .B2(new_n432_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n379_), .B(new_n389_), .C1(new_n434_), .C2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n380_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n369_), .B(new_n365_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n437_), .B(new_n384_), .C1(new_n438_), .C2(new_n381_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n363_), .B1(new_n386_), .B2(new_n380_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n327_), .A2(new_n397_), .A3(new_n328_), .A4(new_n399_), .ZN(new_n442_));
  OAI211_X1 g241(.A(KEYINPUT20), .B(new_n442_), .C1(new_n422_), .C2(new_n293_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n391_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n404_), .A2(new_n392_), .A3(new_n405_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n417_), .A2(KEYINPUT32), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n448_), .B1(new_n431_), .B2(new_n447_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n441_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n343_), .B1(new_n436_), .B2(new_n451_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n439_), .A2(new_n440_), .A3(new_n343_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT97), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n454_), .B1(new_n446_), .B2(new_n416_), .ZN(new_n455_));
  AOI211_X1 g254(.A(KEYINPUT97), .B(new_n417_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n456_));
  OAI211_X1 g255(.A(KEYINPUT27), .B(new_n425_), .C1(new_n455_), .C2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT27), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n417_), .B1(new_n411_), .B2(new_n424_), .ZN(new_n459_));
  AND4_X1   g258(.A1(new_n417_), .A2(new_n424_), .A3(new_n430_), .A4(new_n428_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n458_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n453_), .A2(new_n457_), .A3(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT98), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT98), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n453_), .A2(new_n457_), .A3(new_n461_), .A4(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n271_), .B1(new_n452_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT99), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n441_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n271_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n343_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n457_), .A2(new_n461_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  OAI211_X1 g274(.A(KEYINPUT99), .B(new_n271_), .C1(new_n452_), .C2(new_n466_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n469_), .A2(new_n475_), .A3(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G229gat), .A2(G233gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G1gat), .B(G8gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(KEYINPUT75), .B(G15gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(G22gat), .ZN(new_n482_));
  INV_X1    g281(.A(G1gat), .ZN(new_n483_));
  INV_X1    g282(.A(G8gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT14), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(KEYINPUT76), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT76), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n482_), .A2(new_n488_), .A3(new_n485_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n480_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n487_), .A2(new_n480_), .A3(new_n489_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G29gat), .B(G36gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT71), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G43gat), .B(G50gat), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT71), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n493_), .B(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(new_n495_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n491_), .A2(new_n492_), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n501_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n479_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n492_), .ZN(new_n506_));
  NOR2_X1   g305(.A1(new_n506_), .A2(new_n490_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n508_), .B1(new_n497_), .B2(new_n500_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n499_), .A2(new_n495_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n494_), .A2(new_n496_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT15), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n509_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n507_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n501_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(new_n506_), .B2(new_n490_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n516_), .A3(new_n478_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n505_), .A2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G113gat), .B(G141gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G169gat), .B(G197gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n519_), .B(new_n520_), .Z(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n505_), .A2(new_n517_), .A3(new_n521_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n477_), .A2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(KEYINPUT78), .B(KEYINPUT17), .Z(new_n527_));
  XOR2_X1   g326(.A(G127gat), .B(G155gat), .Z(new_n528_));
  XNOR2_X1  g327(.A(G183gat), .B(G211gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT77), .B(KEYINPUT16), .Z(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n507_), .A2(G231gat), .A3(G233gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G231gat), .A2(G233gat), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n506_), .B2(new_n490_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G57gat), .B(G64gat), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n537_), .A2(KEYINPUT11), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(KEYINPUT11), .ZN(new_n539_));
  XOR2_X1   g338(.A(G71gat), .B(G78gat), .Z(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n539_), .A2(new_n540_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n536_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n527_), .B(new_n532_), .C1(new_n544_), .C2(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n547_), .A2(KEYINPUT79), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(KEYINPUT79), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT68), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n541_), .A2(new_n550_), .A3(new_n542_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n550_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n536_), .B(new_n554_), .Z(new_n555_));
  XOR2_X1   g354(.A(new_n532_), .B(KEYINPUT17), .Z(new_n556_));
  AOI22_X1  g355(.A1(new_n548_), .A2(new_n549_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G230gat), .A2(G233gat), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT65), .B(G85gat), .ZN(new_n561_));
  INV_X1    g360(.A(G92gat), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  OAI22_X1  g362(.A1(KEYINPUT64), .A2(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n564_), .B1(KEYINPUT64), .B2(KEYINPUT9), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n560_), .B1(new_n563_), .B2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT6), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(G106gat), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT10), .B(G99gat), .Z(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n566_), .A2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT66), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n566_), .A2(new_n572_), .A3(KEYINPUT66), .ZN(new_n576_));
  XOR2_X1   g375(.A(G85gat), .B(G92gat), .Z(new_n577_));
  NOR2_X1   g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT7), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n577_), .B1(new_n580_), .B2(new_n569_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT8), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n582_), .A2(KEYINPUT67), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n581_), .A2(new_n583_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n575_), .A2(new_n576_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n554_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n586_), .A2(new_n554_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n559_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT12), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n591_), .B1(new_n586_), .B2(new_n554_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n575_), .A2(new_n576_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n584_), .A2(new_n585_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n545_), .A2(KEYINPUT12), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n592_), .A2(new_n598_), .A3(new_n558_), .A4(new_n587_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G120gat), .B(G148gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT5), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G176gat), .B(G204gat), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(new_n602_), .Z(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n590_), .A2(new_n599_), .A3(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT69), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT69), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n590_), .A2(new_n599_), .A3(new_n607_), .A4(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n590_), .A2(new_n599_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(new_n603_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT70), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n612_), .B1(new_n613_), .B2(KEYINPUT13), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n613_), .A2(KEYINPUT13), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n613_), .A2(KEYINPUT13), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n609_), .B(new_n611_), .C1(new_n615_), .C2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n509_), .A2(new_n512_), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT73), .B1(new_n619_), .B2(new_n586_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G232gat), .A2(G233gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT34), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n622_), .A2(KEYINPUT35), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n622_), .A2(KEYINPUT35), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n624_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT72), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n628_), .B1(new_n595_), .B2(new_n501_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n586_), .A2(KEYINPUT72), .A3(new_n515_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n513_), .A2(new_n595_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n629_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n627_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n629_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(new_n624_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(G190gat), .B(G218gat), .ZN(new_n636_));
  XNOR2_X1  g435(.A(G134gat), .B(G162gat), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n638_), .A2(KEYINPUT36), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n633_), .A2(new_n635_), .A3(new_n639_), .ZN(new_n640_));
  AND2_X1   g439(.A1(new_n634_), .A2(new_n624_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n625_), .B1(new_n620_), .B2(new_n623_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(new_n634_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT74), .B1(new_n641_), .B2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n638_), .A2(KEYINPUT36), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n635_), .B1(new_n634_), .B2(new_n642_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n648_), .A2(KEYINPUT74), .A3(new_n645_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n640_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT37), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n640_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n648_), .A2(KEYINPUT74), .A3(new_n645_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n645_), .B1(new_n648_), .B2(KEYINPUT74), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n653_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(KEYINPUT37), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n557_), .A2(new_n618_), .A3(new_n652_), .A4(new_n657_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n526_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT100), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT100), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n659_), .A2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n470_), .A2(new_n483_), .ZN(new_n665_));
  XOR2_X1   g464(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  OR3_X1    g466(.A1(new_n664_), .A2(new_n665_), .A3(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n656_), .B(KEYINPUT102), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n477_), .A2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n618_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n525_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n557_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n671_), .A2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G1gat), .B1(new_n677_), .B2(new_n441_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n668_), .A2(new_n669_), .A3(new_n678_), .ZN(G1324gat));
  NAND4_X1  g478(.A1(new_n661_), .A2(new_n484_), .A3(new_n473_), .A4(new_n663_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT39), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n671_), .A2(new_n473_), .A3(new_n676_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(G8gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n681_), .A3(G8gat), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n680_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n680_), .B(KEYINPUT40), .C1(new_n683_), .C2(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1325gat));
  INV_X1    g489(.A(new_n271_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n660_), .A2(new_n203_), .A3(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n671_), .A2(new_n691_), .A3(new_n676_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT41), .B1(new_n693_), .B2(G15gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n692_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT103), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(G1326gat));
  OAI21_X1  g498(.A(G22gat), .B1(new_n677_), .B2(new_n472_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT42), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n472_), .A2(G22gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n659_), .B2(new_n702_), .ZN(G1327gat));
  INV_X1    g502(.A(new_n557_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(new_n656_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n705_), .A2(new_n672_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n477_), .A2(new_n525_), .A3(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(G29gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n470_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n652_), .A2(new_n657_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n476_), .A2(new_n475_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT93), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n713_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n378_), .B1(new_n714_), .B2(new_n433_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n450_), .B1(new_n715_), .B2(new_n389_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n463_), .B(new_n465_), .C1(new_n716_), .C2(new_n343_), .ZN(new_n717_));
  AOI21_X1  g516(.A(KEYINPUT99), .B1(new_n717_), .B2(new_n271_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n711_), .B1(new_n712_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT43), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n477_), .A2(new_n721_), .A3(new_n711_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  OAI211_X1 g522(.A(new_n674_), .B(new_n704_), .C1(KEYINPUT105), .C2(KEYINPUT44), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT104), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT105), .B1(new_n727_), .B2(KEYINPUT44), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n726_), .A2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n723_), .A2(new_n725_), .A3(new_n728_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n441_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n710_), .B1(new_n732_), .B2(new_n709_), .ZN(G1328gat));
  INV_X1    g532(.A(KEYINPUT46), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n728_), .B1(new_n723_), .B2(new_n725_), .ZN(new_n735_));
  AOI211_X1 g534(.A(new_n724_), .B(new_n729_), .C1(new_n720_), .C2(new_n722_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n473_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n738_), .A2(G36gat), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n477_), .A2(new_n525_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n474_), .A2(G36gat), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n741_), .A2(new_n742_), .A3(new_n706_), .A4(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n743_), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT45), .B1(new_n707_), .B2(new_n745_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n744_), .A2(new_n746_), .A3(new_n738_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n734_), .B1(new_n740_), .B2(new_n748_), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT46), .B(new_n747_), .C1(new_n737_), .C2(new_n739_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1329gat));
  NAND2_X1  g550(.A1(new_n691_), .A2(G43gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n753_));
  XOR2_X1   g552(.A(KEYINPUT107), .B(G43gat), .Z(new_n754_));
  OAI21_X1  g553(.A(new_n754_), .B1(new_n707_), .B2(new_n271_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  OR3_X1    g555(.A1(new_n753_), .A2(KEYINPUT47), .A3(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT47), .B1(new_n753_), .B2(new_n756_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1330gat));
  AOI21_X1  g558(.A(G50gat), .B1(new_n708_), .B2(new_n343_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n730_), .A2(new_n731_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n343_), .A2(G50gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(G1331gat));
  NAND2_X1  g562(.A1(new_n672_), .A2(new_n673_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n764_), .A2(new_n704_), .ZN(new_n765_));
  XOR2_X1   g564(.A(KEYINPUT108), .B(G57gat), .Z(new_n766_));
  NAND4_X1  g565(.A1(new_n671_), .A2(new_n470_), .A3(new_n765_), .A4(new_n766_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT109), .Z(new_n768_));
  AND2_X1   g567(.A1(new_n477_), .A2(new_n673_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n711_), .A2(new_n704_), .A3(new_n618_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(G57gat), .B1(new_n772_), .B2(new_n470_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n768_), .A2(new_n773_), .ZN(G1332gat));
  NAND2_X1  g573(.A1(new_n671_), .A2(new_n765_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G64gat), .B1(new_n775_), .B2(new_n474_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT48), .ZN(new_n777_));
  OR2_X1    g576(.A1(new_n474_), .A2(G64gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n771_), .B2(new_n778_), .ZN(G1333gat));
  OAI21_X1  g578(.A(G71gat), .B1(new_n775_), .B2(new_n271_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT49), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n271_), .A2(G71gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n781_), .B1(new_n771_), .B2(new_n782_), .ZN(G1334gat));
  OAI21_X1  g582(.A(G78gat), .B1(new_n775_), .B2(new_n472_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(KEYINPUT110), .B(KEYINPUT50), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n784_), .B(new_n785_), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n472_), .A2(G78gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n786_), .B1(new_n771_), .B2(new_n787_), .ZN(G1335gat));
  NOR2_X1   g587(.A1(new_n705_), .A2(new_n618_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n769_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(G85gat), .B1(new_n791_), .B2(new_n470_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n764_), .A2(new_n557_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n723_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n794_), .A2(new_n795_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n441_), .A2(new_n561_), .ZN(new_n799_));
  XOR2_X1   g598(.A(new_n799_), .B(KEYINPUT112), .Z(new_n800_));
  AOI21_X1  g599(.A(new_n792_), .B1(new_n798_), .B2(new_n800_), .ZN(G1336gat));
  NAND3_X1  g600(.A1(new_n791_), .A2(new_n562_), .A3(new_n473_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n796_), .A2(new_n797_), .A3(new_n474_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(new_n562_), .ZN(G1337gat));
  NAND2_X1  g603(.A1(new_n794_), .A2(new_n691_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n691_), .A2(new_n571_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n805_), .A2(G99gat), .B1(new_n791_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n807_), .B(new_n808_), .ZN(G1338gat));
  NAND3_X1  g608(.A1(new_n791_), .A2(new_n570_), .A3(new_n343_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n723_), .A2(new_n343_), .A3(new_n793_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n811_), .A2(new_n812_), .A3(G106gat), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n812_), .B1(new_n811_), .B2(G106gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n810_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT53), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n817_), .B(new_n810_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1339gat));
  NOR2_X1   g618(.A1(new_n711_), .A2(new_n704_), .ZN(new_n820_));
  XNOR2_X1  g619(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n820_), .A2(new_n673_), .A3(new_n618_), .A4(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT54), .ZN(new_n823_));
  OAI211_X1 g622(.A(KEYINPUT113), .B(new_n823_), .C1(new_n658_), .C2(new_n525_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n525_), .A2(new_n609_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(KEYINPUT56), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n599_), .A2(KEYINPUT114), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT55), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n599_), .A2(KEYINPUT114), .A3(new_n831_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n592_), .A2(new_n598_), .A3(new_n587_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n559_), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n830_), .A2(new_n832_), .A3(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n828_), .B1(new_n835_), .B2(new_n604_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n830_), .A2(new_n832_), .A3(new_n834_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n828_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n603_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n826_), .B1(new_n836_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n478_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n841_), .A2(KEYINPUT116), .A3(new_n522_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n514_), .A2(new_n516_), .A3(new_n479_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n479_), .B1(new_n516_), .B2(new_n502_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n521_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n842_), .A2(new_n843_), .A3(new_n846_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n847_), .A2(new_n524_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n848_), .A2(new_n612_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n650_), .B1(new_n840_), .B2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n837_), .A2(new_n603_), .A3(new_n838_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n838_), .B1(new_n837_), .B2(new_n603_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n525_), .B(new_n609_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n848_), .A2(new_n612_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n857_), .A2(KEYINPUT57), .A3(new_n650_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n852_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n647_), .A2(new_n649_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n651_), .B1(new_n861_), .B2(new_n653_), .ZN(new_n862_));
  AOI211_X1 g661(.A(KEYINPUT37), .B(new_n640_), .C1(new_n647_), .C2(new_n649_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n609_), .A2(new_n847_), .A3(new_n524_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT56), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n837_), .B2(new_n603_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n865_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n837_), .A2(new_n866_), .A3(new_n603_), .ZN(new_n869_));
  AOI21_X1  g668(.A(KEYINPUT58), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n860_), .B1(new_n864_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT56), .B1(new_n835_), .B2(new_n604_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n872_), .A2(new_n609_), .A3(new_n848_), .A4(new_n869_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT58), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  AOI22_X1  g674(.A1(new_n657_), .A2(new_n652_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n875_), .B1(new_n876_), .B2(KEYINPUT117), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n859_), .B1(new_n871_), .B2(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n825_), .B1(new_n878_), .B2(new_n557_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n271_), .A2(new_n343_), .A3(new_n473_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(new_n470_), .A3(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT59), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n881_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n673_), .A2(new_n257_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n257_), .B1(new_n881_), .B2(new_n673_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(KEYINPUT118), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n890_), .B(new_n257_), .C1(new_n881_), .C2(new_n673_), .ZN(new_n891_));
  AOI22_X1  g690(.A1(new_n886_), .A2(new_n887_), .B1(new_n889_), .B2(new_n891_), .ZN(G1340gat));
  AOI21_X1  g691(.A(new_n618_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n895_));
  AOI21_X1  g694(.A(G120gat), .B1(new_n672_), .B2(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n255_), .A2(KEYINPUT60), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n894_), .B1(new_n882_), .B2(new_n898_), .ZN(new_n899_));
  NOR4_X1   g698(.A1(new_n881_), .A2(KEYINPUT119), .A3(new_n896_), .A4(new_n897_), .ZN(new_n900_));
  OAI22_X1  g699(.A1(new_n893_), .A2(new_n255_), .B1(new_n899_), .B2(new_n900_), .ZN(G1341gat));
  AOI21_X1  g700(.A(G127gat), .B1(new_n882_), .B2(new_n557_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n557_), .A2(G127gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(KEYINPUT120), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n902_), .B1(new_n886_), .B2(new_n904_), .ZN(G1342gat));
  INV_X1    g704(.A(new_n670_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G134gat), .B1(new_n882_), .B2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n864_), .A2(new_n250_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(KEYINPUT121), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n907_), .B1(new_n886_), .B2(new_n909_), .ZN(G1343gat));
  NOR3_X1   g709(.A1(new_n691_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n879_), .A2(new_n470_), .A3(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n673_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(new_n301_), .ZN(G1344gat));
  NOR2_X1   g713(.A1(new_n912_), .A2(new_n618_), .ZN(new_n915_));
  XOR2_X1   g714(.A(KEYINPUT122), .B(G148gat), .Z(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(G1345gat));
  OAI21_X1  g716(.A(KEYINPUT123), .B1(new_n912_), .B2(new_n704_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n875_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n873_), .A2(new_n874_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n711_), .A2(new_n920_), .A3(KEYINPUT117), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n871_), .A2(new_n919_), .A3(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(KEYINPUT57), .B1(new_n857_), .B2(new_n650_), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n851_), .B(new_n656_), .C1(new_n855_), .C2(new_n856_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n557_), .B1(new_n922_), .B2(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n822_), .A2(new_n824_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n928_), .A2(new_n441_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n929_), .A2(new_n930_), .A3(new_n557_), .A4(new_n911_), .ZN(new_n931_));
  XNOR2_X1  g730(.A(KEYINPUT61), .B(G155gat), .ZN(new_n932_));
  AND3_X1   g731(.A1(new_n918_), .A2(new_n931_), .A3(new_n932_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n932_), .B1(new_n918_), .B2(new_n931_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n933_), .A2(new_n934_), .ZN(G1346gat));
  OAI21_X1  g734(.A(G162gat), .B1(new_n912_), .B2(new_n864_), .ZN(new_n936_));
  OR2_X1    g735(.A1(new_n670_), .A2(G162gat), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n936_), .B1(new_n912_), .B2(new_n937_), .ZN(G1347gat));
  NOR4_X1   g737(.A1(new_n271_), .A2(new_n474_), .A3(new_n343_), .A4(new_n470_), .ZN(new_n939_));
  NAND4_X1  g738(.A1(new_n879_), .A2(KEYINPUT124), .A3(new_n525_), .A4(new_n939_), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n525_), .B(new_n939_), .C1(new_n926_), .C2(new_n927_), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT124), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n940_), .A2(new_n943_), .A3(G169gat), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(KEYINPUT125), .ZN(new_n945_));
  INV_X1    g744(.A(G169gat), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n946_), .B1(new_n941_), .B2(new_n942_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n947_), .A2(new_n948_), .A3(new_n940_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n945_), .A2(KEYINPUT62), .A3(new_n949_), .ZN(new_n950_));
  XOR2_X1   g749(.A(KEYINPUT22), .B(G169gat), .Z(new_n951_));
  NOR2_X1   g750(.A1(new_n941_), .A2(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n948_), .B1(new_n947_), .B2(new_n940_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n952_), .B1(new_n953_), .B2(new_n954_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n950_), .A2(new_n955_), .ZN(G1348gat));
  AND2_X1   g755(.A1(new_n879_), .A2(new_n939_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(new_n672_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g758(.A1(new_n957_), .A2(new_n557_), .ZN(new_n960_));
  AOI21_X1  g759(.A(new_n960_), .B1(new_n223_), .B2(new_n225_), .ZN(new_n961_));
  AOI21_X1  g760(.A(new_n961_), .B1(new_n222_), .B2(new_n960_), .ZN(G1350gat));
  NAND4_X1  g761(.A1(new_n957_), .A2(new_n227_), .A3(new_n229_), .A4(new_n906_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n957_), .A2(new_n711_), .ZN(new_n964_));
  INV_X1    g763(.A(new_n964_), .ZN(new_n965_));
  OAI21_X1  g764(.A(new_n963_), .B1(new_n965_), .B2(new_n226_), .ZN(G1351gat));
  NAND3_X1  g765(.A1(new_n271_), .A2(new_n473_), .A3(new_n453_), .ZN(new_n967_));
  NOR2_X1   g766(.A1(new_n928_), .A2(new_n967_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n968_), .A2(new_n525_), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g769(.A1(new_n283_), .A2(new_n284_), .ZN(new_n971_));
  INV_X1    g770(.A(new_n971_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n968_), .A2(new_n672_), .ZN(new_n973_));
  MUX2_X1   g772(.A(new_n972_), .B(G204gat), .S(new_n973_), .Z(G1353gat));
  INV_X1    g773(.A(new_n967_), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n704_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n976_));
  XOR2_X1   g775(.A(new_n976_), .B(KEYINPUT126), .Z(new_n977_));
  NAND3_X1  g776(.A1(new_n879_), .A2(new_n975_), .A3(new_n977_), .ZN(new_n978_));
  INV_X1    g777(.A(KEYINPUT127), .ZN(new_n979_));
  XNOR2_X1  g778(.A(new_n978_), .B(new_n979_), .ZN(new_n980_));
  NOR2_X1   g779(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n981_));
  NAND2_X1  g780(.A1(new_n980_), .A2(new_n981_), .ZN(new_n982_));
  XNOR2_X1  g781(.A(new_n978_), .B(KEYINPUT127), .ZN(new_n983_));
  INV_X1    g782(.A(new_n981_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n983_), .A2(new_n984_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n982_), .A2(new_n985_), .ZN(G1354gat));
  NAND3_X1  g785(.A1(new_n968_), .A2(new_n272_), .A3(new_n906_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n968_), .A2(new_n711_), .ZN(new_n988_));
  INV_X1    g787(.A(new_n988_), .ZN(new_n989_));
  OAI21_X1  g788(.A(new_n987_), .B1(new_n989_), .B2(new_n272_), .ZN(G1355gat));
endmodule


