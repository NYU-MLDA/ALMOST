//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n793_, new_n794_, new_n795_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n944_, new_n945_, new_n946_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n956_,
    new_n957_, new_n958_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_, new_n970_;
  INV_X1    g000(.A(G22gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT84), .ZN(new_n203_));
  INV_X1    g002(.A(G155gat), .ZN(new_n204_));
  INV_X1    g003(.A(G162gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT1), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n206_), .A2(new_n208_), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT85), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT85), .ZN(new_n212_));
  NAND4_X1  g011(.A1(new_n206_), .A2(new_n208_), .A3(new_n212_), .A4(new_n209_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n211_), .B(new_n213_), .C1(KEYINPUT1), .C2(new_n207_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(G141gat), .ZN(new_n216_));
  INV_X1    g015(.A(G148gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT29), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n206_), .A2(new_n209_), .A3(new_n207_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT87), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT87), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n206_), .A2(new_n223_), .A3(new_n209_), .A4(new_n207_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n216_), .A2(new_n217_), .A3(KEYINPUT86), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227_));
  AOI22_X1  g026(.A1(new_n226_), .A2(KEYINPUT3), .B1(new_n227_), .B2(new_n215_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n228_), .B(new_n229_), .C1(KEYINPUT3), .C2(new_n226_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT88), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n225_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n231_), .B1(new_n225_), .B2(new_n230_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n219_), .B(new_n220_), .C1(new_n232_), .C2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT28), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n225_), .A2(new_n230_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT88), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n225_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT28), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n239_), .A2(new_n240_), .A3(new_n220_), .A4(new_n219_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n202_), .B1(new_n235_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n235_), .A2(new_n241_), .A3(new_n202_), .ZN(new_n244_));
  AOI21_X1  g043(.A(G50gat), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n244_), .ZN(new_n246_));
  INV_X1    g045(.A(G50gat), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n242_), .ZN(new_n248_));
  OAI21_X1  g047(.A(KEYINPUT89), .B1(new_n245_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT90), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT21), .ZN(new_n251_));
  INV_X1    g050(.A(G204gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G197gat), .ZN(new_n253_));
  INV_X1    g052(.A(G197gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(G204gat), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n251_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G211gat), .B(G218gat), .Z(new_n257_));
  AOI21_X1  g056(.A(new_n250_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n256_), .A2(new_n257_), .A3(new_n250_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n253_), .A2(new_n255_), .A3(new_n251_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n256_), .A2(new_n257_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n259_), .A2(new_n260_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n239_), .A2(new_n219_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(KEYINPUT29), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G228gat), .A2(G233gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n220_), .B1(new_n239_), .B2(new_n219_), .ZN(new_n268_));
  OAI211_X1 g067(.A(G228gat), .B(G233gat), .C1(new_n268_), .C2(new_n263_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n267_), .A2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT91), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G78gat), .B(G106gat), .Z(new_n273_));
  INV_X1    g072(.A(new_n273_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n267_), .A2(KEYINPUT91), .A3(new_n269_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n272_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n270_), .A2(new_n271_), .A3(new_n273_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n243_), .A2(G50gat), .A3(new_n244_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n247_), .B1(new_n246_), .B2(new_n242_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT89), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n249_), .A2(new_n276_), .A3(new_n277_), .A4(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G226gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT19), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT23), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n287_), .B(new_n288_), .C1(G183gat), .C2(G190gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT22), .ZN(new_n291_));
  INV_X1    g090(.A(G169gat), .ZN(new_n292_));
  INV_X1    g091(.A(G176gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n291_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n289_), .A2(new_n290_), .A3(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n292_), .A2(new_n293_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n287_), .B(new_n288_), .C1(new_n296_), .C2(KEYINPUT24), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n297_), .B(KEYINPUT81), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT25), .B(G183gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT26), .B(G190gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(G169gat), .A2(G176gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n296_), .A2(KEYINPUT24), .A3(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n295_), .B1(new_n298_), .B2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT20), .B1(new_n306_), .B2(new_n263_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n262_), .A2(new_n261_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n260_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n308_), .B1(new_n309_), .B2(new_n258_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n291_), .A2(new_n292_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT94), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT94), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n311_), .A2(new_n315_), .A3(new_n312_), .ZN(new_n316_));
  AOI21_X1  g115(.A(G176gat), .B1(new_n314_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n289_), .A2(new_n302_), .ZN(new_n318_));
  OAI22_X1  g117(.A1(new_n317_), .A2(new_n318_), .B1(new_n304_), .B2(new_n297_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n310_), .A2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n284_), .B1(new_n307_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n306_), .A2(new_n263_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT95), .ZN(new_n323_));
  AND3_X1   g122(.A1(new_n310_), .A2(new_n319_), .A3(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n323_), .B1(new_n310_), .B2(new_n319_), .ZN(new_n325_));
  OAI211_X1 g124(.A(KEYINPUT20), .B(new_n322_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n284_), .B(KEYINPUT93), .Z(new_n327_));
  OAI21_X1  g126(.A(new_n321_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT99), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G64gat), .B(G92gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n328_), .A2(new_n329_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n326_), .A2(new_n327_), .ZN(new_n337_));
  OR3_X1    g136(.A1(new_n307_), .A2(new_n284_), .A3(new_n320_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n334_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n329_), .B1(new_n328_), .B2(new_n335_), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT27), .B1(new_n340_), .B2(new_n341_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n337_), .A2(new_n338_), .A3(new_n334_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n334_), .B1(new_n337_), .B2(new_n338_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT27), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n342_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n270_), .A2(KEYINPUT92), .A3(new_n274_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n274_), .A2(KEYINPUT92), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n267_), .A2(new_n269_), .A3(new_n350_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n349_), .A2(new_n351_), .A3(new_n278_), .A4(new_n279_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n282_), .A2(new_n348_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT100), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(KEYINPUT97), .B(G85gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(G1gat), .B(G29gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT0), .B(G57gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361_));
  INV_X1    g160(.A(G113gat), .ZN(new_n362_));
  OR2_X1    g161(.A1(G127gat), .A2(G134gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(G127gat), .A2(G134gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT82), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT82), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n363_), .A2(new_n367_), .A3(new_n364_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n362_), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n366_), .A2(new_n362_), .A3(new_n368_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n370_), .A2(G120gat), .A3(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(G120gat), .B1(new_n370_), .B2(new_n371_), .ZN(new_n373_));
  OR2_X1    g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n264_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n372_), .A2(new_n373_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n376_), .A2(new_n239_), .A3(new_n219_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n375_), .A2(KEYINPUT4), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT4), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n264_), .A3(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n361_), .B1(new_n378_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n361_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n375_), .B2(new_n377_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n360_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n381_), .A2(new_n360_), .A3(new_n383_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n306_), .B(KEYINPUT30), .ZN(new_n388_));
  XOR2_X1   g187(.A(G71gat), .B(G99gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT83), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n388_), .B(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(G15gat), .B(G43gat), .Z(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(KEYINPUT31), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n391_), .B(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(G227gat), .A2(G233gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n374_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n394_), .B(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n282_), .A2(new_n348_), .A3(KEYINPUT100), .A4(new_n352_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n355_), .A2(new_n387_), .A3(new_n397_), .A4(new_n398_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n343_), .A2(new_n344_), .A3(KEYINPUT27), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n328_), .A2(new_n335_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT99), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(new_n339_), .A3(new_n336_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n400_), .B1(new_n403_), .B2(KEYINPUT27), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n282_), .B2(new_n352_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n282_), .A2(new_n352_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n328_), .A2(KEYINPUT32), .A3(new_n334_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n334_), .A2(KEYINPUT32), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n337_), .A2(new_n338_), .A3(new_n408_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n407_), .B(new_n409_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT33), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n384_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n378_), .A2(new_n361_), .A3(new_n380_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT98), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n360_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n375_), .A2(new_n382_), .A3(new_n377_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n378_), .A2(KEYINPUT98), .A3(new_n361_), .A4(new_n380_), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n415_), .A2(new_n416_), .A3(new_n417_), .A4(new_n418_), .ZN(new_n419_));
  OAI211_X1 g218(.A(KEYINPUT33), .B(new_n360_), .C1(new_n381_), .C2(new_n383_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n412_), .A2(new_n419_), .A3(new_n345_), .A4(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n410_), .A2(new_n421_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n405_), .A2(new_n387_), .B1(new_n406_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n399_), .B1(new_n423_), .B2(new_n397_), .ZN(new_n424_));
  OAI21_X1  g223(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  AND3_X1   g227(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n429_));
  AOI21_X1  g228(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT67), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G99gat), .A2(G106gat), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT67), .ZN(new_n435_));
  NAND3_X1  g234(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n428_), .A2(new_n431_), .A3(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(G85gat), .A2(G92gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G85gat), .A2(G92gat), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT8), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT8), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT66), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n446_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n434_), .A2(KEYINPUT66), .A3(new_n436_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n428_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n443_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n447_), .A2(new_n448_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT10), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n453_), .A2(G99gat), .ZN(new_n454_));
  INV_X1    g253(.A(G99gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(KEYINPUT10), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT64), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(KEYINPUT10), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n453_), .A2(G99gat), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT64), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n457_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G106gat), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n452_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n440_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT65), .B1(new_n465_), .B2(KEYINPUT9), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(KEYINPUT9), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT65), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT9), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n440_), .A2(new_n468_), .A3(new_n469_), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n466_), .A2(new_n467_), .A3(new_n470_), .A4(new_n439_), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT70), .B1(new_n464_), .B2(new_n471_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n460_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n463_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n447_), .A2(new_n448_), .ZN(new_n476_));
  AND4_X1   g275(.A1(KEYINPUT70), .A2(new_n475_), .A3(new_n476_), .A4(new_n471_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n451_), .B1(new_n472_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT69), .ZN(new_n479_));
  INV_X1    g278(.A(G78gat), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n480_), .A2(G71gat), .ZN(new_n481_));
  INV_X1    g280(.A(G71gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n482_), .A2(G78gat), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n479_), .B(KEYINPUT11), .C1(new_n481_), .C2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G71gat), .B(G78gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT11), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT69), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(G57gat), .A2(G64gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G57gat), .A2(G64gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(KEYINPUT68), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT68), .ZN(new_n491_));
  AND2_X1   g290(.A1(G57gat), .A2(G64gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(G57gat), .A2(G64gat), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  NOR3_X1   g294(.A1(new_n481_), .A2(new_n483_), .A3(KEYINPUT11), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n484_), .B(new_n487_), .C1(new_n495_), .C2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n487_), .A2(new_n484_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n490_), .A2(new_n494_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n501_), .A2(KEYINPUT12), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n478_), .A2(new_n502_), .ZN(new_n503_));
  AOI22_X1  g302(.A1(new_n442_), .A2(KEYINPUT8), .B1(new_n449_), .B2(new_n445_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n475_), .A2(new_n476_), .A3(new_n471_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n501_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G230gat), .A2(G233gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n504_), .A2(new_n506_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n501_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n503_), .A2(new_n509_), .A3(new_n510_), .A4(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT72), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  AOI22_X1  g315(.A1(new_n478_), .A2(new_n502_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n517_), .A2(KEYINPUT72), .A3(new_n510_), .A4(new_n509_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n513_), .A2(new_n507_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(G230gat), .A3(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G120gat), .B(G148gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT5), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(G176gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(new_n252_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n519_), .A2(new_n521_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n526_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT13), .Z(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(G29gat), .ZN(new_n533_));
  INV_X1    g332(.A(G36gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(G43gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G29gat), .A2(G36gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n536_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n247_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n535_), .A2(new_n537_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(G43gat), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(G50gat), .A3(new_n538_), .ZN(new_n544_));
  AND3_X1   g343(.A1(new_n541_), .A2(KEYINPUT15), .A3(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(KEYINPUT15), .B1(new_n541_), .B2(new_n544_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(KEYINPUT75), .B(G8gat), .Z(new_n549_));
  INV_X1    g348(.A(G1gat), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT14), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G15gat), .B(G22gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(G1gat), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n554_), .A2(G8gat), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(G8gat), .ZN(new_n557_));
  INV_X1    g356(.A(new_n555_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n550_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n557_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n548_), .A2(new_n556_), .A3(new_n560_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n539_), .A2(new_n247_), .A3(new_n540_), .ZN(new_n562_));
  AOI21_X1  g361(.A(G50gat), .B1(new_n543_), .B2(new_n538_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n558_), .A2(new_n559_), .A3(new_n557_), .ZN(new_n565_));
  AOI21_X1  g364(.A(G8gat), .B1(new_n554_), .B2(new_n555_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G229gat), .A2(G233gat), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n561_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT80), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT79), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT78), .ZN(new_n572_));
  INV_X1    g371(.A(new_n564_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n560_), .A2(new_n556_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n560_), .B2(new_n556_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n572_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n560_), .A2(new_n556_), .A3(new_n573_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n567_), .A2(KEYINPUT78), .A3(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n568_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n571_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  AOI211_X1 g380(.A(KEYINPUT79), .B(new_n568_), .C1(new_n576_), .C2(new_n578_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n570_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G113gat), .B(G141gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n292_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(new_n254_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n586_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n570_), .B(new_n588_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n532_), .A2(new_n591_), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n424_), .A2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT34), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n464_), .A2(KEYINPUT70), .A3(new_n471_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT70), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n505_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n547_), .B1(new_n599_), .B2(new_n451_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT73), .ZN(new_n601_));
  OAI211_X1 g400(.A(KEYINPUT35), .B(new_n595_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n478_), .A2(new_n548_), .B1(new_n511_), .B2(new_n564_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n602_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n478_), .A2(new_n548_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(KEYINPUT73), .ZN(new_n607_));
  NAND4_X1  g406(.A1(new_n607_), .A2(KEYINPUT35), .A3(new_n603_), .A4(new_n595_), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n595_), .A2(KEYINPUT35), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n605_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G190gat), .B(G218gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(G134gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(new_n205_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT36), .ZN(new_n615_));
  OR2_X1    g414(.A1(new_n610_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT74), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n614_), .A2(KEYINPUT36), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n610_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n618_), .B1(new_n610_), .B2(new_n617_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n616_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT37), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  OAI211_X1 g423(.A(KEYINPUT37), .B(new_n616_), .C1(new_n620_), .C2(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n560_), .A2(new_n556_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(new_n512_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G127gat), .B(G155gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT16), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G183gat), .B(G211gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n634_), .B(new_n635_), .Z(new_n636_));
  INV_X1    g435(.A(KEYINPUT17), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n636_), .A2(new_n637_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n630_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n638_), .B2(new_n630_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n626_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n593_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n387_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(new_n550_), .A3(new_n646_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n647_), .A2(KEYINPUT101), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(KEYINPUT101), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT38), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n622_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n424_), .A2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT102), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n655_), .A2(new_n641_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n592_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G1gat), .B1(new_n657_), .B2(new_n387_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n648_), .A2(KEYINPUT38), .A3(new_n649_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n652_), .A2(new_n658_), .A3(new_n659_), .ZN(G1324gat));
  NAND3_X1  g459(.A1(new_n645_), .A2(new_n549_), .A3(new_n404_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n655_), .A2(new_n592_), .A3(new_n641_), .A4(new_n404_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT39), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(new_n663_), .A3(G8gat), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n663_), .B1(new_n662_), .B2(G8gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n661_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n668_));
  INV_X1    g467(.A(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n669_), .ZN(new_n670_));
  OAI211_X1 g469(.A(new_n661_), .B(new_n668_), .C1(new_n665_), .C2(new_n666_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1325gat));
  INV_X1    g471(.A(new_n397_), .ZN(new_n673_));
  OR3_X1    g472(.A1(new_n644_), .A2(G15gat), .A3(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n656_), .A2(new_n592_), .A3(new_n397_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(KEYINPUT104), .B(KEYINPUT41), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT105), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n675_), .A2(G15gat), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n677_), .B1(new_n675_), .B2(G15gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n674_), .B1(new_n679_), .B2(new_n680_), .ZN(G1326gat));
  INV_X1    g480(.A(new_n406_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n645_), .A2(new_n202_), .A3(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n656_), .A2(new_n592_), .A3(new_n682_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT42), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(G22gat), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n685_), .B1(new_n684_), .B2(G22gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n683_), .B1(new_n687_), .B2(new_n688_), .ZN(G1327gat));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n691_));
  INV_X1    g490(.A(new_n626_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n424_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695_));
  INV_X1    g494(.A(new_n621_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n619_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT37), .B1(new_n697_), .B2(new_n616_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n625_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n624_), .A2(KEYINPUT106), .A3(new_n625_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n405_), .A2(new_n387_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n406_), .A2(new_n422_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(new_n673_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n702_), .B1(new_n706_), .B2(new_n399_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT107), .B1(new_n707_), .B2(new_n691_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n700_), .A2(new_n701_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n424_), .A2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n710_), .A2(new_n711_), .A3(KEYINPUT43), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n694_), .B1(new_n708_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n641_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n592_), .A2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n690_), .B1(new_n713_), .B2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n711_), .B1(new_n710_), .B2(KEYINPUT43), .ZN(new_n717_));
  AOI211_X1 g516(.A(KEYINPUT107), .B(new_n691_), .C1(new_n424_), .C2(new_n709_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n693_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n715_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(KEYINPUT44), .A3(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n716_), .A2(new_n721_), .A3(new_n646_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n722_), .A2(KEYINPUT108), .A3(G29gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT108), .B1(new_n722_), .B2(G29gat), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n653_), .A2(new_n641_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n424_), .A2(new_n592_), .A3(new_n725_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n726_), .A2(KEYINPUT109), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(KEYINPUT109), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n646_), .A2(new_n533_), .ZN(new_n730_));
  OAI22_X1  g529(.A1(new_n723_), .A2(new_n724_), .B1(new_n729_), .B2(new_n730_), .ZN(G1328gat));
  NAND3_X1  g530(.A1(new_n716_), .A2(new_n721_), .A3(new_n404_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(G36gat), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n727_), .A2(new_n534_), .A3(new_n404_), .A4(new_n728_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT45), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n733_), .A2(KEYINPUT46), .A3(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1329gat));
  NAND3_X1  g539(.A1(new_n716_), .A2(new_n721_), .A3(new_n397_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G43gat), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n727_), .A2(new_n536_), .A3(new_n397_), .A4(new_n728_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(KEYINPUT47), .A3(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1330gat));
  AND3_X1   g547(.A1(new_n716_), .A2(new_n721_), .A3(new_n682_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n682_), .A2(new_n247_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT110), .ZN(new_n751_));
  OAI22_X1  g550(.A1(new_n749_), .A2(new_n247_), .B1(new_n729_), .B2(new_n751_), .ZN(G1331gat));
  NOR2_X1   g551(.A1(new_n531_), .A2(new_n590_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n424_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(new_n643_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G57gat), .B1(new_n756_), .B2(new_n646_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n655_), .A2(new_n641_), .A3(new_n753_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n646_), .A2(G57gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n757_), .B1(new_n758_), .B2(new_n759_), .ZN(G1332gat));
  OR3_X1    g559(.A1(new_n755_), .A2(G64gat), .A3(new_n348_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n758_), .A2(new_n404_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT48), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(G64gat), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n763_), .B1(new_n762_), .B2(G64gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n761_), .B1(new_n765_), .B2(new_n766_), .ZN(G1333gat));
  NAND3_X1  g566(.A1(new_n756_), .A2(new_n482_), .A3(new_n397_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n482_), .B1(new_n758_), .B2(new_n397_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT49), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n769_), .A2(new_n770_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n768_), .B1(new_n772_), .B2(new_n773_), .ZN(G1334gat));
  NAND3_X1  g573(.A1(new_n756_), .A2(new_n480_), .A3(new_n682_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n480_), .B1(new_n758_), .B2(new_n682_), .ZN(new_n776_));
  XOR2_X1   g575(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n776_), .A2(new_n777_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n775_), .B1(new_n779_), .B2(new_n780_), .ZN(G1335gat));
  NOR3_X1   g580(.A1(new_n531_), .A2(new_n590_), .A3(new_n641_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n719_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n646_), .A2(G85gat), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT112), .Z(new_n785_));
  AND2_X1   g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT113), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n754_), .A2(new_n725_), .ZN(new_n788_));
  AOI21_X1  g587(.A(G85gat), .B1(new_n788_), .B2(new_n646_), .ZN(new_n789_));
  OR3_X1    g588(.A1(new_n786_), .A2(new_n787_), .A3(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n787_), .B1(new_n786_), .B2(new_n789_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1336gat));
  AOI21_X1  g591(.A(G92gat), .B1(new_n788_), .B2(new_n404_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n404_), .A2(G92gat), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(KEYINPUT114), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n793_), .B1(new_n783_), .B2(new_n795_), .ZN(G1337gat));
  NAND3_X1  g595(.A1(new_n788_), .A2(new_n462_), .A3(new_n397_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n783_), .A2(new_n397_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n798_), .B2(new_n455_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT51), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(new_n797_), .C1(new_n798_), .C2(new_n455_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1338gat));
  NAND3_X1  g602(.A1(new_n788_), .A2(new_n463_), .A3(new_n682_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n719_), .A2(new_n682_), .A3(new_n782_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(G106gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n805_), .B2(G106gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT53), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n811_), .B(new_n804_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1339gat));
  AND3_X1   g612(.A1(new_n355_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n579_), .A2(new_n568_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n561_), .A2(new_n567_), .A3(new_n580_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n586_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n589_), .A2(new_n817_), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n530_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n519_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT115), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n514_), .A2(new_n820_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n517_), .A2(new_n509_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(G230gat), .A3(G233gat), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n519_), .A2(KEYINPUT115), .A3(new_n820_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n823_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n830_), .A2(KEYINPUT116), .A3(new_n525_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832_));
  AOI21_X1  g631(.A(KEYINPUT56), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n528_), .B1(new_n587_), .B2(new_n589_), .ZN(new_n834_));
  AOI21_X1  g633(.A(KEYINPUT115), .B1(new_n519_), .B2(new_n820_), .ZN(new_n835_));
  AOI211_X1 g634(.A(new_n822_), .B(KEYINPUT55), .C1(new_n516_), .C2(new_n518_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n526_), .B1(new_n837_), .B2(new_n828_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n832_), .B2(KEYINPUT56), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n834_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n819_), .B1(new_n833_), .B2(new_n841_), .ZN(new_n842_));
  AND3_X1   g641(.A1(new_n842_), .A2(KEYINPUT57), .A3(new_n653_), .ZN(new_n843_));
  AOI21_X1  g642(.A(KEYINPUT57), .B1(new_n842_), .B2(new_n653_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT56), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n528_), .B1(new_n838_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n830_), .A2(new_n525_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n818_), .B1(new_n848_), .B2(KEYINPUT56), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(new_n849_), .A3(KEYINPUT118), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT58), .B1(new_n850_), .B2(KEYINPUT119), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(KEYINPUT119), .B2(KEYINPUT58), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n692_), .B1(new_n851_), .B2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n641_), .B1(new_n845_), .B2(new_n855_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n531_), .A2(new_n591_), .A3(new_n641_), .A4(new_n626_), .ZN(new_n857_));
  XOR2_X1   g656(.A(new_n857_), .B(KEYINPUT54), .Z(new_n858_));
  OAI211_X1 g657(.A(new_n646_), .B(new_n814_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n362_), .B1(new_n859_), .B2(new_n591_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT120), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT120), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n862_), .B(new_n362_), .C1(new_n859_), .C2(new_n591_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n859_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(KEYINPUT59), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n859_), .B2(KEYINPUT121), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n591_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n864_), .B1(G113gat), .B2(new_n870_), .ZN(G1340gat));
  INV_X1    g670(.A(KEYINPUT60), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n531_), .B2(G120gat), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n865_), .B(new_n873_), .C1(new_n872_), .C2(G120gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n531_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n875_));
  INV_X1    g674(.A(G120gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n874_), .B1(new_n875_), .B2(new_n876_), .ZN(G1341gat));
  AOI21_X1  g676(.A(G127gat), .B1(new_n865_), .B2(new_n641_), .ZN(new_n878_));
  INV_X1    g677(.A(G127gat), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT122), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n641_), .B2(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n881_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n879_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n878_), .B1(new_n882_), .B2(new_n883_), .ZN(G1342gat));
  AOI21_X1  g683(.A(G134gat), .B1(new_n865_), .B2(new_n622_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n626_), .B1(new_n867_), .B2(new_n869_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(G134gat), .ZN(G1343gat));
  OAI211_X1 g686(.A(new_n646_), .B(new_n348_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n406_), .A2(new_n397_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n888_), .A2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n590_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n532_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g694(.A1(new_n891_), .A2(new_n641_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(KEYINPUT61), .B(G155gat), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1346gat));
  AOI21_X1  g697(.A(G162gat), .B1(new_n891_), .B2(new_n622_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n702_), .A2(new_n205_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(KEYINPUT123), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n899_), .B1(new_n891_), .B2(new_n901_), .ZN(G1347gat));
  OAI211_X1 g701(.A(new_n406_), .B(new_n404_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n673_), .A2(new_n646_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n903_), .A2(new_n591_), .A3(new_n905_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n906_), .A2(new_n292_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n314_), .A2(new_n316_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NOR4_X1   g708(.A1(new_n903_), .A2(new_n591_), .A3(new_n909_), .A4(new_n905_), .ZN(new_n910_));
  OAI21_X1  g709(.A(KEYINPUT62), .B1(new_n907_), .B2(new_n910_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n912_), .B1(new_n906_), .B2(new_n292_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n913_), .ZN(G1348gat));
  NOR2_X1   g713(.A1(new_n903_), .A2(new_n905_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n532_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g716(.A1(new_n915_), .A2(new_n641_), .A3(new_n299_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n842_), .A2(new_n653_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT57), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n842_), .A2(KEYINPUT57), .A3(new_n653_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n835_), .A2(new_n836_), .A3(new_n827_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT56), .B1(new_n924_), .B2(new_n526_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n818_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n830_), .A2(new_n846_), .A3(new_n525_), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n925_), .A2(new_n527_), .A3(new_n926_), .A4(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT119), .B1(new_n928_), .B2(new_n852_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT58), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n854_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n626_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n714_), .B1(new_n923_), .B2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n858_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n348_), .B1(new_n934_), .B2(new_n935_), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n936_), .A2(new_n641_), .A3(new_n406_), .A4(new_n904_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(G183gat), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n918_), .A2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(KEYINPUT124), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n918_), .A2(new_n941_), .A3(new_n938_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n940_), .A2(new_n942_), .ZN(G1350gat));
  INV_X1    g742(.A(new_n915_), .ZN(new_n944_));
  OAI21_X1  g743(.A(G190gat), .B1(new_n944_), .B2(new_n626_), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n915_), .A2(new_n622_), .A3(new_n300_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n945_), .A2(new_n946_), .ZN(G1351gat));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948_));
  OAI211_X1 g747(.A(new_n387_), .B(new_n404_), .C1(new_n856_), .C2(new_n858_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n949_), .B2(new_n890_), .ZN(new_n950_));
  NAND4_X1  g749(.A1(new_n936_), .A2(KEYINPUT125), .A3(new_n387_), .A4(new_n889_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(new_n951_), .ZN(new_n952_));
  AOI21_X1  g751(.A(G197gat), .B1(new_n952_), .B2(new_n590_), .ZN(new_n953_));
  AOI211_X1 g752(.A(new_n254_), .B(new_n591_), .C1(new_n950_), .C2(new_n951_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(new_n953_), .A2(new_n954_), .ZN(G1352gat));
  NAND2_X1  g754(.A1(new_n952_), .A2(new_n532_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(G204gat), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n952_), .A2(new_n252_), .A3(new_n532_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(G1353gat));
  AOI21_X1  g758(.A(new_n714_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n952_), .A2(new_n960_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n962_));
  XNOR2_X1  g761(.A(new_n962_), .B(KEYINPUT126), .ZN(new_n963_));
  INV_X1    g762(.A(new_n963_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n961_), .A2(new_n964_), .ZN(new_n965_));
  NAND3_X1  g764(.A1(new_n952_), .A2(new_n963_), .A3(new_n960_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n965_), .A2(new_n966_), .ZN(G1354gat));
  AOI21_X1  g766(.A(G218gat), .B1(new_n952_), .B2(new_n622_), .ZN(new_n968_));
  INV_X1    g767(.A(G218gat), .ZN(new_n969_));
  AOI211_X1 g768(.A(new_n969_), .B(new_n626_), .C1(new_n950_), .C2(new_n951_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(new_n968_), .A2(new_n970_), .ZN(G1355gat));
endmodule


