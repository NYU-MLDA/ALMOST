//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n787_, new_n788_, new_n789_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n903_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n931_, new_n933_, new_n934_, new_n936_, new_n937_,
    new_n938_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n951_;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G155gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G211gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT16), .B(G183gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT17), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT70), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G231gat), .A2(G233gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n209_), .A2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n209_), .A2(new_n211_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT68), .B(G71gat), .ZN(new_n214_));
  INV_X1    g013(.A(G78gat), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n215_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G57gat), .B(G64gat), .Z(new_n218_));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n216_), .A2(new_n217_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT69), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT69), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n216_), .A2(new_n220_), .A3(new_n223_), .A4(new_n217_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n218_), .A2(new_n219_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n222_), .A2(new_n226_), .A3(new_n224_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  OR3_X1    g029(.A1(new_n212_), .A2(new_n213_), .A3(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(G1gat), .B(G8gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT76), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(G15gat), .ZN(new_n235_));
  INV_X1    g034(.A(G22gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G15gat), .A2(G22gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G1gat), .A2(G8gat), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n237_), .A2(new_n238_), .B1(KEYINPUT14), .B2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(new_n234_), .B(new_n240_), .Z(new_n241_));
  OAI21_X1  g040(.A(new_n230_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n231_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n207_), .A2(new_n208_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n241_), .B1(new_n231_), .B2(new_n242_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n202_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n246_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n248_), .A2(KEYINPUT77), .A3(new_n244_), .A4(new_n243_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G85gat), .B(G92gat), .ZN(new_n251_));
  INV_X1    g050(.A(G92gat), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n251_), .B1(KEYINPUT9), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(KEYINPUT9), .B2(new_n251_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n253_), .B(KEYINPUT66), .C1(KEYINPUT9), .C2(new_n251_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G99gat), .A2(G106gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n259_), .B(KEYINPUT6), .Z(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT10), .B(G99gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n261_), .A2(G106gat), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n258_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT67), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n251_), .A2(new_n266_), .ZN(new_n267_));
  OR3_X1    g066(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n267_), .B1(new_n260_), .B2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT8), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n265_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G29gat), .B(G36gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G43gat), .B(G50gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n274_), .B(new_n275_), .Z(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G232gat), .A2(G233gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT34), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(KEYINPUT75), .B(KEYINPUT35), .Z(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n273_), .A2(new_n277_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  AOI211_X1 g082(.A(KEYINPUT71), .B(new_n263_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT71), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(new_n258_), .B2(new_n264_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n272_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n276_), .B(KEYINPUT15), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n283_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n280_), .A2(new_n282_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G190gat), .B(G218gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G134gat), .B(G162gat), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n293_), .B(new_n294_), .Z(new_n295_));
  INV_X1    g094(.A(KEYINPUT36), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n290_), .A2(new_n291_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n292_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n295_), .B(KEYINPUT36), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n303_), .B1(new_n292_), .B2(new_n299_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT37), .B1(new_n301_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT37), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n292_), .A2(new_n299_), .ZN(new_n307_));
  OAI211_X1 g106(.A(new_n306_), .B(new_n300_), .C1(new_n307_), .C2(new_n303_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n305_), .A2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G8gat), .B(G36gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(new_n252_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT18), .B(G64gat), .ZN(new_n312_));
  XOR2_X1   g111(.A(new_n311_), .B(new_n312_), .Z(new_n313_));
  INV_X1    g112(.A(KEYINPUT93), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G226gat), .A2(G233gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G197gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT87), .ZN(new_n321_));
  INV_X1    g120(.A(G204gat), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n321_), .B1(G197gat), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(G204gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n320_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(G211gat), .A2(G218gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT88), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G211gat), .A2(G218gat), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  AND2_X1   g129(.A1(G211gat), .A2(G218gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(G211gat), .A2(G218gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT88), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n330_), .A2(new_n333_), .A3(KEYINPUT21), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n322_), .A2(G197gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n324_), .A2(new_n335_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n330_), .A2(new_n333_), .B1(new_n336_), .B2(KEYINPUT21), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT21), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n338_), .B(new_n320_), .C1(new_n323_), .C2(new_n325_), .ZN(new_n339_));
  AOI22_X1  g138(.A1(new_n326_), .A2(new_n334_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT25), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(G183gat), .ZN(new_n342_));
  INV_X1    g141(.A(G183gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT25), .ZN(new_n344_));
  AND2_X1   g143(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n342_), .B(new_n344_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT24), .ZN(new_n351_));
  INV_X1    g150(.A(G169gat), .ZN(new_n352_));
  INV_X1    g151(.A(G176gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  AND3_X1   g153(.A1(new_n347_), .A2(new_n350_), .A3(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n356_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(KEYINPUT24), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT92), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n360_), .A2(KEYINPUT92), .A3(KEYINPUT24), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n359_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G183gat), .A2(G190gat), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n368_), .B(new_n369_), .C1(G183gat), .C2(G190gat), .ZN(new_n370_));
  INV_X1    g169(.A(new_n360_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT22), .B(G169gat), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(new_n353_), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n355_), .A2(new_n365_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT20), .B1(new_n340_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(KEYINPUT83), .A2(G169gat), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n353_), .B1(new_n376_), .B2(KEYINPUT22), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT22), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(KEYINPUT83), .B2(G169gat), .ZN(new_n379_));
  OR2_X1    g178(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n381_));
  AOI21_X1  g180(.A(G183gat), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n368_), .A2(new_n369_), .ZN(new_n383_));
  OAI221_X1 g182(.A(new_n360_), .B1(new_n377_), .B2(new_n379_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n380_), .A2(KEYINPUT26), .A3(new_n381_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n346_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT80), .B1(new_n343_), .B2(KEYINPUT25), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT80), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n341_), .A3(G183gat), .ZN(new_n390_));
  AND3_X1   g189(.A1(new_n388_), .A2(new_n390_), .A3(new_n344_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n387_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n361_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n359_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n357_), .A2(new_n351_), .A3(new_n358_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n394_), .A2(new_n350_), .A3(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n384_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n337_), .A2(new_n339_), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n326_), .A2(KEYINPUT21), .A3(new_n333_), .A4(new_n330_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n318_), .B1(new_n375_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT20), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n403_), .B1(new_n340_), .B2(new_n374_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n397_), .A2(new_n400_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n404_), .A2(new_n317_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n314_), .B1(new_n402_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n373_), .A2(new_n370_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n365_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n347_), .A2(new_n350_), .A3(new_n354_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n408_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(KEYINPUT20), .B1(new_n400_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n387_), .A2(new_n391_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n383_), .B1(new_n359_), .B2(new_n393_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n395_), .A3(new_n414_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n415_), .A2(new_n384_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n412_), .A2(new_n416_), .A3(new_n318_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n417_), .A2(KEYINPUT93), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n313_), .B1(new_n407_), .B2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n403_), .B1(new_n400_), .B2(new_n411_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n340_), .A2(new_n384_), .A3(new_n415_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n317_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT93), .B1(new_n417_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n313_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n406_), .A2(new_n314_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n419_), .A2(new_n426_), .ZN(new_n427_));
  XOR2_X1   g226(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n420_), .A2(new_n421_), .A3(new_n317_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT98), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n317_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n431_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n432_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n426_), .B(KEYINPUT27), .C1(new_n435_), .C2(new_n424_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n429_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(G155gat), .ZN(new_n439_));
  INV_X1    g238(.A(G162gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(KEYINPUT85), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT85), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n442_), .B1(G155gat), .B2(G162gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G155gat), .A2(G162gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT86), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n447_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT3), .ZN(new_n449_));
  NOR3_X1   g248(.A1(new_n449_), .A2(G141gat), .A3(G148gat), .ZN(new_n450_));
  INV_X1    g249(.A(G141gat), .ZN(new_n451_));
  INV_X1    g250(.A(G148gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT3), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n448_), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT86), .ZN(new_n456_));
  NAND2_X1  g255(.A1(G141gat), .A2(G148gat), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n456_), .B1(new_n458_), .B2(KEYINPUT2), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n446_), .B1(new_n454_), .B2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT29), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n444_), .A2(KEYINPUT1), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT1), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(G155gat), .A3(G162gat), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n441_), .A2(new_n462_), .A3(new_n443_), .A4(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n451_), .A2(new_n452_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n457_), .A3(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n460_), .A2(new_n461_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(G228gat), .ZN(new_n469_));
  INV_X1    g268(.A(G233gat), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n469_), .A2(new_n470_), .A3(KEYINPUT89), .ZN(new_n471_));
  OR2_X1    g270(.A1(new_n468_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n468_), .A2(new_n471_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n474_), .A2(KEYINPUT90), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(KEYINPUT90), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G22gat), .B(G50gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT28), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n449_), .B1(G141gat), .B2(G148gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n451_), .A2(new_n452_), .A3(KEYINPUT3), .ZN(new_n483_));
  AND3_X1   g282(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n484_));
  AOI22_X1  g283(.A1(new_n482_), .A2(new_n483_), .B1(new_n484_), .B2(new_n447_), .ZN(new_n485_));
  AOI21_X1  g284(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n486_), .B1(KEYINPUT86), .B2(new_n455_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n445_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n466_), .A2(new_n457_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n441_), .A2(new_n443_), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n462_), .A2(new_n464_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n489_), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT29), .B1(new_n488_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(new_n400_), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT89), .B1(new_n469_), .B2(new_n470_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n481_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n495_), .ZN(new_n497_));
  AOI211_X1 g296(.A(KEYINPUT28), .B(new_n497_), .C1(new_n493_), .C2(new_n400_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n480_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  XOR2_X1   g298(.A(G78gat), .B(G106gat), .Z(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n461_), .B1(new_n460_), .B2(new_n467_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n495_), .B1(new_n502_), .B2(new_n340_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT28), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n494_), .A2(new_n481_), .A3(new_n495_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(new_n479_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n499_), .A2(new_n501_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n501_), .B1(new_n499_), .B2(new_n506_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n478_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n499_), .A2(new_n506_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n500_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n499_), .A2(new_n501_), .A3(new_n506_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n477_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT30), .B(G15gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT31), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n397_), .B(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(G227gat), .A2(G233gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(G127gat), .A2(G134gat), .ZN(new_n521_));
  INV_X1    g320(.A(G120gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(G113gat), .ZN(new_n523_));
  INV_X1    g322(.A(G113gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(G120gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G127gat), .A2(G134gat), .ZN(new_n526_));
  AND4_X1   g325(.A1(new_n521_), .A2(new_n523_), .A3(new_n525_), .A4(new_n526_), .ZN(new_n527_));
  AOI22_X1  g326(.A1(new_n523_), .A2(new_n525_), .B1(new_n521_), .B2(new_n526_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT84), .B(G43gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G71gat), .B(G99gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n520_), .B(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n515_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n521_), .A2(new_n526_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n523_), .A2(new_n525_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n488_), .B2(new_n492_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n460_), .A2(new_n529_), .A3(new_n467_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n539_), .A2(new_n540_), .B1(G225gat), .B2(G233gat), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n539_), .A2(new_n540_), .A3(KEYINPUT4), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT4), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n538_), .B(new_n544_), .C1(new_n488_), .C2(new_n492_), .ZN(new_n545_));
  AND2_X1   g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G225gat), .A2(G233gat), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n542_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G1gat), .B(G29gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(G85gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT0), .B(G57gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n548_), .B(new_n553_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n438_), .A2(new_n535_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n534_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT99), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n539_), .A2(new_n540_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n552_), .B1(new_n558_), .B2(new_n547_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n559_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n547_), .B1(new_n543_), .B2(new_n545_), .ZN(new_n561_));
  OAI211_X1 g360(.A(KEYINPUT33), .B(new_n553_), .C1(new_n561_), .C2(new_n541_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n560_), .B1(new_n562_), .B2(KEYINPUT94), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT94), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n548_), .A2(new_n564_), .A3(KEYINPUT33), .A4(new_n553_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n419_), .A2(new_n563_), .A3(new_n426_), .A4(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n553_), .B1(new_n561_), .B2(new_n541_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT95), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(KEYINPUT95), .B(new_n553_), .C1(new_n561_), .C2(new_n541_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT96), .B(KEYINPUT33), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AND4_X1   g372(.A1(new_n567_), .A2(new_n570_), .A3(new_n571_), .A4(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n572_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n567_), .B1(new_n575_), .B2(new_n571_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n566_), .A2(new_n574_), .A3(new_n576_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n424_), .A2(KEYINPUT32), .ZN(new_n578_));
  OR3_X1    g377(.A1(new_n407_), .A2(new_n418_), .A3(new_n578_), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n432_), .B(new_n578_), .C1(new_n433_), .C2(new_n434_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n554_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n557_), .B(new_n515_), .C1(new_n577_), .C2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n554_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n437_), .A2(new_n514_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  AND3_X1   g385(.A1(new_n419_), .A2(new_n565_), .A3(new_n426_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n575_), .A2(new_n567_), .A3(new_n571_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n570_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT97), .ZN(new_n590_));
  NAND4_X1  g389(.A1(new_n587_), .A2(new_n588_), .A3(new_n590_), .A4(new_n563_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n581_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n557_), .B1(new_n592_), .B2(new_n515_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n556_), .B1(new_n586_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT101), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n555_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n596_));
  OAI211_X1 g395(.A(KEYINPUT101), .B(new_n556_), .C1(new_n586_), .C2(new_n593_), .ZN(new_n597_));
  AOI211_X1 g396(.A(new_n250_), .B(new_n309_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n234_), .B(new_n240_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n289_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G229gat), .A2(G233gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n277_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n601_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n241_), .A2(new_n276_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n605_), .A2(KEYINPUT78), .A3(new_n602_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT78), .B1(new_n605_), .B2(new_n602_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n604_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n603_), .A2(new_n608_), .ZN(new_n609_));
  XOR2_X1   g408(.A(G169gat), .B(G197gat), .Z(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT79), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G113gat), .B(G141gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n611_), .B(new_n612_), .Z(new_n613_));
  XNOR2_X1  g412(.A(new_n609_), .B(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT70), .ZN(new_n619_));
  INV_X1    g418(.A(new_n229_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n226_), .B1(new_n222_), .B2(new_n224_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n619_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n228_), .A2(KEYINPUT70), .A3(new_n229_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n622_), .A2(new_n273_), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n273_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n618_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n622_), .A2(new_n273_), .A3(new_n623_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n228_), .A2(KEYINPUT12), .A3(new_n229_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n287_), .A2(new_n628_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n627_), .B(new_n629_), .C1(new_n625_), .C2(KEYINPUT12), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n626_), .B1(new_n630_), .B2(new_n618_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G120gat), .B(G148gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT73), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n631_), .A2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n626_), .B(new_n636_), .C1(new_n630_), .C2(new_n618_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n640_), .A2(KEYINPUT13), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(KEYINPUT13), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT74), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n598_), .A2(new_n615_), .A3(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(G1gat), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n554_), .B(KEYINPUT102), .Z(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n646_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT38), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n594_), .A2(new_n595_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n555_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n597_), .A3(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n643_), .A2(new_n614_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n301_), .A2(new_n304_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n250_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G1gat), .B1(new_n661_), .B2(new_n584_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n650_), .A2(new_n651_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n652_), .A2(new_n662_), .A3(new_n663_), .ZN(G1324gat));
  INV_X1    g463(.A(G8gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n646_), .A2(new_n665_), .A3(new_n438_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n655_), .A2(new_n438_), .A3(new_n659_), .A4(new_n656_), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n667_), .A2(KEYINPUT103), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n665_), .B1(new_n667_), .B2(KEYINPUT103), .ZN(new_n670_));
  AND3_X1   g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n669_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n666_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT40), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(G1325gat));
  OAI21_X1  g474(.A(G15gat), .B1(new_n661_), .B2(new_n556_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n676_), .A2(KEYINPUT41), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(KEYINPUT41), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n646_), .A2(new_n235_), .A3(new_n534_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(G1326gat));
  AOI21_X1  g479(.A(new_n236_), .B1(new_n660_), .B2(new_n514_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT42), .Z(new_n682_));
  NAND3_X1  g481(.A1(new_n646_), .A2(new_n236_), .A3(new_n514_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(G1327gat));
  NAND2_X1  g483(.A1(new_n250_), .A2(new_n658_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT104), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n657_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G29gat), .B1(new_n688_), .B2(new_n554_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n656_), .A2(new_n250_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n305_), .A2(new_n308_), .ZN(new_n692_));
  AOI211_X1 g491(.A(KEYINPUT43), .B(new_n692_), .C1(new_n596_), .C2(new_n597_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n655_), .B2(new_n309_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n691_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n698_), .A2(G29gat), .A3(new_n649_), .ZN(new_n699_));
  AND4_X1   g498(.A1(new_n514_), .A2(new_n584_), .A3(new_n429_), .A4(new_n436_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n514_), .B1(new_n591_), .B2(new_n581_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(new_n557_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n577_), .A2(new_n582_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT99), .B1(new_n703_), .B2(new_n514_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n534_), .B1(new_n702_), .B2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n654_), .B1(new_n705_), .B2(KEYINPUT101), .ZN(new_n706_));
  INV_X1    g505(.A(new_n597_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n309_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT43), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n655_), .A2(new_n694_), .A3(new_n309_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n690_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT44), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n689_), .B1(new_n699_), .B2(new_n712_), .ZN(G1328gat));
  NAND2_X1  g512(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(G36gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n437_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n719_), .B2(new_n712_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n657_), .A2(new_n718_), .A3(new_n438_), .A4(new_n686_), .ZN(new_n721_));
  XOR2_X1   g520(.A(KEYINPUT105), .B(KEYINPUT45), .Z(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n721_), .B(new_n723_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n714_), .B(new_n717_), .C1(new_n720_), .C2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n438_), .B1(new_n711_), .B2(KEYINPUT44), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n696_), .A2(new_n697_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G36gat), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n721_), .B(new_n722_), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n728_), .A2(new_n715_), .A3(new_n716_), .A4(new_n729_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n725_), .A2(new_n730_), .ZN(G1329gat));
  INV_X1    g530(.A(G43gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n732_), .B1(new_n687_), .B2(new_n556_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n698_), .A2(G43gat), .A3(new_n534_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n727_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT47), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT47), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n737_), .B(new_n733_), .C1(new_n734_), .C2(new_n727_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1330gat));
  NAND3_X1  g538(.A1(new_n712_), .A2(new_n698_), .A3(new_n514_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n740_), .A2(KEYINPUT107), .A3(G50gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT107), .B1(new_n740_), .B2(G50gat), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n515_), .A2(G50gat), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT108), .ZN(new_n744_));
  OAI22_X1  g543(.A1(new_n741_), .A2(new_n742_), .B1(new_n687_), .B2(new_n744_), .ZN(G1331gat));
  AND2_X1   g544(.A1(new_n641_), .A2(new_n642_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n746_), .A2(new_n615_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n598_), .A2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G57gat), .B1(new_n748_), .B2(new_n649_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n655_), .A2(new_n644_), .A3(new_n614_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(new_n659_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n750_), .A2(KEYINPUT109), .A3(new_n659_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n554_), .A2(G57gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n749_), .B1(new_n755_), .B2(new_n756_), .ZN(G1332gat));
  INV_X1    g556(.A(G64gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n748_), .A2(new_n758_), .A3(new_n438_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n753_), .A2(new_n438_), .A3(new_n754_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT48), .ZN(new_n761_));
  AND3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(G64gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n760_), .B2(G64gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(G1333gat));
  INV_X1    g563(.A(G71gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n748_), .A2(new_n765_), .A3(new_n534_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n753_), .A2(new_n534_), .A3(new_n754_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT49), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n767_), .A2(new_n768_), .A3(G71gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n767_), .B2(G71gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(G1334gat));
  NAND3_X1  g570(.A1(new_n748_), .A2(new_n215_), .A3(new_n514_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n753_), .A2(new_n514_), .A3(new_n754_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT50), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(G78gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(G78gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(G1335gat));
  NAND2_X1  g576(.A1(new_n750_), .A2(new_n686_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  AOI21_X1  g578(.A(G85gat), .B1(new_n779_), .B2(new_n649_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n709_), .A2(new_n710_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n747_), .A2(new_n250_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT110), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n554_), .A2(G85gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n780_), .B1(new_n784_), .B2(new_n785_), .ZN(G1336gat));
  AOI21_X1  g585(.A(G92gat), .B1(new_n779_), .B2(new_n438_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n438_), .A2(G92gat), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT111), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n787_), .B1(new_n784_), .B2(new_n789_), .ZN(G1337gat));
  NOR2_X1   g589(.A1(new_n556_), .A2(new_n261_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  OR3_X1    g591(.A1(new_n778_), .A2(KEYINPUT113), .A3(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT113), .B1(new_n778_), .B2(new_n792_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n781_), .A2(new_n534_), .A3(new_n783_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n796_), .A2(new_n797_), .A3(G99gat), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n796_), .B2(G99gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT51), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n802_), .B(new_n795_), .C1(new_n798_), .C2(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(G1338gat));
  OR3_X1    g603(.A1(new_n778_), .A2(G106gat), .A3(new_n515_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n781_), .A2(new_n514_), .A3(new_n783_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n806_), .A2(new_n807_), .A3(G106gat), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n806_), .B2(G106gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n805_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n805_), .B(new_n811_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(G1339gat));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816_));
  INV_X1    g615(.A(new_n250_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n817_), .A2(new_n692_), .A3(new_n614_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n816_), .B1(new_n819_), .B2(new_n746_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n818_), .A2(new_n643_), .A3(KEYINPUT54), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT55), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n630_), .B2(new_n618_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n630_), .A2(new_n618_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n630_), .A2(new_n823_), .A3(new_n618_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n637_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT56), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n830_), .B(new_n637_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n829_), .A2(new_n615_), .A3(new_n639_), .A4(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n613_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n608_), .A2(new_n603_), .A3(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n600_), .A2(new_n835_), .A3(new_n602_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n601_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n601_), .B1(new_n606_), .B2(new_n607_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(new_n613_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n834_), .B1(new_n838_), .B2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT116), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n832_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n658_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n639_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n849_), .B1(new_n828_), .B2(KEYINPUT56), .ZN(new_n850_));
  INV_X1    g649(.A(new_n841_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n831_), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n850_), .A2(KEYINPUT58), .A3(new_n831_), .A4(new_n851_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n309_), .A3(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n844_), .A2(KEYINPUT57), .A3(new_n845_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n848_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n822_), .B1(new_n858_), .B2(new_n250_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n649_), .A2(new_n437_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n860_), .A2(new_n535_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n859_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(G113gat), .B1(new_n863_), .B2(new_n615_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n863_), .B2(new_n866_), .ZN(new_n867_));
  OAI211_X1 g666(.A(KEYINPUT117), .B(KEYINPUT59), .C1(new_n859_), .C2(new_n862_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT119), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n862_), .A2(KEYINPUT118), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n862_), .A2(KEYINPUT118), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n870_), .A2(new_n866_), .A3(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n869_), .B1(new_n859_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n872_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n658_), .B1(new_n832_), .B2(new_n843_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n847_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n817_), .B1(new_n876_), .B2(new_n856_), .ZN(new_n877_));
  OAI211_X1 g676(.A(KEYINPUT119), .B(new_n874_), .C1(new_n877_), .C2(new_n822_), .ZN(new_n878_));
  AOI22_X1  g677(.A1(new_n867_), .A2(new_n868_), .B1(new_n873_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n615_), .A2(G113gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT120), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n864_), .B1(new_n879_), .B2(new_n881_), .ZN(G1340gat));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n873_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n861_), .B1(new_n877_), .B2(new_n822_), .ZN(new_n884_));
  AOI21_X1  g683(.A(KEYINPUT117), .B1(new_n884_), .B2(KEYINPUT59), .ZN(new_n885_));
  INV_X1    g684(.A(new_n868_), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n644_), .B(new_n883_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G120gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n522_), .B1(new_n746_), .B2(KEYINPUT60), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n863_), .B(new_n889_), .C1(KEYINPUT60), .C2(new_n522_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n890_), .ZN(G1341gat));
  AOI21_X1  g690(.A(G127gat), .B1(new_n863_), .B2(new_n817_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n817_), .A2(G127gat), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT121), .Z(new_n894_));
  AOI21_X1  g693(.A(new_n892_), .B1(new_n879_), .B2(new_n894_), .ZN(G1342gat));
  AOI21_X1  g694(.A(G134gat), .B1(new_n863_), .B2(new_n658_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n309_), .A2(G134gat), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n896_), .B1(new_n879_), .B2(new_n897_), .ZN(G1343gat));
  NOR4_X1   g697(.A1(new_n859_), .A2(new_n534_), .A3(new_n515_), .A4(new_n860_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n615_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT122), .B(G141gat), .Z(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1344gat));
  NAND2_X1  g701(.A1(new_n899_), .A2(new_n644_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n903_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g703(.A1(new_n899_), .A2(new_n817_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(KEYINPUT61), .B(G155gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n905_), .B(new_n906_), .ZN(G1346gat));
  AOI21_X1  g706(.A(G162gat), .B1(new_n899_), .B2(new_n658_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n692_), .A2(new_n440_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n899_), .B2(new_n909_), .ZN(G1347gat));
  NOR2_X1   g709(.A1(new_n859_), .A2(new_n514_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n649_), .A2(new_n437_), .A3(new_n556_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n911_), .A2(new_n615_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(G169gat), .ZN(new_n914_));
  OR2_X1    g713(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n915_));
  NAND2_X1  g714(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n913_), .A2(KEYINPUT123), .A3(KEYINPUT62), .A4(G169gat), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n911_), .A2(new_n912_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n615_), .A2(new_n372_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT124), .ZN(new_n921_));
  OAI211_X1 g720(.A(new_n917_), .B(new_n918_), .C1(new_n919_), .C2(new_n921_), .ZN(G1348gat));
  OR2_X1    g721(.A1(new_n911_), .A2(KEYINPUT125), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n911_), .A2(KEYINPUT125), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n645_), .A2(new_n353_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n923_), .A2(new_n912_), .A3(new_n924_), .A4(new_n925_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n353_), .B1(new_n919_), .B2(new_n746_), .ZN(new_n927_));
  AND2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1349gat));
  AND2_X1   g727(.A1(new_n342_), .A2(new_n344_), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n919_), .A2(new_n929_), .A3(new_n250_), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n923_), .A2(new_n817_), .A3(new_n912_), .A4(new_n924_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n931_), .B2(new_n343_), .ZN(G1350gat));
  OAI21_X1  g731(.A(G190gat), .B1(new_n919_), .B2(new_n692_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n658_), .B1(new_n346_), .B2(new_n345_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n919_), .B2(new_n934_), .ZN(G1351gat));
  NAND4_X1  g734(.A1(new_n438_), .A2(new_n556_), .A3(new_n514_), .A4(new_n584_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n859_), .A2(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n615_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n644_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n322_), .A2(KEYINPUT126), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n940_), .B(new_n941_), .ZN(G1353gat));
  NAND2_X1  g741(.A1(new_n937_), .A2(new_n817_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n944_));
  AND2_X1   g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n943_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n946_), .B1(new_n943_), .B2(new_n944_), .ZN(G1354gat));
  NAND3_X1  g746(.A1(new_n937_), .A2(G218gat), .A3(new_n309_), .ZN(new_n948_));
  NOR3_X1   g747(.A1(new_n859_), .A2(new_n845_), .A3(new_n936_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n949_), .B2(G218gat), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n950_), .B(new_n951_), .ZN(G1355gat));
endmodule


