//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n780_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n816_, new_n817_, new_n818_, new_n819_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n925_, new_n926_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n934_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n967_, new_n968_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n976_,
    new_n977_, new_n978_;
  INV_X1    g000(.A(KEYINPUT74), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT36), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G190gat), .B(G218gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(G134gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G162gat), .ZN(new_n206_));
  INV_X1    g005(.A(G134gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n204_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G162gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n203_), .B1(new_n206_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n206_), .A2(new_n210_), .A3(new_n203_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n202_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n213_), .ZN(new_n215_));
  NOR3_X1   g014(.A1(new_n215_), .A2(new_n211_), .A3(KEYINPUT74), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G232gat), .A2(G233gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT34), .ZN(new_n219_));
  AND3_X1   g018(.A1(new_n219_), .A2(KEYINPUT70), .A3(KEYINPUT35), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT70), .B1(new_n219_), .B2(KEYINPUT35), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT72), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT10), .B(G99gat), .Z(new_n225_));
  INV_X1    g024(.A(G106gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n228_), .A2(KEYINPUT9), .ZN(new_n229_));
  OR2_X1    g028(.A1(G85gat), .A2(G92gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n230_), .A2(KEYINPUT9), .A3(new_n228_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G99gat), .A2(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT6), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n227_), .A2(new_n229_), .A3(new_n231_), .A4(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT7), .ZN(new_n238_));
  INV_X1    g037(.A(G99gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n238_), .A2(new_n239_), .A3(new_n226_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n240_), .A2(new_n234_), .A3(new_n235_), .A4(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT8), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n230_), .A2(new_n228_), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n242_), .B2(new_n244_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n237_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(KEYINPUT65), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n237_), .B(new_n249_), .C1(new_n245_), .C2(new_n246_), .ZN(new_n250_));
  INV_X1    g049(.A(G50gat), .ZN(new_n251_));
  OR2_X1    g050(.A1(G29gat), .A2(G36gat), .ZN(new_n252_));
  INV_X1    g051(.A(G43gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G29gat), .A2(G36gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n253_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n251_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n257_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(G50gat), .A3(new_n255_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n258_), .A2(new_n260_), .A3(KEYINPUT15), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n260_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT15), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n248_), .A2(new_n250_), .B1(new_n261_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT34), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n218_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT35), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n223_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n271_), .B(new_n272_), .C1(new_n247_), .C2(new_n262_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n224_), .B1(new_n265_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n264_), .A2(new_n261_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n246_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n249_), .B1(new_n278_), .B2(new_n237_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n250_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n275_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n224_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n273_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n217_), .A2(new_n274_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT75), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT75), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n217_), .A2(new_n274_), .A3(new_n284_), .A4(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n274_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT73), .B1(new_n289_), .B2(new_n215_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n291_));
  AOI211_X1 g090(.A(new_n291_), .B(new_n213_), .C1(new_n284_), .C2(new_n274_), .ZN(new_n292_));
  OAI211_X1 g091(.A(new_n286_), .B(new_n288_), .C1(new_n290_), .C2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT76), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT37), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n293_), .B2(KEYINPUT37), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n290_), .A2(new_n292_), .ZN(new_n297_));
  NOR3_X1   g096(.A1(new_n289_), .A2(new_n215_), .A3(new_n211_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n297_), .A2(KEYINPUT37), .A3(new_n298_), .ZN(new_n299_));
  NOR3_X1   g098(.A1(new_n295_), .A2(new_n296_), .A3(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT16), .B(G183gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(G211gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G127gat), .B(G155gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(G8gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(KEYINPUT77), .B(G1gat), .Z(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT14), .B1(new_n306_), .B2(new_n305_), .ZN(new_n307_));
  INV_X1    g106(.A(G1gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G15gat), .B(G22gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n308_), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n308_), .B1(new_n307_), .B2(new_n309_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n305_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n312_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(G8gat), .A3(new_n310_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G57gat), .B(G64gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT11), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G71gat), .B(G78gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(G57gat), .ZN(new_n321_));
  INV_X1    g120(.A(G64gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT11), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G57gat), .A2(G64gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n318_), .A2(new_n320_), .A3(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n317_), .A2(new_n319_), .A3(KEYINPUT11), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G231gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n316_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT78), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n304_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT17), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n335_), .A2(new_n336_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n333_), .A2(new_n304_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n300_), .A2(new_n340_), .ZN(new_n341_));
  XOR2_X1   g140(.A(new_n341_), .B(KEYINPUT79), .Z(new_n342_));
  INV_X1    g141(.A(new_n329_), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n343_), .A2(KEYINPUT12), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n345_));
  AOI21_X1  g144(.A(KEYINPUT12), .B1(new_n247_), .B2(new_n343_), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n329_), .B(new_n237_), .C1(new_n246_), .C2(new_n245_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n346_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G230gat), .A2(G233gat), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n345_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G120gat), .B(G148gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT66), .B(KEYINPUT5), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G176gat), .B(G204gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n247_), .A2(new_n343_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(KEYINPUT64), .A3(new_n347_), .ZN(new_n358_));
  OR3_X1    g157(.A1(new_n247_), .A2(new_n343_), .A3(KEYINPUT64), .ZN(new_n359_));
  INV_X1    g158(.A(new_n350_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n351_), .A2(new_n356_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT68), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n351_), .A2(KEYINPUT68), .A3(new_n356_), .A4(new_n361_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n356_), .B(KEYINPUT67), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n367_), .B1(new_n351_), .B2(new_n361_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n366_), .A2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT69), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT13), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n366_), .A2(KEYINPUT69), .A3(new_n369_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n372_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(KEYINPUT69), .B1(new_n366_), .B2(new_n369_), .ZN(new_n376_));
  AOI211_X1 g175(.A(new_n371_), .B(new_n368_), .C1(new_n364_), .C2(new_n365_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT13), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G127gat), .B(G134gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G113gat), .A2(G120gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G113gat), .A2(G120gat), .ZN(new_n385_));
  NOR3_X1   g184(.A1(new_n384_), .A2(new_n385_), .A3(KEYINPUT85), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n387_));
  OR2_X1    g186(.A1(G113gat), .A2(G120gat), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(new_n383_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n382_), .B1(new_n386_), .B2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT85), .B1(new_n384_), .B2(new_n385_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n388_), .A2(new_n387_), .A3(new_n383_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n381_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT31), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT83), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(G15gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G71gat), .B(G99gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(G43gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n399_), .B(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G169gat), .A2(G176gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT22), .B(G169gat), .ZN(new_n405_));
  INV_X1    g204(.A(G176gat), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n404_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G183gat), .A2(G190gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT23), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT23), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(G183gat), .A3(G190gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  OR2_X1    g211(.A1(G183gat), .A2(G190gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n407_), .A2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(G169gat), .A2(G176gat), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT24), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(G169gat), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n406_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(KEYINPUT24), .A3(new_n403_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(KEYINPUT81), .A2(G183gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT25), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT25), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(KEYINPUT81), .A3(G183gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n427_));
  NOR2_X1   g226(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n418_), .B(new_n421_), .C1(new_n426_), .C2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT82), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n411_), .A2(new_n431_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n410_), .A2(KEYINPUT82), .A3(G183gat), .A4(G190gat), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n432_), .A2(new_n409_), .A3(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n415_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n435_), .A2(KEYINPUT30), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT30), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n426_), .A2(new_n429_), .ZN(new_n438_));
  AND2_X1   g237(.A1(new_n421_), .A2(new_n418_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n432_), .A2(new_n409_), .A3(new_n433_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n437_), .B1(new_n441_), .B2(new_n415_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n436_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n402_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n443_), .A2(new_n444_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT84), .B1(new_n436_), .B2(new_n442_), .ZN(new_n448_));
  AND2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n402_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n396_), .B(new_n446_), .C1(new_n449_), .C2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n395_), .B1(new_n452_), .B2(new_n445_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT0), .B(G57gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(G85gat), .ZN(new_n456_));
  XOR2_X1   g255(.A(G1gat), .B(G29gat), .Z(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(new_n457_), .Z(new_n458_));
  INV_X1    g257(.A(G141gat), .ZN(new_n459_));
  INV_X1    g258(.A(G148gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n461_));
  OAI211_X1 g260(.A(new_n459_), .B(new_n460_), .C1(new_n461_), .C2(KEYINPUT3), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT3), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n463_), .B(KEYINPUT87), .C1(G141gat), .C2(G148gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G141gat), .A2(G148gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT86), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT86), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(G141gat), .A3(G148gat), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT2), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n465_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G155gat), .A2(G162gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G155gat), .A2(G162gat), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n473_), .A2(new_n478_), .ZN(new_n479_));
  NOR3_X1   g278(.A1(new_n475_), .A2(new_n476_), .A3(KEYINPUT1), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n467_), .A2(new_n469_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT1), .ZN(new_n482_));
  OAI22_X1  g281(.A1(new_n474_), .A2(new_n482_), .B1(G141gat), .B2(G148gat), .ZN(new_n483_));
  OR3_X1    g282(.A1(new_n480_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n394_), .A2(new_n479_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n472_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n486_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n477_), .B1(new_n487_), .B2(new_n471_), .ZN(new_n488_));
  NOR3_X1   g287(.A1(new_n480_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n393_), .B(new_n390_), .C1(new_n488_), .C2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n485_), .A2(new_n490_), .A3(KEYINPUT4), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n479_), .A2(new_n484_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT4), .ZN(new_n493_));
  NAND4_X1  g292(.A1(new_n492_), .A2(new_n493_), .A3(new_n393_), .A4(new_n390_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n491_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G225gat), .A2(G233gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n497_), .B1(new_n485_), .B2(new_n490_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n458_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n496_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n458_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(new_n502_), .A2(new_n503_), .A3(new_n499_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n501_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT27), .ZN(new_n506_));
  XOR2_X1   g305(.A(G197gat), .B(G204gat), .Z(new_n507_));
  OR2_X1    g306(.A1(G211gat), .A2(G218gat), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT21), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G211gat), .A2(G218gat), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n508_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(G211gat), .A2(G218gat), .ZN(new_n512_));
  NOR2_X1   g311(.A1(G211gat), .A2(G218gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT21), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n507_), .A2(new_n511_), .A3(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G197gat), .B(G204gat), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n516_), .B(KEYINPUT21), .C1(new_n513_), .C2(new_n512_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n417_), .A2(KEYINPUT92), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT92), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT24), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n416_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n420_), .A2(new_n519_), .A3(new_n521_), .A4(new_n403_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n412_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(G183gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT25), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n424_), .A2(G183gat), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OR2_X1    g328(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(KEYINPUT91), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT91), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n529_), .B1(new_n532_), .B2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n525_), .A2(new_n535_), .ZN(new_n536_));
  AND2_X1   g335(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n406_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(new_n403_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n540_), .B1(new_n440_), .B2(new_n413_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n518_), .B1(new_n536_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n518_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(new_n441_), .A3(new_n415_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G226gat), .A2(G233gat), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n545_), .B(KEYINPUT90), .Z(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT19), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n542_), .A2(new_n544_), .A3(KEYINPUT20), .A4(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT20), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n435_), .B2(new_n518_), .ZN(new_n551_));
  AOI22_X1  g350(.A1(new_n522_), .A2(new_n416_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n552_));
  NOR3_X1   g351(.A1(new_n427_), .A2(new_n428_), .A3(new_n533_), .ZN(new_n553_));
  AOI21_X1  g352(.A(KEYINPUT91), .B1(new_n530_), .B2(new_n531_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n552_), .B(new_n524_), .C1(new_n555_), .C2(new_n529_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n440_), .A2(new_n413_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(new_n407_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n543_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n547_), .B1(new_n551_), .B2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G8gat), .B(G36gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G64gat), .B(G92gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  NOR3_X1   g364(.A1(new_n549_), .A2(new_n560_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n565_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n551_), .A2(new_n559_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n547_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n567_), .B1(new_n570_), .B2(new_n548_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n506_), .B1(new_n566_), .B2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n565_), .B1(new_n549_), .B2(new_n560_), .ZN(new_n573_));
  AND4_X1   g372(.A1(KEYINPUT20), .A2(new_n542_), .A3(new_n569_), .A4(new_n544_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n515_), .A2(new_n517_), .A3(KEYINPUT88), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT88), .B1(new_n515_), .B2(new_n517_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n556_), .B(new_n558_), .C1(new_n575_), .C2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(KEYINPUT95), .B(KEYINPUT20), .Z(new_n578_));
  AOI21_X1  g377(.A(new_n578_), .B1(new_n435_), .B2(new_n518_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n569_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n567_), .B1(new_n574_), .B2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n573_), .A2(new_n581_), .A3(KEYINPUT27), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n505_), .A2(new_n572_), .A3(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G78gat), .B(G106gat), .Z(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(G228gat), .ZN(new_n586_));
  INV_X1    g385(.A(G233gat), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n492_), .A2(KEYINPUT29), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n575_), .A2(new_n576_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n589_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT29), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n593_), .B1(new_n479_), .B2(new_n484_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n518_), .A2(new_n589_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n585_), .B1(new_n592_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT88), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n518_), .A2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n515_), .A2(new_n517_), .A3(KEYINPUT88), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n588_), .B1(new_n601_), .B2(new_n594_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n602_), .B(new_n584_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT89), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n488_), .A2(new_n489_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G22gat), .B(G50gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT28), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n605_), .A2(new_n593_), .A3(new_n607_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n605_), .B2(new_n593_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND4_X1  g410(.A1(new_n597_), .A2(new_n603_), .A3(new_n604_), .A4(new_n611_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n610_), .B(new_n585_), .C1(new_n592_), .C2(new_n596_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n592_), .A2(new_n596_), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n614_), .B(new_n584_), .C1(KEYINPUT89), .C2(new_n610_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n612_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n454_), .B1(new_n583_), .B2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n498_), .A2(new_n458_), .A3(new_n500_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n503_), .B1(new_n502_), .B2(new_n499_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n565_), .A2(KEYINPUT32), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(new_n549_), .B2(new_n560_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n621_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n623_), .B1(new_n574_), .B2(new_n580_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT96), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT96), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n626_), .B(new_n623_), .C1(new_n574_), .C2(new_n580_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n620_), .A2(new_n622_), .A3(new_n625_), .A4(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n612_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT94), .B1(new_n495_), .B2(new_n497_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n485_), .A2(new_n490_), .A3(new_n497_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT94), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n491_), .A2(new_n632_), .A3(new_n496_), .A4(new_n494_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n630_), .A2(new_n631_), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n503_), .B1(new_n634_), .B2(KEYINPUT33), .ZN(new_n635_));
  OR3_X1    g434(.A1(new_n502_), .A2(KEYINPUT33), .A3(new_n499_), .ZN(new_n636_));
  OAI211_X1 g435(.A(KEYINPUT33), .B(new_n503_), .C1(new_n502_), .C2(new_n499_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n570_), .A2(new_n548_), .A3(new_n567_), .ZN(new_n638_));
  NAND4_X1  g437(.A1(new_n636_), .A2(new_n637_), .A3(new_n573_), .A4(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n628_), .B(new_n629_), .C1(new_n635_), .C2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n617_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n641_), .A2(KEYINPUT97), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT97), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n617_), .A2(new_n640_), .A3(new_n643_), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n629_), .A2(new_n505_), .A3(new_n572_), .A4(new_n582_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n454_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT98), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n572_), .A2(new_n582_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(new_n616_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT98), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n649_), .A2(new_n650_), .A3(new_n505_), .A4(new_n454_), .ZN(new_n651_));
  AOI22_X1  g450(.A1(new_n642_), .A2(new_n644_), .B1(new_n647_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT80), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n262_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(G229gat), .A2(G233gat), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n275_), .A2(new_n315_), .A3(new_n313_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n656_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n313_), .A2(new_n315_), .A3(new_n262_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n659_), .B1(new_n660_), .B2(new_n654_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(G113gat), .B(G141gat), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(new_n419_), .ZN(new_n663_));
  INV_X1    g462(.A(G197gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n658_), .A2(new_n661_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(new_n658_), .B2(new_n661_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n653_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n669_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n671_), .A2(KEYINPUT80), .A3(new_n667_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT99), .B1(new_n652_), .B2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n651_), .A2(new_n647_), .ZN(new_n676_));
  AND3_X1   g475(.A1(new_n617_), .A2(new_n640_), .A3(new_n643_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n643_), .B1(new_n617_), .B2(new_n640_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n676_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n679_), .A2(new_n680_), .A3(new_n673_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n380_), .B1(new_n675_), .B2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n342_), .A2(new_n683_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT100), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n620_), .A3(new_n306_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n379_), .B2(new_n673_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n379_), .A2(new_n689_), .A3(new_n673_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n297_), .A2(new_n298_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n340_), .A2(new_n693_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n691_), .A2(new_n679_), .A3(new_n692_), .A4(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(G1gat), .B1(new_n695_), .B2(new_n505_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n686_), .A2(new_n687_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n688_), .A2(new_n696_), .A3(new_n697_), .ZN(G1324gat));
  NAND3_X1  g497(.A1(new_n685_), .A2(new_n305_), .A3(new_n648_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n648_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G8gat), .B1(new_n695_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT103), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT39), .B1(new_n701_), .B2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n702_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n699_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT40), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n699_), .A2(new_n705_), .A3(KEYINPUT40), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1325gat));
  INV_X1    g509(.A(new_n684_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n711_), .A2(G15gat), .A3(new_n646_), .ZN(new_n712_));
  OAI21_X1  g511(.A(G15gat), .B1(new_n695_), .B2(new_n646_), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n713_), .B(KEYINPUT41), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1326gat));
  OAI21_X1  g514(.A(G22gat), .B1(new_n695_), .B2(new_n629_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT42), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n629_), .A2(G22gat), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT104), .Z(new_n719_));
  OAI21_X1  g518(.A(new_n717_), .B1(new_n711_), .B2(new_n719_), .ZN(G1327gat));
  NAND2_X1  g519(.A1(new_n340_), .A2(new_n693_), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n380_), .B(new_n721_), .C1(new_n675_), .C2(new_n681_), .ZN(new_n722_));
  AOI21_X1  g521(.A(G29gat), .B1(new_n722_), .B2(new_n620_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n293_), .A2(KEYINPUT37), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT76), .ZN(new_n725_));
  INV_X1    g524(.A(new_n299_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n293_), .A2(new_n294_), .A3(KEYINPUT37), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n725_), .A2(new_n726_), .A3(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(KEYINPUT43), .B1(new_n652_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n679_), .A2(new_n300_), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  AOI211_X1 g531(.A(KEYINPUT102), .B(new_n674_), .C1(new_n375_), .C2(new_n378_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n340_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n690_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n732_), .A2(new_n735_), .A3(KEYINPUT44), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT105), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT105), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n732_), .A2(new_n735_), .A3(new_n738_), .A4(KEYINPUT44), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT44), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n679_), .A2(new_n730_), .A3(new_n300_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n730_), .B1(new_n679_), .B2(new_n300_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n691_), .A2(new_n692_), .A3(new_n340_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n740_), .A2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(new_n505_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n723_), .B1(new_n748_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g548(.A(G36gat), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n732_), .A2(new_n735_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n700_), .B1(new_n751_), .B2(new_n741_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n750_), .B1(new_n740_), .B2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n721_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n682_), .A2(new_n750_), .A3(new_n648_), .A4(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT45), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT45), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n722_), .A2(new_n757_), .A3(new_n750_), .A4(new_n648_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT106), .B1(new_n753_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n756_), .A2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n746_), .A2(new_n648_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n737_), .B2(new_n739_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n761_), .B(new_n762_), .C1(new_n764_), .C2(new_n750_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT46), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n760_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT107), .ZN(new_n768_));
  OAI211_X1 g567(.A(KEYINPUT46), .B(new_n762_), .C1(new_n764_), .C2(new_n750_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT107), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n760_), .A2(new_n765_), .A3(new_n770_), .A4(new_n766_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(new_n769_), .A3(new_n771_), .ZN(G1329gat));
  NAND2_X1  g571(.A1(new_n454_), .A2(G43gat), .ZN(new_n773_));
  INV_X1    g572(.A(new_n722_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n774_), .A2(new_n646_), .ZN(new_n775_));
  OAI22_X1  g574(.A1(new_n747_), .A2(new_n773_), .B1(G43gat), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g576(.A(G50gat), .B1(new_n747_), .B2(new_n629_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n616_), .A2(new_n251_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT108), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n778_), .B1(new_n774_), .B2(new_n780_), .ZN(G1331gat));
  NOR2_X1   g580(.A1(new_n379_), .A2(new_n673_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n679_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(new_n694_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n785_), .A2(new_n321_), .A3(new_n505_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n342_), .A2(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n620_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n786_), .B1(new_n788_), .B2(new_n321_), .ZN(G1332gat));
  OAI21_X1  g588(.A(G64gat), .B1(new_n785_), .B2(new_n700_), .ZN(new_n790_));
  XNOR2_X1  g589(.A(new_n790_), .B(KEYINPUT48), .ZN(new_n791_));
  INV_X1    g590(.A(new_n787_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n648_), .A2(new_n322_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT109), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n791_), .B1(new_n792_), .B2(new_n794_), .ZN(G1333gat));
  OR3_X1    g594(.A1(new_n792_), .A2(G71gat), .A3(new_n646_), .ZN(new_n796_));
  OAI21_X1  g595(.A(G71gat), .B1(new_n785_), .B2(new_n646_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n797_), .A2(KEYINPUT110), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n797_), .A2(KEYINPUT110), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n799_), .A2(KEYINPUT49), .A3(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT49), .B1(new_n799_), .B2(new_n800_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n796_), .B1(new_n801_), .B2(new_n802_), .ZN(G1334gat));
  OAI21_X1  g602(.A(G78gat), .B1(new_n785_), .B2(new_n629_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n804_), .B(KEYINPUT50), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n629_), .A2(G78gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n792_), .B2(new_n806_), .ZN(G1335gat));
  NAND3_X1  g606(.A1(new_n784_), .A2(KEYINPUT111), .A3(new_n754_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT111), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n783_), .B2(new_n721_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(G85gat), .B1(new_n811_), .B2(new_n620_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n732_), .A2(new_n782_), .A3(new_n340_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n505_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n812_), .B1(G85gat), .B2(new_n814_), .ZN(G1336gat));
  AOI21_X1  g614(.A(G92gat), .B1(new_n811_), .B2(new_n648_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n648_), .A2(G92gat), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT112), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n816_), .B1(new_n817_), .B2(new_n819_), .ZN(G1337gat));
  OAI21_X1  g619(.A(G99gat), .B1(new_n813_), .B2(new_n646_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT113), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n811_), .A2(new_n454_), .A3(new_n225_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n824_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g624(.A(G106gat), .B1(new_n813_), .B2(new_n629_), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n826_), .B(KEYINPUT52), .Z(new_n827_));
  AOI21_X1  g626(.A(G106gat), .B1(new_n808_), .B2(new_n810_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n616_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n829_), .B(KEYINPUT114), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n827_), .A2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(G1339gat));
  NAND3_X1  g632(.A1(new_n649_), .A2(new_n620_), .A3(new_n454_), .ZN(new_n834_));
  XOR2_X1   g633(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n351_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(KEYINPUT55), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n345_), .A2(new_n349_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n360_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT55), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n351_), .A2(new_n837_), .A3(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n839_), .A2(new_n841_), .A3(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n367_), .ZN(new_n845_));
  AOI21_X1  g644(.A(KEYINPUT56), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(KEYINPUT56), .A3(new_n845_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n655_), .A2(new_n659_), .A3(new_n657_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n656_), .B1(new_n660_), .B2(new_n654_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n665_), .A3(new_n851_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n667_), .A2(new_n852_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n853_), .A2(new_n366_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n836_), .B1(new_n849_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(KEYINPUT118), .B1(new_n855_), .B2(new_n728_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857_));
  INV_X1    g656(.A(new_n848_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n854_), .B1(new_n858_), .B2(new_n846_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n835_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n300_), .A2(new_n857_), .A3(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n849_), .A2(KEYINPUT58), .A3(new_n854_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n856_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT119), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT119), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n856_), .A2(new_n861_), .A3(new_n865_), .A4(new_n862_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n673_), .B(new_n366_), .C1(new_n858_), .C2(new_n846_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n853_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n693_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT120), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n869_), .A2(new_n870_), .A3(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n871_), .A2(new_n872_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n875_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n869_), .A2(new_n870_), .A3(new_n877_), .A4(new_n873_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n876_), .A2(new_n878_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n864_), .A2(new_n866_), .A3(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n340_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n882_));
  NAND4_X1  g681(.A1(new_n728_), .A2(new_n379_), .A3(new_n674_), .A4(new_n734_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n883_), .A2(KEYINPUT115), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(KEYINPUT115), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n882_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n883_), .A2(KEYINPUT115), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n883_), .A2(KEYINPUT115), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n887_), .A2(KEYINPUT54), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n886_), .A2(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n834_), .B1(new_n881_), .B2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(G113gat), .B1(new_n891_), .B2(new_n673_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n886_), .A2(new_n889_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n734_), .B1(new_n879_), .B2(new_n863_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n834_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n895_), .A2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n900_), .B1(new_n891_), .B2(new_n897_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n880_), .A2(new_n340_), .B1(new_n886_), .B2(new_n889_), .ZN(new_n902_));
  OAI211_X1 g701(.A(KEYINPUT121), .B(KEYINPUT59), .C1(new_n902_), .C2(new_n834_), .ZN(new_n903_));
  AOI211_X1 g702(.A(new_n674_), .B(new_n899_), .C1(new_n901_), .C2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n892_), .B1(new_n904_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g704(.A(G120gat), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n906_), .B1(new_n379_), .B2(KEYINPUT60), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n891_), .B(new_n907_), .C1(KEYINPUT60), .C2(new_n906_), .ZN(new_n908_));
  AOI211_X1 g707(.A(new_n379_), .B(new_n899_), .C1(new_n901_), .C2(new_n903_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n906_), .ZN(G1341gat));
  AOI21_X1  g709(.A(G127gat), .B1(new_n891_), .B2(new_n734_), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n340_), .B(new_n899_), .C1(new_n901_), .C2(new_n903_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n911_), .B1(new_n912_), .B2(G127gat), .ZN(G1342gat));
  AOI22_X1  g712(.A1(new_n863_), .A2(KEYINPUT119), .B1(new_n876_), .B2(new_n878_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n734_), .B1(new_n914_), .B2(new_n866_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n693_), .B(new_n896_), .C1(new_n893_), .C2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(new_n207_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT122), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n916_), .A2(KEYINPUT122), .A3(new_n207_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n920_), .ZN(new_n921_));
  XOR2_X1   g720(.A(KEYINPUT123), .B(G134gat), .Z(new_n922_));
  AOI211_X1 g721(.A(new_n922_), .B(new_n899_), .C1(new_n901_), .C2(new_n903_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n923_), .B2(new_n300_), .ZN(G1343gat));
  NOR3_X1   g723(.A1(new_n902_), .A2(new_n629_), .A3(new_n454_), .ZN(new_n925_));
  NAND4_X1  g724(.A1(new_n925_), .A2(new_n620_), .A3(new_n700_), .A4(new_n673_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g726(.A1(new_n925_), .A2(new_n620_), .A3(new_n700_), .A4(new_n380_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g728(.A1(new_n925_), .A2(new_n620_), .A3(new_n700_), .A4(new_n734_), .ZN(new_n930_));
  XOR2_X1   g729(.A(KEYINPUT61), .B(G155gat), .Z(new_n931_));
  XNOR2_X1  g730(.A(new_n931_), .B(KEYINPUT124), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n930_), .B(new_n932_), .ZN(G1346gat));
  AND4_X1   g732(.A1(G162gat), .A2(new_n925_), .A3(new_n620_), .A4(new_n700_), .ZN(new_n934_));
  NAND4_X1  g733(.A1(new_n925_), .A2(new_n620_), .A3(new_n700_), .A4(new_n693_), .ZN(new_n935_));
  AOI22_X1  g734(.A1(new_n934_), .A2(new_n300_), .B1(new_n209_), .B2(new_n935_), .ZN(G1347gat));
  NOR2_X1   g735(.A1(new_n700_), .A2(new_n620_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n454_), .ZN(new_n938_));
  NOR3_X1   g737(.A1(new_n895_), .A2(new_n616_), .A3(new_n938_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n939_), .A2(new_n405_), .A3(new_n673_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n674_), .A2(new_n938_), .ZN(new_n941_));
  XOR2_X1   g740(.A(new_n941_), .B(KEYINPUT125), .Z(new_n942_));
  OAI211_X1 g741(.A(new_n629_), .B(new_n942_), .C1(new_n893_), .C2(new_n894_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n944_));
  AND3_X1   g743(.A1(new_n943_), .A2(new_n944_), .A3(G169gat), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n943_), .B2(G169gat), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n940_), .B1(new_n945_), .B2(new_n946_), .ZN(G1348gat));
  NOR3_X1   g746(.A1(new_n902_), .A2(new_n616_), .A3(new_n938_), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n948_), .A2(G176gat), .A3(new_n380_), .ZN(new_n949_));
  AND2_X1   g748(.A1(new_n949_), .A2(KEYINPUT126), .ZN(new_n950_));
  NOR2_X1   g749(.A1(new_n949_), .A2(KEYINPUT126), .ZN(new_n951_));
  AOI21_X1  g750(.A(G176gat), .B1(new_n939_), .B2(new_n380_), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n950_), .A2(new_n951_), .A3(new_n952_), .ZN(G1349gat));
  AOI21_X1  g752(.A(G183gat), .B1(new_n948_), .B2(new_n734_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n340_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n954_), .B1(new_n939_), .B2(new_n955_), .ZN(G1350gat));
  NAND2_X1  g755(.A1(new_n939_), .A2(new_n300_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(G190gat), .ZN(new_n958_));
  OAI211_X1 g757(.A(new_n939_), .B(new_n693_), .C1(new_n554_), .C2(new_n553_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n958_), .A2(new_n959_), .ZN(G1351gat));
  NAND2_X1  g759(.A1(new_n925_), .A2(new_n937_), .ZN(new_n961_));
  INV_X1    g760(.A(new_n961_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n962_), .A2(new_n664_), .A3(new_n673_), .ZN(new_n963_));
  OAI21_X1  g762(.A(G197gat), .B1(new_n961_), .B2(new_n674_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n963_), .A2(new_n964_), .ZN(G1352gat));
  AOI21_X1  g764(.A(G204gat), .B1(new_n962_), .B2(new_n380_), .ZN(new_n966_));
  INV_X1    g765(.A(G204gat), .ZN(new_n967_));
  NOR3_X1   g766(.A1(new_n961_), .A2(new_n967_), .A3(new_n379_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n966_), .A2(new_n968_), .ZN(G1353gat));
  NOR2_X1   g768(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n970_));
  XNOR2_X1  g769(.A(new_n970_), .B(KEYINPUT127), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n340_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n971_), .B1(new_n962_), .B2(new_n972_), .ZN(new_n973_));
  AND4_X1   g772(.A1(new_n925_), .A2(new_n937_), .A3(new_n972_), .A4(new_n971_), .ZN(new_n974_));
  NOR2_X1   g773(.A1(new_n973_), .A2(new_n974_), .ZN(G1354gat));
  INV_X1    g774(.A(G218gat), .ZN(new_n976_));
  NOR3_X1   g775(.A1(new_n961_), .A2(new_n976_), .A3(new_n728_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n962_), .A2(new_n693_), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n977_), .B1(new_n976_), .B2(new_n978_), .ZN(G1355gat));
endmodule


