//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n915_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n950_, new_n951_, new_n953_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_;
  NAND2_X1  g000(.A1(G232gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT34), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT74), .B1(new_n203_), .B2(KEYINPUT35), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT65), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n206_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n207_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(new_n213_), .A3(KEYINPUT65), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n211_), .A2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n220_), .A2(KEYINPUT9), .ZN(new_n221_));
  INV_X1    g020(.A(G85gat), .ZN(new_n222_));
  INV_X1    g021(.A(G92gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(KEYINPUT9), .A3(new_n220_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n215_), .A2(new_n219_), .A3(new_n221_), .A4(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227_));
  AND2_X1   g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G85gat), .A2(G92gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n227_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n224_), .A2(KEYINPUT66), .A3(new_n220_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT8), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT7), .ZN(new_n234_));
  INV_X1    g033(.A(G99gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(new_n217_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n233_), .B1(new_n215_), .B2(new_n239_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n230_), .A2(new_n231_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n236_), .B(new_n237_), .C1(new_n208_), .C2(new_n210_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n232_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n226_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G29gat), .B(G36gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G43gat), .B(G50gat), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n245_), .A2(new_n246_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n205_), .B1(new_n244_), .B2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n219_), .A2(new_n225_), .A3(new_n221_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n252_), .B1(new_n214_), .B2(new_n211_), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n212_), .A2(new_n213_), .A3(KEYINPUT65), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT65), .B1(new_n212_), .B2(new_n213_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n239_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n233_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n212_), .A2(new_n213_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n259_), .A2(new_n238_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n230_), .A2(new_n231_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT8), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n253_), .B1(new_n258_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT15), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n249_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n247_), .A2(KEYINPUT15), .A3(new_n248_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n263_), .A2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT71), .B1(new_n251_), .B2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n204_), .B1(new_n263_), .B2(new_n249_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n244_), .A2(new_n266_), .A3(new_n265_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n269_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n203_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT35), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n269_), .A2(new_n277_), .A3(new_n273_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G190gat), .B(G218gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT72), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G134gat), .B(G162gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n284_), .B(new_n285_), .Z(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n282_), .A2(KEYINPUT36), .A3(new_n287_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n269_), .A2(new_n277_), .A3(new_n273_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n277_), .B1(new_n269_), .B2(new_n273_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n286_), .B1(new_n291_), .B2(new_n280_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n279_), .A2(new_n281_), .A3(new_n286_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT36), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n288_), .B1(new_n292_), .B2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT75), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT37), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n282_), .A2(new_n287_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(new_n294_), .A3(new_n293_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(KEYINPUT75), .A2(KEYINPUT37), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n298_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n288_), .A4(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n299_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT77), .ZN(new_n306_));
  INV_X1    g105(.A(G1gat), .ZN(new_n307_));
  INV_X1    g106(.A(G8gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT14), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT76), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT76), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n311_), .B(KEYINPUT14), .C1(new_n307_), .C2(new_n308_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G15gat), .B(G22gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G1gat), .B(G8gat), .Z(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n310_), .A2(new_n315_), .A3(new_n312_), .A4(new_n313_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n319_), .A2(G231gat), .A3(G233gat), .ZN(new_n320_));
  INV_X1    g119(.A(G231gat), .ZN(new_n321_));
  INV_X1    g120(.A(G233gat), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n317_), .B(new_n318_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G71gat), .B(G78gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G57gat), .B(G64gat), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n324_), .B1(KEYINPUT11), .B2(new_n325_), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n325_), .A2(KEYINPUT11), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n325_), .A2(new_n324_), .A3(KEYINPUT11), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n320_), .A2(new_n323_), .A3(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n331_), .B1(new_n320_), .B2(new_n323_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n306_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n334_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n336_), .A2(KEYINPUT77), .A3(new_n332_), .ZN(new_n337_));
  XOR2_X1   g136(.A(G127gat), .B(G155gat), .Z(new_n338_));
  XNOR2_X1  g137(.A(new_n338_), .B(KEYINPUT16), .ZN(new_n339_));
  XNOR2_X1  g138(.A(G183gat), .B(G211gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT17), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n335_), .A2(new_n337_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n336_), .A2(KEYINPUT78), .A3(new_n332_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n341_), .B(KEYINPUT17), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n344_), .A2(new_n349_), .ZN(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT12), .B1(new_n263_), .B2(new_n330_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT12), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n244_), .A2(new_n352_), .A3(new_n331_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n330_), .B(new_n226_), .C1(new_n240_), .C2(new_n243_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G230gat), .A2(G233gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n356_), .B(KEYINPUT64), .Z(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n355_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT68), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n355_), .A2(KEYINPUT68), .A3(new_n358_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n354_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n244_), .A2(new_n331_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(KEYINPUT67), .A3(new_n355_), .ZN(new_n365_));
  OR3_X1    g164(.A1(new_n263_), .A2(KEYINPUT67), .A3(new_n330_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(new_n357_), .ZN(new_n367_));
  XOR2_X1   g166(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT70), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G120gat), .B(G148gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G176gat), .B(G204gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  AND3_X1   g172(.A1(new_n363_), .A2(new_n367_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n373_), .B1(new_n363_), .B2(new_n367_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT13), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT13), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n378_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n305_), .A2(new_n350_), .A3(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT79), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT88), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G113gat), .B(G120gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT87), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G127gat), .B(G134gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n388_), .ZN(new_n390_));
  OR2_X1    g189(.A1(new_n385_), .A2(new_n386_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n385_), .A2(new_n386_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n390_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n384_), .B1(new_n389_), .B2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n385_), .B(KEYINPUT87), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n384_), .B1(new_n395_), .B2(new_n390_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT31), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT89), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G71gat), .B(G99gat), .ZN(new_n401_));
  INV_X1    g200(.A(G43gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT30), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G183gat), .A2(G190gat), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT23), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(KEYINPUT85), .ZN(new_n408_));
  OR3_X1    g207(.A1(new_n405_), .A2(KEYINPUT85), .A3(KEYINPUT23), .ZN(new_n409_));
  XOR2_X1   g208(.A(KEYINPUT82), .B(G183gat), .Z(new_n410_));
  INV_X1    g209(.A(G190gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n408_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT86), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT86), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n408_), .A2(new_n415_), .A3(new_n409_), .A4(new_n412_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G169gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n414_), .A2(new_n416_), .A3(new_n418_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n420_));
  INV_X1    g219(.A(G169gat), .ZN(new_n421_));
  INV_X1    g220(.A(G176gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT24), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n423_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n424_));
  AOI211_X1 g223(.A(new_n420_), .B(new_n407_), .C1(new_n424_), .C2(KEYINPUT84), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT25), .ZN(new_n426_));
  INV_X1    g225(.A(G183gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n428_), .B1(new_n410_), .B2(new_n426_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT26), .ZN(new_n430_));
  OR3_X1    g229(.A1(new_n430_), .A2(KEYINPUT83), .A3(G190gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(G190gat), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT83), .B1(new_n430_), .B2(G190gat), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n429_), .A2(new_n431_), .A3(new_n432_), .A4(new_n433_), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n424_), .A2(KEYINPUT84), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n425_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n404_), .B1(new_n419_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n419_), .A2(new_n436_), .A3(new_n404_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G227gat), .A2(G233gat), .ZN(new_n441_));
  INV_X1    g240(.A(G15gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n400_), .B1(new_n440_), .B2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n438_), .A2(new_n443_), .A3(new_n439_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n399_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n439_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n444_), .B1(new_n448_), .B2(new_n437_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n446_), .A3(KEYINPUT89), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(KEYINPUT31), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n398_), .B1(new_n447_), .B2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n445_), .A2(new_n399_), .A3(new_n446_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n450_), .A2(KEYINPUT31), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n387_), .A2(new_n388_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n395_), .A2(new_n390_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n396_), .B1(new_n457_), .B2(new_n384_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(new_n454_), .A3(new_n458_), .ZN(new_n459_));
  AND2_X1   g258(.A1(new_n452_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G211gat), .B(G218gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT94), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G197gat), .B(G204gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n463_), .B(KEYINPUT21), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n463_), .A2(KEYINPUT96), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(KEYINPUT96), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n466_), .A2(KEYINPUT21), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n462_), .ZN(new_n469_));
  AOI22_X1  g268(.A1(new_n465_), .A2(KEYINPUT95), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT95), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n462_), .A2(new_n464_), .A3(new_n471_), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n470_), .A2(new_n419_), .A3(new_n472_), .A4(new_n436_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n465_), .A2(KEYINPUT95), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n468_), .A2(new_n469_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n472_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n408_), .A2(new_n409_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(KEYINPUT25), .B(G183gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT26), .B(G190gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n424_), .A2(new_n420_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n477_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT22), .B(G169gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT101), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n422_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n407_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n427_), .A2(new_n411_), .ZN(new_n488_));
  AOI22_X1  g287(.A1(new_n487_), .A2(new_n488_), .B1(G169gat), .B2(G176gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n486_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n482_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n476_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n473_), .A2(new_n492_), .A3(KEYINPUT20), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G226gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT19), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(new_n476_), .A2(new_n491_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n419_), .A2(new_n436_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n476_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n495_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n497_), .A2(KEYINPUT20), .A3(new_n499_), .A4(new_n500_), .ZN(new_n501_));
  XOR2_X1   g300(.A(G8gat), .B(G36gat), .Z(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT18), .ZN(new_n503_));
  XNOR2_X1  g302(.A(G64gat), .B(G92gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n496_), .A2(new_n501_), .A3(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT20), .B1(new_n476_), .B2(new_n491_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n472_), .A2(new_n470_), .B1(new_n419_), .B2(new_n436_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n495_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n473_), .A2(new_n492_), .A3(KEYINPUT20), .A4(new_n500_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n510_), .A2(new_n512_), .ZN(new_n513_));
  OAI211_X1 g312(.A(KEYINPUT27), .B(new_n506_), .C1(new_n513_), .C2(new_n505_), .ZN(new_n514_));
  XOR2_X1   g313(.A(KEYINPUT106), .B(KEYINPUT27), .Z(new_n515_));
  AND3_X1   g314(.A1(new_n496_), .A2(new_n505_), .A3(new_n501_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n505_), .B1(new_n496_), .B2(new_n501_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n515_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n460_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G141gat), .A2(G148gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT92), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT2), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT2), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n521_), .A2(KEYINPUT92), .A3(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(G141gat), .A2(G148gat), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT3), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n523_), .A2(new_n525_), .A3(new_n528_), .A4(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G155gat), .B(G162gat), .Z(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT93), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n530_), .A2(KEYINPUT93), .A3(new_n531_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G155gat), .A2(G162gat), .ZN(new_n536_));
  NOR2_X1   g335(.A1(G155gat), .A2(G162gat), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n536_), .B1(new_n537_), .B2(KEYINPUT1), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT90), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(KEYINPUT90), .B(new_n536_), .C1(new_n537_), .C2(KEYINPUT1), .ZN(new_n541_));
  OR3_X1    g340(.A1(new_n536_), .A2(KEYINPUT91), .A3(KEYINPUT1), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT91), .B1(new_n536_), .B2(KEYINPUT1), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n540_), .A2(new_n541_), .A3(new_n542_), .A4(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n521_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n545_), .A2(new_n526_), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n534_), .A2(new_n535_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT29), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT28), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n549_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G22gat), .B(G50gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n549_), .B(KEYINPUT28), .ZN(new_n554_));
  INV_X1    g353(.A(new_n552_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G78gat), .B(G106gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT99), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT97), .B1(new_n547_), .B2(new_n548_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n544_), .A2(new_n546_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n535_), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT93), .B1(new_n530_), .B2(new_n531_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n561_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT97), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n565_), .A3(KEYINPUT29), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(new_n566_), .A3(new_n476_), .ZN(new_n567_));
  INV_X1    g366(.A(G228gat), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n568_), .A2(new_n322_), .ZN(new_n569_));
  AOI21_X1  g368(.A(KEYINPUT98), .B1(new_n567_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n567_), .A2(KEYINPUT98), .A3(new_n569_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  OAI221_X1 g372(.A(new_n476_), .B1(new_n568_), .B2(new_n322_), .C1(new_n548_), .C2(new_n547_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n559_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n567_), .A2(KEYINPUT98), .A3(new_n569_), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n559_), .B(new_n574_), .C1(new_n576_), .C2(new_n570_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n557_), .B1(new_n575_), .B2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n574_), .B1(new_n576_), .B2(new_n570_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n557_), .B1(new_n580_), .B2(new_n558_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n573_), .A2(KEYINPUT100), .A3(new_n559_), .A4(new_n574_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT100), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n577_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n581_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n579_), .A2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G1gat), .B(G29gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT103), .B(KEYINPUT0), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G57gat), .B(G85gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n547_), .A2(new_n457_), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n593_), .B(KEYINPUT4), .C1(new_n398_), .C2(new_n547_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G225gat), .A2(G233gat), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT4), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n458_), .A2(new_n597_), .A3(new_n564_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n594_), .A2(KEYINPUT102), .A3(new_n596_), .A4(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n458_), .A2(new_n564_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(new_n593_), .A3(new_n595_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n598_), .A2(new_n596_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT102), .B1(new_n603_), .B2(new_n594_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n592_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT102), .ZN(new_n606_));
  INV_X1    g405(.A(new_n594_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n598_), .A2(new_n596_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n609_), .A2(new_n591_), .A3(new_n601_), .A4(new_n599_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n605_), .A2(new_n610_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n520_), .A2(new_n586_), .A3(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n611_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n586_), .A2(new_n613_), .A3(new_n519_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT105), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n505_), .A2(KEYINPUT32), .ZN(new_n616_));
  AOI211_X1 g415(.A(new_n615_), .B(new_n616_), .C1(new_n509_), .C2(new_n511_), .ZN(new_n617_));
  OAI211_X1 g416(.A(KEYINPUT32), .B(new_n505_), .C1(new_n510_), .C2(new_n512_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n496_), .A2(new_n501_), .A3(new_n616_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT105), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n617_), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(new_n611_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n610_), .A2(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n599_), .A2(new_n601_), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n625_), .A2(KEYINPUT33), .A3(new_n591_), .A4(new_n609_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n516_), .A2(new_n517_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n600_), .A2(new_n593_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n591_), .B1(new_n629_), .B2(new_n596_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT104), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n598_), .A2(new_n595_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n631_), .B1(new_n632_), .B2(new_n594_), .ZN(new_n633_));
  AND4_X1   g432(.A1(new_n631_), .A2(new_n594_), .A3(new_n595_), .A4(new_n598_), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n630_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n624_), .A2(new_n626_), .A3(new_n627_), .A4(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n622_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n579_), .A3(new_n585_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n614_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n460_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n612_), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n319_), .A2(new_n265_), .A3(new_n266_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n317_), .A2(new_n249_), .A3(new_n318_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(G229gat), .A2(G233gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n644_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n317_), .A2(new_n249_), .A3(new_n318_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n249_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n646_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G113gat), .B(G141gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT80), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G169gat), .B(G197gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n645_), .A2(new_n649_), .A3(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT81), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n653_), .B1(new_n645_), .B2(new_n649_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n656_), .B(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n641_), .A2(new_n658_), .ZN(new_n659_));
  AND2_X1   g458(.A1(new_n383_), .A2(new_n659_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n613_), .B(KEYINPUT107), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n660_), .A2(new_n307_), .A3(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT108), .B(KEYINPUT38), .ZN(new_n663_));
  INV_X1    g462(.A(new_n296_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n641_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n657_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n656_), .B(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n380_), .A2(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(new_n350_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n665_), .A2(new_n611_), .A3(new_n669_), .ZN(new_n670_));
  AOI22_X1  g469(.A1(new_n662_), .A2(new_n663_), .B1(G1gat), .B2(new_n670_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n662_), .A2(new_n663_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n672_), .A2(KEYINPUT109), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(KEYINPUT109), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n671_), .B1(new_n673_), .B2(new_n674_), .ZN(G1324gat));
  AOI21_X1  g474(.A(new_n460_), .B1(new_n614_), .B2(new_n638_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n296_), .B(new_n669_), .C1(new_n676_), .C2(new_n612_), .ZN(new_n677_));
  OAI21_X1  g476(.A(G8gat), .B1(new_n677_), .B2(new_n519_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n678_), .A2(KEYINPUT39), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT39), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n680_), .B(G8gat), .C1(new_n677_), .C2(new_n519_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n519_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n659_), .A2(new_n383_), .A3(new_n308_), .A4(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(KEYINPUT110), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT110), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n682_), .A2(new_n687_), .A3(new_n684_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(KEYINPUT111), .B(KEYINPUT40), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n686_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n689_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1325gat));
  NAND3_X1  g491(.A1(new_n660_), .A2(new_n442_), .A3(new_n460_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n665_), .A2(new_n460_), .A3(new_n669_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n694_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT41), .B1(new_n694_), .B2(G15gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(G1326gat));
  XOR2_X1   g497(.A(new_n586_), .B(KEYINPUT112), .Z(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G22gat), .B1(new_n677_), .B2(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT42), .ZN(new_n702_));
  INV_X1    g501(.A(G22gat), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n660_), .A2(new_n703_), .A3(new_n699_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n704_), .ZN(G1327gat));
  NAND2_X1  g504(.A1(new_n664_), .A2(new_n350_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n706_), .A2(new_n381_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n659_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G29gat), .B1(new_n709_), .B2(new_n611_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n305_), .ZN(new_n711_));
  OAI21_X1  g510(.A(KEYINPUT43), .B1(new_n641_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n713_), .B(new_n305_), .C1(new_n676_), .C2(new_n612_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n344_), .A2(new_n349_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n668_), .A2(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(KEYINPUT44), .B1(new_n715_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n719_));
  INV_X1    g518(.A(new_n717_), .ZN(new_n720_));
  AOI211_X1 g519(.A(new_n719_), .B(new_n720_), .C1(new_n712_), .C2(new_n714_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n718_), .A2(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n661_), .A2(G29gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n710_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  INV_X1    g524(.A(G36gat), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n726_), .B1(new_n722_), .B2(new_n683_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n519_), .A2(G36gat), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OR3_X1    g528(.A1(new_n708_), .A2(KEYINPUT45), .A3(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(KEYINPUT45), .B1(new_n708_), .B2(new_n729_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n725_), .B1(new_n727_), .B2(new_n733_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n718_), .A2(new_n721_), .A3(new_n519_), .ZN(new_n735_));
  OAI211_X1 g534(.A(KEYINPUT46), .B(new_n732_), .C1(new_n735_), .C2(new_n726_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1329gat));
  NOR2_X1   g536(.A1(new_n640_), .A2(new_n402_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n722_), .A2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n402_), .B1(new_n708_), .B2(new_n640_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT47), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n739_), .A2(new_n743_), .A3(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1330gat));
  OR3_X1    g544(.A1(new_n708_), .A2(G50gat), .A3(new_n700_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n722_), .A2(KEYINPUT113), .A3(new_n586_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G50gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(KEYINPUT113), .B1(new_n722_), .B2(new_n586_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n748_), .B2(new_n749_), .ZN(G1331gat));
  NOR2_X1   g549(.A1(new_n380_), .A2(new_n667_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n665_), .A2(new_n716_), .A3(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G57gat), .B1(new_n752_), .B2(new_n613_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n641_), .A2(new_n667_), .A3(new_n380_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n711_), .A3(new_n716_), .ZN(new_n755_));
  INV_X1    g554(.A(G57gat), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n661_), .A2(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n755_), .B2(new_n757_), .ZN(G1332gat));
  OAI21_X1  g557(.A(G64gat), .B1(new_n752_), .B2(new_n519_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT48), .ZN(new_n760_));
  OR2_X1    g559(.A1(new_n519_), .A2(G64gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n755_), .B2(new_n761_), .ZN(G1333gat));
  OAI21_X1  g561(.A(G71gat), .B1(new_n752_), .B2(new_n640_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n763_), .B(KEYINPUT49), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n640_), .A2(G71gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n755_), .B2(new_n765_), .ZN(G1334gat));
  OAI21_X1  g565(.A(G78gat), .B1(new_n752_), .B2(new_n700_), .ZN(new_n767_));
  XOR2_X1   g566(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(new_n769_));
  OR2_X1    g568(.A1(new_n700_), .A2(G78gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n769_), .B1(new_n755_), .B2(new_n770_), .ZN(G1335gat));
  NAND2_X1  g570(.A1(new_n751_), .A2(new_n350_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n772_), .B1(new_n712_), .B2(new_n714_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G85gat), .B1(new_n774_), .B2(new_n613_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n706_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n754_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n222_), .A3(new_n661_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n775_), .A2(new_n779_), .ZN(G1336gat));
  OAI21_X1  g579(.A(G92gat), .B1(new_n774_), .B2(new_n519_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(new_n223_), .A3(new_n683_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(G1337gat));
  OAI21_X1  g582(.A(G99gat), .B1(new_n774_), .B2(new_n640_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n460_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n777_), .B2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g586(.A1(new_n778_), .A2(new_n217_), .A3(new_n586_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n773_), .A2(new_n586_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(G106gat), .ZN(new_n791_));
  AOI211_X1 g590(.A(KEYINPUT52), .B(new_n217_), .C1(new_n773_), .C2(new_n586_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT53), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n795_), .B(new_n788_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(G1339gat));
  INV_X1    g596(.A(new_n661_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n798_), .A2(new_n586_), .A3(new_n520_), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n374_), .A2(new_n375_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n319_), .A2(new_n250_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n646_), .B1(new_n801_), .B2(new_n643_), .ZN(new_n802_));
  OAI21_X1  g601(.A(KEYINPUT119), .B1(new_n802_), .B2(new_n653_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n644_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n805_));
  INV_X1    g604(.A(new_n653_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n803_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n642_), .A2(new_n643_), .A3(new_n646_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(KEYINPUT120), .A3(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n654_), .ZN(new_n811_));
  AOI21_X1  g610(.A(KEYINPUT120), .B1(new_n808_), .B2(new_n809_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT121), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n800_), .A2(new_n813_), .A3(new_n814_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n802_), .A2(KEYINPUT119), .A3(new_n653_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n805_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n809_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n820_), .A2(new_n654_), .A3(new_n810_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT121), .B1(new_n376_), .B2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n815_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n263_), .A2(KEYINPUT12), .A3(new_n330_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n352_), .B1(new_n244_), .B2(new_n331_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n355_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  AOI22_X1  g627(.A1(new_n363_), .A2(new_n825_), .B1(new_n828_), .B2(new_n357_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n357_), .B1(new_n263_), .B2(new_n330_), .ZN(new_n830_));
  AOI22_X1  g629(.A1(new_n351_), .A2(new_n353_), .B1(new_n830_), .B2(KEYINPUT68), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT117), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(KEYINPUT55), .A4(new_n361_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n354_), .A2(new_n361_), .A3(KEYINPUT55), .A4(new_n362_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(KEYINPUT117), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n829_), .A2(new_n833_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n373_), .ZN(new_n837_));
  AND3_X1   g636(.A1(new_n836_), .A2(KEYINPUT56), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(KEYINPUT56), .B1(new_n836_), .B2(new_n837_), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n838_), .A2(new_n839_), .A3(KEYINPUT118), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n836_), .A2(new_n837_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT56), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n841_), .A2(KEYINPUT118), .A3(new_n842_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n658_), .A2(new_n374_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n824_), .B1(new_n840_), .B2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(KEYINPUT57), .A3(new_n296_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT57), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n841_), .A2(new_n842_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n836_), .A2(KEYINPUT56), .A3(new_n837_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n850_), .A2(new_n851_), .A3(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n844_), .B1(new_n839_), .B2(KEYINPUT118), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n823_), .B1(new_n853_), .B2(new_n854_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n849_), .B1(new_n855_), .B2(new_n664_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n821_), .A2(new_n374_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n857_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(KEYINPUT58), .B(new_n857_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n305_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n848_), .A2(new_n856_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(new_n350_), .ZN(new_n864_));
  OAI21_X1  g663(.A(KEYINPUT115), .B1(new_n667_), .B2(new_n350_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT115), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n716_), .A2(new_n866_), .A3(new_n658_), .ZN(new_n867_));
  AND4_X1   g666(.A1(new_n379_), .A2(new_n865_), .A3(new_n377_), .A4(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n299_), .A2(new_n868_), .A3(new_n304_), .ZN(new_n869_));
  XOR2_X1   g668(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n869_), .A2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n299_), .A2(new_n868_), .A3(new_n304_), .A4(new_n870_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(KEYINPUT122), .B1(new_n864_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877_));
  AOI211_X1 g676(.A(new_n877_), .B(new_n874_), .C1(new_n863_), .C2(new_n350_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n799_), .B1(new_n876_), .B2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(G113gat), .B1(new_n880_), .B2(new_n667_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n874_), .B1(new_n863_), .B2(new_n350_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT59), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n799_), .A2(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n884_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n879_), .B2(KEYINPUT59), .ZN(new_n886_));
  INV_X1    g685(.A(G113gat), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n658_), .A2(new_n887_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT123), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n881_), .B1(new_n886_), .B2(new_n889_), .ZN(G1340gat));
  OR2_X1    g689(.A1(new_n876_), .A2(new_n878_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n380_), .A2(KEYINPUT60), .ZN(new_n892_));
  INV_X1    g691(.A(G120gat), .ZN(new_n893_));
  MUX2_X1   g692(.A(KEYINPUT60), .B(new_n892_), .S(new_n893_), .Z(new_n894_));
  NAND3_X1  g693(.A1(new_n891_), .A2(new_n799_), .A3(new_n894_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n381_), .B1(new_n882_), .B2(new_n884_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n896_), .B1(new_n879_), .B2(KEYINPUT59), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n895_), .B1(new_n897_), .B2(new_n893_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(KEYINPUT124), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT124), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n900_), .B(new_n895_), .C1(new_n897_), .C2(new_n893_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n901_), .ZN(G1341gat));
  INV_X1    g701(.A(G127gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n880_), .A2(new_n903_), .A3(new_n716_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n886_), .A2(new_n716_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n903_), .ZN(G1342gat));
  INV_X1    g705(.A(G134gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n880_), .A2(new_n907_), .A3(new_n664_), .ZN(new_n908_));
  AND2_X1   g707(.A1(new_n886_), .A2(new_n305_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n907_), .ZN(G1343gat));
  INV_X1    g709(.A(new_n586_), .ZN(new_n911_));
  NOR4_X1   g710(.A1(new_n798_), .A2(new_n911_), .A3(new_n683_), .A4(new_n460_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n891_), .A2(new_n667_), .A3(new_n912_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g713(.A1(new_n891_), .A2(new_n381_), .A3(new_n912_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g715(.A1(new_n891_), .A2(new_n716_), .A3(new_n912_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT61), .B(G155gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1346gat));
  NAND2_X1  g718(.A1(new_n891_), .A2(new_n912_), .ZN(new_n920_));
  OAI21_X1  g719(.A(G162gat), .B1(new_n920_), .B2(new_n711_), .ZN(new_n921_));
  OR2_X1    g720(.A1(new_n296_), .A2(G162gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n920_), .B2(new_n922_), .ZN(G1347gat));
  INV_X1    g722(.A(new_n882_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n683_), .A2(new_n460_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n661_), .A2(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n924_), .A2(new_n700_), .A3(new_n926_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  AOI211_X1 g727(.A(KEYINPUT62), .B(new_n421_), .C1(new_n928_), .C2(new_n667_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n928_), .A2(new_n667_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n931_), .B2(G169gat), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n928_), .A2(new_n667_), .A3(new_n485_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n929_), .B1(new_n932_), .B2(new_n933_), .ZN(G1348gat));
  AOI21_X1  g733(.A(G176gat), .B1(new_n928_), .B2(new_n381_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n891_), .A2(new_n911_), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  NOR4_X1   g736(.A1(new_n661_), .A2(new_n925_), .A3(new_n422_), .A4(new_n380_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n935_), .B1(new_n937_), .B2(new_n938_), .ZN(G1349gat));
  NOR3_X1   g738(.A1(new_n927_), .A2(new_n478_), .A3(new_n350_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT125), .ZN(new_n941_));
  OR2_X1    g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n926_), .A2(new_n716_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n410_), .B1(new_n936_), .B2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n940_), .A2(new_n941_), .ZN(new_n945_));
  AND3_X1   g744(.A1(new_n942_), .A2(new_n944_), .A3(new_n945_), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n927_), .B2(new_n711_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n664_), .A2(new_n479_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n947_), .B1(new_n927_), .B2(new_n948_), .ZN(G1351gat));
  NOR4_X1   g748(.A1(new_n911_), .A2(new_n611_), .A3(new_n519_), .A4(new_n460_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n891_), .A2(new_n667_), .A3(new_n950_), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g751(.A1(new_n891_), .A2(new_n381_), .A3(new_n950_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(new_n953_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g753(.A(new_n350_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(KEYINPUT126), .ZN(new_n956_));
  NAND3_X1  g755(.A1(new_n891_), .A2(new_n950_), .A3(new_n956_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n958_));
  XOR2_X1   g757(.A(new_n957_), .B(new_n958_), .Z(G1354gat));
  OAI211_X1 g758(.A(new_n664_), .B(new_n950_), .C1(new_n876_), .C2(new_n878_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n960_), .A2(KEYINPUT127), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n961_), .A2(G218gat), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n960_), .A2(KEYINPUT127), .ZN(new_n963_));
  AND2_X1   g762(.A1(new_n891_), .A2(new_n950_), .ZN(new_n964_));
  AND2_X1   g763(.A1(new_n305_), .A2(G218gat), .ZN(new_n965_));
  AOI22_X1  g764(.A1(new_n962_), .A2(new_n963_), .B1(new_n964_), .B2(new_n965_), .ZN(G1355gat));
endmodule


