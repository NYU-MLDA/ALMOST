//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 0 1 1 0 0 0 1 1 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n925_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT69), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G134gat), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n204_), .A2(G162gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT36), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(G162gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(G29gat), .B(G36gat), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(G43gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(G43gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(G50gat), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  AOI21_X1  g013(.A(G50gat), .B1(new_n211_), .B2(new_n212_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OR2_X1    g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  AND2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G99gat), .A2(G106gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT6), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT6), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(G99gat), .A3(G106gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  INV_X1    g024(.A(G99gat), .ZN(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n219_), .B1(new_n224_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT8), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n233_), .B(new_n219_), .C1(new_n224_), .C2(new_n230_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n218_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT9), .ZN(new_n237_));
  AOI22_X1  g036(.A1(new_n221_), .A2(new_n223_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n226_), .A2(KEYINPUT10), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n226_), .A2(KEYINPUT10), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n227_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n217_), .A2(KEYINPUT9), .A3(new_n218_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n238_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n216_), .A2(new_n235_), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n238_), .A2(new_n241_), .A3(KEYINPUT65), .A4(new_n242_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n235_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n249_), .A2(new_n235_), .A3(KEYINPUT66), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT15), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n255_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n215_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(new_n213_), .A3(KEYINPUT15), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n245_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(G232gat), .A2(G233gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT34), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT35), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n263_), .A2(new_n264_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n260_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n249_), .A2(new_n235_), .A3(KEYINPUT66), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT66), .B1(new_n249_), .B2(new_n235_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n259_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(new_n244_), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT68), .B1(new_n272_), .B2(new_n265_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n274_));
  AOI211_X1 g073(.A(new_n274_), .B(new_n266_), .C1(new_n271_), .C2(new_n244_), .ZN(new_n275_));
  OAI211_X1 g074(.A(new_n209_), .B(new_n268_), .C1(new_n273_), .C2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n260_), .B2(new_n266_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n272_), .A2(KEYINPUT68), .A3(new_n265_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n272_), .A2(new_n265_), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n277_), .A2(new_n278_), .B1(new_n279_), .B2(new_n267_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n204_), .B(G162gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(KEYINPUT36), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n208_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT70), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(new_n285_), .A3(new_n208_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n276_), .B1(new_n280_), .B2(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(KEYINPUT71), .B1(new_n288_), .B2(KEYINPUT37), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(KEYINPUT37), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT37), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n276_), .B(new_n291_), .C1(new_n280_), .C2(new_n283_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n289_), .B1(new_n293_), .B2(KEYINPUT71), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G127gat), .B(G155gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G183gat), .B(G211gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n297_), .B(new_n298_), .Z(new_n299_));
  XOR2_X1   g098(.A(new_n299_), .B(KEYINPUT17), .Z(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT72), .B(G15gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(G22gat), .ZN(new_n302_));
  INV_X1    g101(.A(G1gat), .ZN(new_n303_));
  INV_X1    g102(.A(G8gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT14), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT73), .B(KEYINPUT74), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G1gat), .B(G8gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n306_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n306_), .A2(new_n309_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G71gat), .B(G78gat), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G57gat), .B(G64gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT11), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n315_), .A2(KEYINPUT11), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n313_), .A2(KEYINPUT11), .A3(new_n315_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G231gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n312_), .B(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n300_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n299_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(KEYINPUT17), .A3(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n294_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(KEYINPUT25), .B(G183gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT26), .B(G190gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT23), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(G169gat), .ZN(new_n337_));
  INV_X1    g136(.A(G176gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n339_), .A2(KEYINPUT24), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n339_), .A2(KEYINPUT24), .A3(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n331_), .A2(new_n336_), .A3(new_n340_), .A4(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT22), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n345_), .B1(new_n346_), .B2(G169gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n337_), .A2(KEYINPUT78), .A3(KEYINPUT22), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(G169gat), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n338_), .A4(new_n349_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n350_), .A2(KEYINPUT79), .A3(new_n341_), .ZN(new_n351_));
  AOI21_X1  g150(.A(KEYINPUT79), .B1(new_n350_), .B2(new_n341_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n334_), .A2(new_n354_), .A3(new_n335_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT80), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n344_), .B1(new_n353_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT86), .ZN(new_n359_));
  INV_X1    g158(.A(G197gat), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n360_), .A2(G204gat), .ZN(new_n361_));
  INV_X1    g160(.A(G204gat), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n362_), .A2(G197gat), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n359_), .B(KEYINPUT21), .C1(new_n361_), .C2(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G197gat), .B(G204gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT21), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G211gat), .B(G218gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n364_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n365_), .ZN(new_n370_));
  XOR2_X1   g169(.A(G211gat), .B(G218gat), .Z(new_n371_));
  NAND4_X1  g170(.A1(new_n370_), .A2(new_n371_), .A3(new_n359_), .A4(KEYINPUT21), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n369_), .A2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT87), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n369_), .A2(new_n372_), .A3(KEYINPUT87), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT92), .B1(new_n358_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n376_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT87), .B1(new_n369_), .B2(new_n372_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n350_), .A2(KEYINPUT79), .A3(new_n341_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n350_), .A2(new_n341_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n357_), .A2(new_n382_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n343_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT92), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n381_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n378_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n373_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n355_), .A2(KEYINPUT91), .ZN(new_n392_));
  INV_X1    g191(.A(new_n341_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT22), .B(G169gat), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n393_), .B1(new_n394_), .B2(new_n338_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT91), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n334_), .A2(new_n354_), .A3(new_n396_), .A4(new_n335_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n392_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n391_), .A2(new_n343_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G226gat), .A2(G233gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT19), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n399_), .A2(KEYINPUT20), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n390_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT18), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G64gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(new_n408_), .B(G92gat), .Z(new_n409_));
  NAND2_X1  g208(.A1(new_n398_), .A2(new_n343_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n373_), .ZN(new_n411_));
  OAI211_X1 g210(.A(KEYINPUT20), .B(new_n411_), .C1(new_n381_), .C2(new_n387_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(new_n401_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n405_), .A2(new_n409_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n409_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n403_), .B1(new_n378_), .B2(new_n389_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT20), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n358_), .B2(new_n377_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n402_), .B1(new_n418_), .B2(new_n411_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n415_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT27), .B1(new_n414_), .B2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(KEYINPUT95), .B1(new_n398_), .B2(new_n343_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n398_), .A2(KEYINPUT95), .A3(new_n343_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n423_), .A2(new_n391_), .A3(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n425_), .A2(KEYINPUT96), .A3(KEYINPUT20), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT96), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n398_), .A2(KEYINPUT95), .A3(new_n343_), .ZN(new_n428_));
  NOR3_X1   g227(.A1(new_n428_), .A2(new_n422_), .A3(new_n373_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n427_), .B1(new_n429_), .B2(new_n417_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n390_), .A2(new_n426_), .A3(new_n430_), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n431_), .A2(new_n401_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n412_), .A2(new_n401_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n415_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT27), .ZN(new_n435_));
  AOI22_X1  g234(.A1(new_n390_), .A2(new_n404_), .B1(new_n401_), .B2(new_n412_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n436_), .B2(new_n409_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n421_), .B1(new_n434_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT97), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G225gat), .A2(G233gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n442_));
  AND3_X1   g241(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT84), .B1(G155gat), .B2(G162gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT1), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G155gat), .A2(G162gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT84), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT1), .ZN(new_n449_));
  NAND3_X1  g248(.A1(KEYINPUT84), .A2(G155gat), .A3(G162gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(G155gat), .A2(G162gat), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n445_), .A2(new_n451_), .A3(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(G141gat), .B(G148gat), .Z(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT3), .ZN(new_n457_));
  INV_X1    g256(.A(G141gat), .ZN(new_n458_));
  INV_X1    g257(.A(G148gat), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G141gat), .A2(G148gat), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT2), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n460_), .A2(new_n463_), .A3(new_n464_), .A4(new_n465_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n452_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n466_), .A2(KEYINPUT85), .A3(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(KEYINPUT85), .B1(new_n466_), .B2(new_n467_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n456_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT81), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G127gat), .A2(G134gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(G127gat), .A2(G134gat), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n471_), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  XOR2_X1   g274(.A(G113gat), .B(G120gat), .Z(new_n476_));
  INV_X1    g275(.A(G127gat), .ZN(new_n477_));
  INV_X1    g276(.A(G134gat), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(KEYINPUT81), .A3(new_n472_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n475_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n476_), .B1(new_n475_), .B2(new_n480_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT82), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT82), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n470_), .A2(new_n484_), .A3(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n475_), .A2(new_n480_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G113gat), .B(G120gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n481_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n491_), .B(new_n456_), .C1(new_n469_), .C2(new_n468_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n442_), .B1(new_n487_), .B2(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n481_), .A2(new_n485_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n494_), .B1(KEYINPUT82), .B2(new_n491_), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT4), .B1(new_n495_), .B2(new_n470_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n441_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(KEYINPUT93), .B(G85gat), .Z(new_n498_));
  XNOR2_X1  g297(.A(G1gat), .B(G29gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT0), .B(G57gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n487_), .A2(new_n440_), .A3(new_n492_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n497_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n502_), .B1(new_n497_), .B2(new_n503_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n439_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n497_), .A2(new_n503_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n502_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n497_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n509_), .A2(KEYINPUT97), .A3(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n506_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT89), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n466_), .A2(new_n467_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT85), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n466_), .A2(new_n467_), .A3(KEYINPUT85), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n516_), .A2(new_n517_), .B1(new_n455_), .B2(new_n454_), .ZN(new_n518_));
  XOR2_X1   g317(.A(KEYINPUT88), .B(KEYINPUT29), .Z(new_n519_));
  OAI21_X1  g318(.A(new_n513_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n519_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n470_), .A2(KEYINPUT89), .A3(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n373_), .A3(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(G228gat), .A2(G233gat), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n524_), .B1(new_n470_), .B2(KEYINPUT29), .ZN(new_n525_));
  AOI22_X1  g324(.A1(new_n523_), .A2(new_n524_), .B1(new_n381_), .B2(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G78gat), .B(G106gat), .Z(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT90), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  OR3_X1    g327(.A1(new_n470_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT28), .B1(new_n470_), .B2(KEYINPUT29), .ZN(new_n530_));
  XOR2_X1   g329(.A(G22gat), .B(G50gat), .Z(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n531_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n523_), .A2(new_n524_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n525_), .A2(new_n381_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n536_), .A2(new_n527_), .A3(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n527_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n539_));
  OAI22_X1  g338(.A1(new_n528_), .A2(new_n535_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n536_), .A2(new_n537_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n527_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n533_), .A2(new_n534_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n526_), .A2(new_n527_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n543_), .A2(new_n544_), .A3(KEYINPUT90), .A4(new_n545_), .ZN(new_n546_));
  XOR2_X1   g345(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n547_));
  NAND2_X1  g346(.A1(G227gat), .A2(G233gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G15gat), .B(G43gat), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n549_), .B(new_n550_), .Z(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G71gat), .B(G99gat), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n553_), .B(KEYINPUT30), .Z(new_n554_));
  NOR2_X1   g353(.A1(new_n358_), .A2(new_n554_), .ZN(new_n555_));
  AND3_X1   g354(.A1(new_n386_), .A2(new_n554_), .A3(new_n343_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n495_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR3_X1   g357(.A1(new_n555_), .A2(new_n556_), .A3(new_n495_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n552_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n559_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(new_n557_), .A3(new_n551_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n540_), .A2(new_n546_), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n563_), .B1(new_n540_), .B2(new_n546_), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n438_), .B(new_n512_), .C1(new_n564_), .C2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n433_), .B1(new_n431_), .B2(new_n401_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n409_), .A2(KEYINPUT32), .ZN(new_n568_));
  OAI22_X1  g367(.A1(new_n567_), .A2(new_n568_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n436_), .A2(new_n568_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT33), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n510_), .A2(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n497_), .A2(KEYINPUT33), .A3(new_n502_), .A4(new_n503_), .ZN(new_n573_));
  NAND4_X1  g372(.A1(new_n572_), .A2(new_n414_), .A3(new_n420_), .A4(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n487_), .A2(new_n492_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT94), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n441_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n440_), .B1(new_n493_), .B2(new_n496_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n577_), .A2(new_n508_), .A3(new_n578_), .ZN(new_n579_));
  OAI22_X1  g378(.A1(new_n569_), .A2(new_n570_), .B1(new_n574_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n563_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n546_), .B2(new_n540_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n566_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT76), .ZN(new_n585_));
  INV_X1    g384(.A(new_n216_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n312_), .A2(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n310_), .A2(new_n311_), .A3(new_n216_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(G229gat), .A2(G233gat), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n589_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n259_), .A2(new_n312_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(new_n590_), .A3(new_n588_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n585_), .B1(new_n592_), .B2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n585_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G113gat), .B(G141gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT77), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(new_n337_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(new_n360_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n596_), .A2(new_n597_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n597_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n601_), .B1(new_n595_), .B2(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n320_), .A2(KEYINPUT12), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n607_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n320_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n235_), .A2(new_n609_), .A3(new_n243_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT12), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n235_), .A2(new_n243_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n320_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT64), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n608_), .A2(new_n614_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n613_), .A2(new_n610_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n622_));
  XNOR2_X1  g421(.A(G120gat), .B(G148gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G176gat), .B(G204gat), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n624_), .B(new_n625_), .Z(new_n626_));
  NAND2_X1  g425(.A1(new_n621_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n626_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n618_), .A2(new_n620_), .A3(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT13), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n627_), .A2(KEYINPUT13), .A3(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n606_), .A2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n584_), .A2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n328_), .A2(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT98), .Z(new_n638_));
  INV_X1    g437(.A(new_n512_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n303_), .A3(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT38), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n276_), .B1(new_n280_), .B2(new_n283_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(new_n327_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n636_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(new_n639_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(G1gat), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n641_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT99), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT99), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n641_), .A2(new_n650_), .A3(new_n647_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(G1324gat));
  INV_X1    g451(.A(new_n438_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n304_), .B1(new_n645_), .B2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(KEYINPUT100), .B(KEYINPUT39), .Z(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n438_), .A2(G8gat), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n638_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT40), .ZN(G1325gat));
  INV_X1    g458(.A(G15gat), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n638_), .A2(new_n660_), .A3(new_n581_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT101), .Z(new_n662_));
  AOI21_X1  g461(.A(new_n660_), .B1(new_n645_), .B2(new_n581_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT41), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n662_), .A2(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n540_), .A2(new_n546_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n666_), .B1(new_n645_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT42), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n667_), .A2(G22gat), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n638_), .B2(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n672_), .B(KEYINPUT102), .ZN(G1327gat));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n584_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n292_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n268_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n677_));
  AND3_X1   g476(.A1(new_n282_), .A2(new_n285_), .A3(new_n208_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n285_), .B1(new_n282_), .B2(new_n208_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n677_), .A2(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n291_), .B1(new_n681_), .B2(new_n276_), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT71), .B1(new_n676_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n289_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT106), .B1(new_n675_), .B2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT43), .B1(new_n566_), .B2(new_n583_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n294_), .A3(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690_));
  INV_X1    g489(.A(new_n421_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n437_), .B1(new_n567_), .B2(new_n409_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n512_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n565_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n540_), .A2(new_n546_), .A3(new_n563_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n693_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n580_), .A2(new_n582_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n690_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n566_), .A2(new_n583_), .A3(KEYINPUT105), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(new_n294_), .A3(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n701_));
  AOI22_X1  g500(.A1(new_n686_), .A2(new_n689_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n635_), .A2(new_n327_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT103), .Z(new_n704_));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705_));
  OAI22_X1  g504(.A1(new_n702_), .A2(new_n704_), .B1(new_n705_), .B2(KEYINPUT44), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n698_), .A2(new_n294_), .A3(new_n699_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n701_), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n687_), .A2(new_n294_), .A3(new_n688_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n688_), .B1(new_n687_), .B2(new_n294_), .ZN(new_n710_));
  OAI22_X1  g509(.A1(new_n707_), .A2(new_n708_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n705_), .A2(KEYINPUT44), .ZN(new_n712_));
  INV_X1    g511(.A(new_n704_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n711_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n706_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G29gat), .B1(new_n716_), .B2(new_n512_), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n636_), .A2(new_n643_), .A3(new_n327_), .ZN(new_n718_));
  INV_X1    g517(.A(G29gat), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n639_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n717_), .A2(new_n720_), .ZN(G1328gat));
  INV_X1    g520(.A(G36gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n715_), .B2(new_n653_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n718_), .A2(new_n722_), .A3(new_n653_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT45), .Z(new_n725_));
  NOR2_X1   g524(.A1(new_n723_), .A2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT46), .ZN(G1329gat));
  NAND3_X1  g526(.A1(new_n715_), .A2(G43gat), .A3(new_n581_), .ZN(new_n728_));
  AOI21_X1  g527(.A(G43gat), .B1(new_n718_), .B2(new_n581_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT108), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n715_), .B2(new_n668_), .ZN(new_n734_));
  AOI211_X1 g533(.A(KEYINPUT109), .B(new_n667_), .C1(new_n706_), .C2(new_n714_), .ZN(new_n735_));
  INV_X1    g534(.A(G50gat), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n718_), .A2(new_n736_), .A3(new_n668_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT110), .B1(new_n737_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n734_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n715_), .A2(new_n733_), .A3(new_n668_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(G50gat), .A3(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT110), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(new_n738_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n740_), .A2(new_n745_), .ZN(G1331gat));
  INV_X1    g545(.A(new_n606_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n634_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n584_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n328_), .A2(new_n750_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT111), .Z(new_n752_));
  AOI21_X1  g551(.A(G57gat), .B1(new_n752_), .B2(new_n639_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n750_), .A2(new_n644_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT112), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n639_), .A2(G57gat), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n753_), .B1(new_n755_), .B2(new_n756_), .ZN(G1332gat));
  INV_X1    g556(.A(G64gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n755_), .B2(new_n653_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT48), .Z(new_n760_));
  NAND3_X1  g559(.A1(new_n752_), .A2(new_n758_), .A3(new_n653_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1333gat));
  INV_X1    g561(.A(G71gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n755_), .B2(new_n581_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT49), .Z(new_n765_));
  NAND3_X1  g564(.A1(new_n752_), .A2(new_n763_), .A3(new_n581_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1334gat));
  INV_X1    g566(.A(G78gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n755_), .B2(new_n668_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT50), .Z(new_n770_));
  NAND3_X1  g569(.A1(new_n752_), .A2(new_n768_), .A3(new_n668_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1335gat));
  NAND2_X1  g571(.A1(new_n749_), .A2(new_n327_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n686_), .A2(new_n689_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n700_), .A2(new_n701_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n773_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n776_), .A2(G85gat), .A3(new_n639_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n750_), .A2(new_n643_), .A3(new_n327_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n778_), .A2(new_n639_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n777_), .B1(G85gat), .B2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT113), .ZN(G1336gat));
  NAND3_X1  g580(.A1(new_n776_), .A2(G92gat), .A3(new_n653_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n778_), .A2(new_n653_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n782_), .B1(G92gat), .B2(new_n783_), .ZN(new_n784_));
  XOR2_X1   g583(.A(new_n784_), .B(KEYINPUT114), .Z(G1337gat));
  OAI211_X1 g584(.A(new_n778_), .B(new_n581_), .C1(new_n239_), .C2(new_n240_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT115), .Z(new_n787_));
  NOR3_X1   g586(.A1(new_n702_), .A2(new_n563_), .A3(new_n773_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n787_), .B1(new_n788_), .B2(new_n226_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g589(.A1(new_n778_), .A2(new_n227_), .A3(new_n668_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(new_n776_), .B2(new_n668_), .ZN(new_n794_));
  NOR4_X1   g593(.A1(new_n702_), .A2(KEYINPUT116), .A3(new_n667_), .A4(new_n773_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n792_), .B1(new_n796_), .B2(G106gat), .ZN(new_n797_));
  NOR4_X1   g596(.A1(new_n794_), .A2(new_n795_), .A3(KEYINPUT52), .A4(new_n227_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n791_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT53), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(new_n791_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1339gat));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n618_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n608_), .A2(new_n614_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n808_), .A2(new_n617_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n805_), .B1(new_n618_), .B2(new_n804_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n807_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  OAI22_X1  g610(.A1(new_n811_), .A2(new_n628_), .B1(KEYINPUT118), .B2(KEYINPUT56), .ZN(new_n812_));
  INV_X1    g611(.A(new_n629_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n813_), .B1(new_n603_), .B2(new_n605_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n618_), .A2(new_n804_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(KEYINPUT55), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n816_), .B(new_n806_), .C1(new_n617_), .C2(new_n808_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n626_), .A3(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n812_), .A2(new_n814_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n589_), .A2(new_n590_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n593_), .A2(new_n591_), .A3(new_n588_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n601_), .A3(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n603_), .A2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n630_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n820_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT57), .B1(new_n826_), .B2(new_n642_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT57), .ZN(new_n828_));
  AOI211_X1 g627(.A(new_n828_), .B(new_n643_), .C1(new_n820_), .C2(new_n825_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT56), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n817_), .A2(new_n831_), .A3(new_n626_), .ZN(new_n832_));
  AND2_X1   g631(.A1(new_n832_), .A2(new_n629_), .ZN(new_n833_));
  OAI21_X1  g632(.A(KEYINPUT56), .B1(new_n811_), .B2(new_n628_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n833_), .A2(KEYINPUT58), .A3(new_n824_), .A4(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n824_), .A2(new_n834_), .A3(new_n629_), .A4(new_n832_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT58), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n294_), .A2(new_n835_), .A3(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n294_), .A2(new_n835_), .A3(new_n838_), .A4(KEYINPUT119), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n830_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n327_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n327_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n685_), .A2(new_n606_), .A3(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT54), .B1(new_n846_), .B2(new_n634_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848_));
  NAND4_X1  g647(.A1(new_n328_), .A2(new_n848_), .A3(new_n606_), .A4(new_n748_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n844_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n438_), .A2(new_n639_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n852_), .A2(new_n694_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT59), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n830_), .A2(new_n839_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n850_), .B1(new_n856_), .B2(new_n845_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n857_), .A2(new_n858_), .A3(new_n853_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n855_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(G113gat), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n860_), .A2(new_n861_), .A3(new_n606_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n854_), .B2(new_n606_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n863_), .A2(KEYINPUT120), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n863_), .A2(KEYINPUT120), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n862_), .A2(new_n864_), .A3(new_n865_), .ZN(G1340gat));
  AOI22_X1  g665(.A1(new_n843_), .A2(new_n327_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n867_), .A2(new_n694_), .A3(new_n852_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n748_), .A2(G120gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(KEYINPUT60), .B2(new_n869_), .ZN(new_n870_));
  AND4_X1   g669(.A1(new_n634_), .A2(new_n870_), .A3(new_n855_), .A4(new_n859_), .ZN(new_n871_));
  INV_X1    g670(.A(G120gat), .ZN(new_n872_));
  OAI22_X1  g671(.A1(new_n871_), .A2(new_n872_), .B1(KEYINPUT60), .B2(new_n870_), .ZN(G1341gat));
  AOI21_X1  g672(.A(G127gat), .B1(new_n868_), .B2(new_n845_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n860_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n327_), .A2(new_n477_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT121), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n874_), .B1(new_n875_), .B2(new_n877_), .ZN(G1342gat));
  AOI21_X1  g677(.A(G134gat), .B1(new_n868_), .B2(new_n643_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n685_), .A2(new_n478_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n875_), .B2(new_n880_), .ZN(G1343gat));
  NAND2_X1  g680(.A1(new_n851_), .A2(new_n564_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n882_), .A2(new_n852_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n747_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n634_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g686(.A1(new_n883_), .A2(new_n845_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT61), .B(G155gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1346gat));
  AOI21_X1  g689(.A(G162gat), .B1(new_n883_), .B2(new_n643_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n294_), .A2(G162gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n883_), .B2(new_n892_), .ZN(G1347gat));
  NOR2_X1   g692(.A1(new_n438_), .A2(new_n639_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n581_), .ZN(new_n895_));
  XOR2_X1   g694(.A(new_n895_), .B(KEYINPUT122), .Z(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n857_), .A2(new_n667_), .A3(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n898_), .A2(KEYINPUT123), .A3(new_n747_), .ZN(new_n899_));
  NAND4_X1  g698(.A1(new_n857_), .A2(new_n747_), .A3(new_n667_), .A4(new_n897_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n899_), .A2(G169gat), .A3(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n898_), .A2(new_n747_), .A3(new_n394_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n899_), .A2(KEYINPUT62), .A3(G169gat), .A4(new_n902_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(G1348gat));
  NOR2_X1   g707(.A1(new_n867_), .A2(new_n668_), .ZN(new_n909_));
  AND4_X1   g708(.A1(G176gat), .A2(new_n909_), .A3(new_n634_), .A4(new_n897_), .ZN(new_n910_));
  AOI21_X1  g709(.A(G176gat), .B1(new_n898_), .B2(new_n634_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT124), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(KEYINPUT124), .B1(new_n910_), .B2(new_n911_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1349gat));
  INV_X1    g715(.A(new_n329_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n896_), .A2(new_n327_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n857_), .A2(new_n667_), .A3(new_n917_), .A4(new_n918_), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n919_), .B(KEYINPUT125), .Z(new_n920_));
  AOI21_X1  g719(.A(G183gat), .B1(new_n909_), .B2(new_n918_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1350gat));
  INV_X1    g721(.A(new_n898_), .ZN(new_n923_));
  OAI21_X1  g722(.A(G190gat), .B1(new_n923_), .B2(new_n685_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n898_), .A2(new_n330_), .A3(new_n643_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(G1351gat));
  INV_X1    g725(.A(new_n894_), .ZN(new_n927_));
  NOR4_X1   g726(.A1(new_n867_), .A2(new_n606_), .A3(new_n695_), .A4(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(KEYINPUT127), .B1(new_n928_), .B2(KEYINPUT126), .ZN(new_n929_));
  AOI21_X1  g728(.A(G197gat), .B1(new_n928_), .B2(KEYINPUT126), .ZN(new_n930_));
  NAND4_X1  g729(.A1(new_n851_), .A2(new_n747_), .A3(new_n564_), .A4(new_n894_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT126), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n931_), .A2(new_n932_), .A3(new_n933_), .ZN(new_n934_));
  AND3_X1   g733(.A1(new_n929_), .A2(new_n930_), .A3(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n930_), .B1(new_n934_), .B2(new_n929_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1352gat));
  NOR2_X1   g736(.A1(new_n882_), .A2(new_n927_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n634_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G204gat), .ZN(G1353gat));
  NOR3_X1   g739(.A1(new_n882_), .A2(new_n327_), .A3(new_n927_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n941_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n942_));
  XOR2_X1   g741(.A(KEYINPUT63), .B(G211gat), .Z(new_n943_));
  AOI21_X1  g742(.A(new_n942_), .B1(new_n941_), .B2(new_n943_), .ZN(G1354gat));
  AOI21_X1  g743(.A(G218gat), .B1(new_n938_), .B2(new_n643_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n294_), .A2(G218gat), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(new_n938_), .B2(new_n946_), .ZN(G1355gat));
endmodule


