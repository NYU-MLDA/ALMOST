//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n914_, new_n915_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT21), .ZN(new_n205_));
  NOR3_X1   g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(new_n203_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT98), .ZN(new_n209_));
  AND2_X1   g008(.A1(G197gat), .A2(G204gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G197gat), .A2(G204gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n209_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(new_n205_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n209_), .B(KEYINPUT21), .C1(new_n210_), .C2(new_n211_), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n208_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT99), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  AOI211_X1 g016(.A(KEYINPUT99), .B(new_n208_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n207_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G183gat), .A2(G190gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(KEYINPUT86), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT86), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n222_), .A2(G183gat), .A3(G190gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n223_), .A3(KEYINPUT23), .ZN(new_n224_));
  INV_X1    g023(.A(new_n220_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT93), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n221_), .A2(new_n223_), .A3(KEYINPUT93), .A4(KEYINPUT23), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n228_), .A2(new_n230_), .A3(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G169gat), .A2(G176gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT22), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n235_), .A2(KEYINPUT89), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(KEYINPUT89), .ZN(new_n237_));
  OAI21_X1  g036(.A(G169gat), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT90), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT91), .B(G176gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT22), .B1(KEYINPUT88), .B2(G169gat), .ZN(new_n243_));
  AND2_X1   g042(.A1(KEYINPUT88), .A2(G169gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  OAI211_X1 g045(.A(KEYINPUT90), .B(G169gat), .C1(new_n236_), .C2(new_n237_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n240_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT92), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n240_), .A2(new_n246_), .A3(KEYINPUT92), .A4(new_n247_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n234_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(G169gat), .ZN(new_n253_));
  INV_X1    g052(.A(G176gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n255_), .A2(KEYINPUT24), .ZN(new_n256_));
  INV_X1    g055(.A(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT23), .B1(new_n221_), .B2(new_n223_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n225_), .A2(new_n226_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n257_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT87), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT87), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n257_), .B(new_n262_), .C1(new_n258_), .C2(new_n259_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT25), .B(G183gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT26), .B(G190gat), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n233_), .A2(KEYINPUT24), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n264_), .A2(new_n265_), .B1(new_n266_), .B2(new_n255_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n261_), .A2(new_n263_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n219_), .B1(new_n252_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT20), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT21), .B1(new_n204_), .B2(new_n209_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n214_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n203_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT99), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n215_), .A2(new_n216_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n206_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  AND2_X1   g076(.A1(new_n267_), .A2(new_n257_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n228_), .A2(new_n231_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n230_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT22), .B(G169gat), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n241_), .A2(new_n281_), .B1(G169gat), .B2(G176gat), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n278_), .A2(new_n279_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n271_), .B1(new_n277_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT100), .B(KEYINPUT19), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G226gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n270_), .A2(new_n284_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n234_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n241_), .B1(new_n244_), .B2(new_n243_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n239_), .B2(new_n238_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT92), .B1(new_n292_), .B2(new_n247_), .ZN(new_n293_));
  AND4_X1   g092(.A1(KEYINPUT92), .A2(new_n240_), .A3(new_n246_), .A4(new_n247_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n290_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n295_), .A2(new_n277_), .A3(new_n268_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n278_), .A2(new_n279_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n280_), .A2(new_n282_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n271_), .B1(new_n219_), .B2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n288_), .B1(new_n296_), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G8gat), .B(G36gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n302_), .B(KEYINPUT18), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G64gat), .B(G92gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n289_), .A2(new_n301_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n305_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n252_), .A2(new_n219_), .A3(new_n269_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT20), .B1(new_n277_), .B2(new_n283_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n287_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n270_), .A2(new_n284_), .A3(new_n288_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n307_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n202_), .B1(new_n306_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT107), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT107), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n315_), .B(new_n202_), .C1(new_n306_), .C2(new_n312_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n310_), .A2(new_n311_), .A3(new_n307_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n296_), .A2(new_n300_), .A3(new_n288_), .ZN(new_n319_));
  AND2_X1   g118(.A1(new_n270_), .A2(new_n284_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n319_), .B1(new_n320_), .B2(new_n288_), .ZN(new_n321_));
  AND3_X1   g120(.A1(new_n321_), .A2(KEYINPUT106), .A3(new_n305_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT106), .B1(new_n321_), .B2(new_n305_), .ZN(new_n323_));
  OAI211_X1 g122(.A(KEYINPUT27), .B(new_n318_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n317_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT95), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(KEYINPUT95), .A2(G155gat), .A3(G162gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(G155gat), .ZN(new_n331_));
  INV_X1    g130(.A(G162gat), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n330_), .A2(KEYINPUT1), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n328_), .A2(new_n334_), .A3(new_n329_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G141gat), .A2(G148gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT94), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT94), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(G141gat), .A3(G148gat), .ZN(new_n340_));
  OR2_X1    g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n338_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n336_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(KEYINPUT96), .A3(KEYINPUT3), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT96), .ZN(new_n346_));
  NOR2_X1   g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT3), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n346_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT2), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n337_), .A2(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(new_n348_), .B2(new_n347_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n338_), .A2(new_n340_), .A3(new_n351_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n350_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n330_), .B1(G155gat), .B2(G162gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n344_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(KEYINPUT29), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n360_), .B(KEYINPUT28), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n277_), .B1(KEYINPUT29), .B2(new_n359_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  AND2_X1   g162(.A1(KEYINPUT97), .A2(G228gat), .ZN(new_n364_));
  NOR2_X1   g163(.A1(KEYINPUT97), .A2(G228gat), .ZN(new_n365_));
  OAI21_X1  g164(.A(G233gat), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(G78gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G106gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G22gat), .B(G50gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n370_), .B(new_n371_), .ZN(new_n372_));
  OR2_X1    g171(.A1(new_n363_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n363_), .A2(new_n372_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n325_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n295_), .A2(new_n268_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G71gat), .B(G99gat), .ZN(new_n379_));
  INV_X1    g178(.A(G43gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n378_), .B(new_n381_), .ZN(new_n382_));
  XOR2_X1   g181(.A(G127gat), .B(G134gat), .Z(new_n383_));
  XOR2_X1   g182(.A(G113gat), .B(G120gat), .Z(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n382_), .B(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(G227gat), .A2(G233gat), .ZN(new_n387_));
  INV_X1    g186(.A(G15gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT30), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT31), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n386_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n386_), .A2(new_n391_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n385_), .ZN(new_n396_));
  OAI22_X1  g195(.A1(new_n341_), .A2(KEYINPUT3), .B1(new_n351_), .B2(new_n337_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n349_), .B2(new_n345_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n356_), .B1(new_n398_), .B2(new_n354_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n342_), .B1(new_n333_), .B2(new_n335_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n396_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n344_), .A2(new_n358_), .A3(new_n385_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G225gat), .A2(G233gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n401_), .A2(KEYINPUT4), .A3(new_n402_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n404_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n359_), .A2(new_n408_), .A3(new_n396_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n406_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G1gat), .B(G29gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G85gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT0), .B(G57gat), .ZN(new_n413_));
  XOR2_X1   g212(.A(new_n412_), .B(new_n413_), .Z(new_n414_));
  NAND3_X1  g213(.A1(new_n405_), .A2(new_n410_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT104), .ZN(new_n416_));
  OR2_X1    g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n416_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n405_), .A2(new_n410_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n414_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n417_), .A2(new_n418_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n395_), .A2(new_n423_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n377_), .A2(new_n424_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n307_), .A2(KEYINPUT32), .ZN(new_n426_));
  OR3_X1    g225(.A1(new_n289_), .A2(new_n301_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n321_), .A2(new_n426_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n422_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT101), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n306_), .B2(new_n312_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n305_), .B1(new_n289_), .B2(new_n301_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(new_n318_), .A3(KEYINPUT101), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n415_), .B(KEYINPUT33), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n431_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n406_), .A2(new_n404_), .A3(new_n409_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(KEYINPUT102), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT102), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n406_), .A2(new_n438_), .A3(new_n404_), .A4(new_n409_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n414_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(KEYINPUT103), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT103), .B1(new_n440_), .B2(new_n441_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n429_), .B1(new_n435_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n376_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT105), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n440_), .A2(new_n441_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT103), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(new_n442_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n452_), .A2(new_n433_), .A3(new_n431_), .A4(new_n434_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n375_), .B1(new_n453_), .B2(new_n429_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT105), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n317_), .A2(new_n324_), .A3(new_n375_), .A4(new_n423_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n448_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n425_), .B1(new_n458_), .B2(new_n394_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G120gat), .B(G148gat), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT5), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G176gat), .B(G204gat), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n461_), .B(new_n462_), .Z(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G230gat), .A2(G233gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(G71gat), .B(G78gat), .Z(new_n466_));
  XNOR2_X1  g265(.A(G57gat), .B(G64gat), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n466_), .B1(KEYINPUT11), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT67), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT67), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n466_), .B(new_n470_), .C1(KEYINPUT11), .C2(new_n467_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n467_), .A2(KEYINPUT11), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n469_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n472_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(G99gat), .B2(G106gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(G99gat), .A2(G106gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n478_), .A2(KEYINPUT6), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(G85gat), .ZN(new_n481_));
  INV_X1    g280(.A(G92gat), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n481_), .A2(new_n482_), .A3(KEYINPUT9), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n480_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(KEYINPUT10), .B(G99gat), .Z(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(new_n369_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G85gat), .B(G92gat), .Z(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT9), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n484_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT8), .ZN(new_n490_));
  NOR2_X1   g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  AND2_X1   g290(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n492_));
  NOR2_X1   g291(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  OAI22_X1  g293(.A1(KEYINPUT64), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n490_), .B(new_n487_), .C1(new_n496_), .C2(new_n480_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT65), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n498_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n478_), .A2(KEYINPUT6), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n476_), .A2(G99gat), .A3(G106gat), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(new_n501_), .A3(KEYINPUT65), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n499_), .A2(new_n502_), .A3(new_n494_), .A4(new_n495_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n490_), .B1(new_n503_), .B2(new_n487_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT66), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n497_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  AOI211_X1 g305(.A(KEYINPUT66), .B(new_n490_), .C1(new_n503_), .C2(new_n487_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n475_), .B(new_n489_), .C1(new_n506_), .C2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT12), .ZN(new_n509_));
  INV_X1    g308(.A(new_n487_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT65), .B1(new_n500_), .B2(new_n501_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n496_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n510_), .B1(new_n512_), .B2(new_n502_), .ZN(new_n513_));
  OAI21_X1  g312(.A(KEYINPUT66), .B1(new_n513_), .B2(new_n490_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n504_), .A2(new_n505_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(new_n497_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n475_), .B1(new_n516_), .B2(new_n489_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n509_), .A2(new_n517_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n489_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT12), .ZN(new_n520_));
  INV_X1    g319(.A(new_n475_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n465_), .B1(new_n518_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n519_), .A2(new_n521_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(KEYINPUT68), .A3(new_n508_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n465_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n526_), .B(new_n527_), .C1(KEYINPUT68), .C2(new_n525_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n464_), .B1(new_n524_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n524_), .A2(new_n528_), .A3(new_n464_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(KEYINPUT13), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT13), .ZN(new_n533_));
  INV_X1    g332(.A(new_n531_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n533_), .B1(new_n534_), .B2(new_n529_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT69), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n532_), .A2(new_n535_), .A3(KEYINPUT69), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G29gat), .B(G36gat), .Z(new_n541_));
  XOR2_X1   g340(.A(G43gat), .B(G50gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G15gat), .B(G22gat), .ZN(new_n546_));
  INV_X1    g345(.A(G1gat), .ZN(new_n547_));
  INV_X1    g346(.A(G8gat), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT14), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT78), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT78), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n546_), .A2(new_n552_), .A3(new_n549_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G1gat), .B(G8gat), .Z(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n551_), .A2(new_n553_), .A3(new_n555_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n545_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n557_), .A2(new_n558_), .A3(new_n543_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(G229gat), .A2(G233gat), .ZN(new_n562_));
  XOR2_X1   g361(.A(new_n562_), .B(KEYINPUT83), .Z(new_n563_));
  NAND3_X1  g362(.A1(new_n560_), .A2(new_n561_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT81), .ZN(new_n565_));
  INV_X1    g364(.A(new_n561_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n543_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n543_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n559_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n570_), .A2(KEYINPUT81), .A3(new_n561_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n562_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT82), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT82), .ZN(new_n575_));
  AOI211_X1 g374(.A(new_n575_), .B(new_n562_), .C1(new_n568_), .C2(new_n571_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n564_), .B1(new_n574_), .B2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G113gat), .B(G141gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT84), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G169gat), .B(G197gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  NAND2_X1  g380(.A1(new_n577_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT85), .ZN(new_n583_));
  INV_X1    g382(.A(new_n581_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n564_), .B(new_n584_), .C1(new_n574_), .C2(new_n576_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n582_), .A2(new_n583_), .A3(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n577_), .A2(KEYINPUT85), .A3(new_n581_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n540_), .A2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n459_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT73), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n592_), .B1(new_n519_), .B2(new_n569_), .ZN(new_n593_));
  XOR2_X1   g392(.A(KEYINPUT70), .B(KEYINPUT34), .Z(new_n594_));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n593_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n519_), .A2(new_n545_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n516_), .A2(new_n543_), .A3(new_n489_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n596_), .A2(new_n597_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n599_), .A2(new_n603_), .ZN(new_n604_));
  NAND4_X1  g403(.A1(new_n600_), .A2(new_n601_), .A3(KEYINPUT73), .A4(new_n598_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G190gat), .B(G218gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT74), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n607_), .B(new_n608_), .Z(new_n609_));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n604_), .A2(new_n605_), .A3(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n609_), .A2(new_n610_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n604_), .A2(new_n605_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT75), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n614_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  AOI211_X1 g416(.A(KEYINPUT75), .B(new_n613_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n612_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT37), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT77), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT77), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(new_n623_), .A3(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n615_), .A2(new_n616_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n613_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n615_), .A2(new_n616_), .A3(new_n614_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT76), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n628_), .A2(new_n629_), .A3(KEYINPUT37), .A4(new_n612_), .ZN(new_n630_));
  OAI211_X1 g429(.A(KEYINPUT37), .B(new_n612_), .C1(new_n617_), .C2(new_n618_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(KEYINPUT76), .ZN(new_n632_));
  AOI22_X1  g431(.A1(new_n622_), .A2(new_n624_), .B1(new_n630_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(G231gat), .A2(G233gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n475_), .B(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n559_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n635_), .B(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(G127gat), .B(G155gat), .Z(new_n638_));
  XNOR2_X1  g437(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G183gat), .B(G211gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT79), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT17), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n642_), .A2(new_n643_), .A3(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n637_), .A2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n642_), .A2(new_n644_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n646_), .B1(new_n637_), .B2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n633_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n591_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(new_n547_), .A3(new_n422_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT38), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n457_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n655_));
  AND3_X1   g454(.A1(new_n446_), .A2(new_n455_), .A3(new_n376_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n394_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  OR2_X1    g456(.A1(new_n377_), .A2(new_n424_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n619_), .B(KEYINPUT108), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n649_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n590_), .ZN(new_n663_));
  AND3_X1   g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n547_), .B1(new_n664_), .B2(new_n422_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n654_), .A2(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n666_), .B1(new_n653_), .B2(new_n652_), .ZN(G1324gat));
  INV_X1    g466(.A(new_n325_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n651_), .A2(new_n548_), .A3(new_n668_), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n661_), .A2(new_n662_), .A3(new_n668_), .A4(new_n663_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT39), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(G8gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n670_), .B2(G8gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n674_), .B(new_n676_), .ZN(G1325gat));
  AOI21_X1  g476(.A(new_n388_), .B1(new_n664_), .B2(new_n395_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT41), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n651_), .A2(new_n388_), .A3(new_n395_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1326gat));
  INV_X1    g480(.A(G22gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n664_), .B2(new_n375_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT42), .Z(new_n684_));
  NAND3_X1  g483(.A1(new_n651_), .A2(new_n682_), .A3(new_n375_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1327gat));
  NOR2_X1   g485(.A1(new_n660_), .A2(new_n662_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n591_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G29gat), .B1(new_n688_), .B2(new_n422_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n622_), .A2(new_n624_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n630_), .A2(new_n632_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT43), .B1(new_n459_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n659_), .A2(new_n694_), .A3(new_n633_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n663_), .A2(new_n649_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT44), .B1(new_n696_), .B2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n700_));
  AOI211_X1 g499(.A(new_n700_), .B(new_n697_), .C1(new_n693_), .C2(new_n695_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n422_), .A2(G29gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n689_), .B1(new_n702_), .B2(new_n703_), .ZN(G1328gat));
  NOR2_X1   g503(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n705_));
  INV_X1    g504(.A(G36gat), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n706_), .B1(new_n702_), .B2(new_n668_), .ZN(new_n707_));
  NAND4_X1  g506(.A1(new_n591_), .A2(new_n706_), .A3(new_n668_), .A4(new_n687_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT45), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n707_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n705_), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n699_), .A2(new_n701_), .A3(new_n325_), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n709_), .B(new_n712_), .C1(new_n713_), .C2(new_n706_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(G1329gat));
  NOR4_X1   g514(.A1(new_n699_), .A2(new_n701_), .A3(new_n380_), .A4(new_n394_), .ZN(new_n716_));
  AOI21_X1  g515(.A(G43gat), .B1(new_n688_), .B2(new_n395_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT47), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n394_), .A2(new_n380_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n717_), .B1(new_n702_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT47), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n718_), .A2(new_n722_), .ZN(G1330gat));
  INV_X1    g522(.A(G50gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n688_), .A2(new_n724_), .A3(new_n375_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n702_), .A2(new_n726_), .A3(new_n375_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(G50gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n726_), .B1(new_n702_), .B2(new_n375_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1331gat));
  NOR3_X1   g529(.A1(new_n633_), .A2(new_n540_), .A3(new_n649_), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n731_), .A2(KEYINPUT112), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n459_), .A2(new_n589_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(KEYINPUT112), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(G57gat), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(new_n737_), .A3(new_n422_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n540_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n649_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n661_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(new_n422_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n738_), .B1(new_n742_), .B2(new_n737_), .ZN(G1332gat));
  INV_X1    g542(.A(G64gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n741_), .B2(new_n668_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT48), .Z(new_n746_));
  NAND3_X1  g545(.A1(new_n736_), .A2(new_n744_), .A3(new_n668_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1333gat));
  INV_X1    g547(.A(G71gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n741_), .B2(new_n395_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT49), .Z(new_n751_));
  NAND3_X1  g550(.A1(new_n736_), .A2(new_n749_), .A3(new_n395_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1334gat));
  NAND3_X1  g552(.A1(new_n736_), .A2(new_n367_), .A3(new_n375_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n741_), .A2(new_n375_), .ZN(new_n755_));
  XOR2_X1   g554(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(G78gat), .A3(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G78gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(G1335gat));
  NAND2_X1  g558(.A1(new_n739_), .A2(new_n649_), .ZN(new_n760_));
  NOR4_X1   g559(.A1(new_n459_), .A2(new_n760_), .A3(new_n589_), .A4(new_n660_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n481_), .A3(new_n422_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n760_), .A2(new_n589_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n696_), .A2(new_n763_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n764_), .A2(new_n422_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n762_), .B1(new_n765_), .B2(new_n481_), .ZN(G1336gat));
  NAND3_X1  g565(.A1(new_n761_), .A2(new_n482_), .A3(new_n668_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n764_), .A2(new_n668_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n482_), .ZN(G1337gat));
  NAND3_X1  g568(.A1(new_n761_), .A2(new_n485_), .A3(new_n395_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n764_), .A2(new_n395_), .ZN(new_n771_));
  INV_X1    g570(.A(G99gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT51), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT51), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n775_), .B(new_n770_), .C1(new_n771_), .C2(new_n772_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n761_), .A2(new_n369_), .A3(new_n375_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n696_), .A2(new_n375_), .A3(new_n763_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n779_), .A2(new_n780_), .A3(G106gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n780_), .B1(new_n779_), .B2(G106gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n778_), .B(new_n785_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  NAND3_X1  g586(.A1(new_n586_), .A2(new_n587_), .A3(new_n531_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n525_), .A2(KEYINPUT12), .A3(new_n508_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n789_), .A2(new_n527_), .A3(new_n522_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT55), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n524_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n527_), .B1(new_n789_), .B2(new_n522_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(KEYINPUT115), .A3(KEYINPUT55), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT55), .B(new_n465_), .C1(new_n518_), .C2(new_n523_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n792_), .A2(new_n794_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n463_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT56), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n463_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n788_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n572_), .A2(new_n563_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n566_), .A2(new_n563_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n584_), .B1(new_n805_), .B2(new_n560_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n585_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n585_), .A2(KEYINPUT116), .A3(new_n807_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n810_), .A2(new_n811_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n660_), .B1(new_n803_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(KEYINPUT57), .B(new_n660_), .C1(new_n803_), .C2(new_n812_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n534_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n817_));
  AND3_X1   g616(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n463_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n463_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n817_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT58), .B(new_n817_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n633_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n815_), .A2(new_n816_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n649_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n740_), .A2(new_n535_), .A3(new_n532_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT114), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n827_), .B(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(KEYINPUT54), .B1(new_n829_), .B2(new_n633_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n827_), .B(KEYINPUT114), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n832_), .A3(new_n692_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n830_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n826_), .A2(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n377_), .A2(new_n394_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n422_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(G113gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n589_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n837_), .A2(new_n841_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n825_), .A2(new_n649_), .B1(new_n830_), .B2(new_n833_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n843_), .A2(new_n423_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(KEYINPUT59), .A3(new_n836_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n588_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n840_), .B1(new_n846_), .B2(new_n839_), .ZN(G1340gat));
  AOI21_X1  g646(.A(new_n540_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n848_));
  INV_X1    g647(.A(G120gat), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT117), .B1(new_n849_), .B2(KEYINPUT60), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT60), .ZN(new_n851_));
  AOI21_X1  g650(.A(G120gat), .B1(new_n739_), .B2(new_n851_), .ZN(new_n852_));
  MUX2_X1   g651(.A(new_n850_), .B(KEYINPUT117), .S(new_n852_), .Z(new_n853_));
  OAI22_X1  g652(.A1(new_n848_), .A2(new_n849_), .B1(new_n837_), .B2(new_n853_), .ZN(G1341gat));
  AOI21_X1  g653(.A(G127gat), .B1(new_n838_), .B2(new_n662_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n842_), .A2(new_n845_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n662_), .A2(G127gat), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT118), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n855_), .B1(new_n856_), .B2(new_n858_), .ZN(G1342gat));
  INV_X1    g658(.A(G134gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n837_), .B2(new_n660_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(KEYINPUT119), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n863_), .B(new_n860_), .C1(new_n837_), .C2(new_n660_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n692_), .A2(new_n860_), .ZN(new_n865_));
  AOI22_X1  g664(.A1(new_n862_), .A2(new_n864_), .B1(new_n856_), .B2(new_n865_), .ZN(G1343gat));
  NOR3_X1   g665(.A1(new_n668_), .A2(new_n376_), .A3(new_n395_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n844_), .A2(new_n589_), .A3(new_n867_), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT120), .B(G141gat), .Z(new_n869_));
  XNOR2_X1  g668(.A(new_n868_), .B(new_n869_), .ZN(G1344gat));
  NAND3_X1  g669(.A1(new_n844_), .A2(new_n739_), .A3(new_n867_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g671(.A1(new_n844_), .A2(new_n662_), .A3(new_n867_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  NOR2_X1   g674(.A1(new_n660_), .A2(G162gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n844_), .A2(new_n867_), .A3(new_n876_), .ZN(new_n877_));
  AND4_X1   g676(.A1(new_n633_), .A2(new_n835_), .A3(new_n422_), .A4(new_n867_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n332_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n879_), .A2(new_n880_), .ZN(new_n881_));
  OAI211_X1 g680(.A(KEYINPUT121), .B(new_n877_), .C1(new_n878_), .C2(new_n332_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1347gat));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n424_), .A2(new_n325_), .A3(new_n375_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n843_), .A2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n589_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n884_), .B1(new_n888_), .B2(G169gat), .ZN(new_n889_));
  AOI211_X1 g688(.A(KEYINPUT62), .B(new_n253_), .C1(new_n887_), .C2(new_n589_), .ZN(new_n890_));
  AOI21_X1  g689(.A(KEYINPUT122), .B1(new_n835_), .B2(new_n885_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n843_), .A2(new_n892_), .A3(new_n886_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n891_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n589_), .A2(new_n281_), .ZN(new_n895_));
  OAI22_X1  g694(.A1(new_n889_), .A2(new_n890_), .B1(new_n894_), .B2(new_n895_), .ZN(G1348gat));
  NAND2_X1  g695(.A1(new_n835_), .A2(new_n885_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n897_), .A2(new_n254_), .A3(new_n540_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n739_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n900_), .A3(new_n241_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n835_), .A2(KEYINPUT122), .A3(new_n885_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n892_), .B1(new_n843_), .B2(new_n886_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n540_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(KEYINPUT123), .B1(new_n904_), .B2(new_n242_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n898_), .B1(new_n901_), .B2(new_n905_), .ZN(G1349gat));
  OR2_X1    g705(.A1(new_n649_), .A2(new_n264_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n907_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n897_), .A2(new_n649_), .ZN(new_n909_));
  OAI22_X1  g708(.A1(new_n908_), .A2(KEYINPUT124), .B1(G183gat), .B2(new_n909_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n908_), .A2(KEYINPUT124), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1350gat));
  OAI21_X1  g711(.A(G190gat), .B1(new_n894_), .B2(new_n692_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n265_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n660_), .A2(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n913_), .B1(new_n894_), .B2(new_n915_), .ZN(G1351gat));
  NOR3_X1   g715(.A1(new_n395_), .A2(new_n376_), .A3(new_n422_), .ZN(new_n917_));
  AND2_X1   g716(.A1(new_n917_), .A2(KEYINPUT125), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(KEYINPUT125), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n918_), .A2(new_n919_), .A3(new_n325_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n835_), .A2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n588_), .ZN(new_n922_));
  XOR2_X1   g721(.A(KEYINPUT126), .B(G197gat), .Z(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1352gat));
  INV_X1    g723(.A(new_n921_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n739_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n921_), .A2(new_n649_), .ZN(new_n929_));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n930_));
  INV_X1    g729(.A(G211gat), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n928_), .B1(new_n929_), .B2(new_n932_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  OAI211_X1 g733(.A(KEYINPUT127), .B(new_n934_), .C1(new_n921_), .C2(new_n649_), .ZN(new_n935_));
  XOR2_X1   g734(.A(KEYINPUT63), .B(G211gat), .Z(new_n936_));
  AOI22_X1  g735(.A1(new_n933_), .A2(new_n935_), .B1(new_n929_), .B2(new_n936_), .ZN(G1354gat));
  OAI21_X1  g736(.A(G218gat), .B1(new_n921_), .B2(new_n692_), .ZN(new_n938_));
  OR2_X1    g737(.A1(new_n660_), .A2(G218gat), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n921_), .B2(new_n939_), .ZN(G1355gat));
endmodule


