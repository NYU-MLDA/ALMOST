//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:29 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n836_, new_n837_,
    new_n838_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n907_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_;
  XNOR2_X1  g000(.A(G120gat), .B(G148gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT5), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G176gat), .B(G204gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  XOR2_X1   g004(.A(new_n205_), .B(KEYINPUT72), .Z(new_n206_));
  NAND4_X1  g005(.A1(KEYINPUT66), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT10), .B(G99gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n208_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G85gat), .B(G92gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT9), .ZN(new_n214_));
  AOI21_X1  g013(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n215_), .A2(KEYINPUT66), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G99gat), .A2(G106gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT6), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n212_), .A2(new_n217_), .A3(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G57gat), .B(G64gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT11), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G71gat), .B(G78gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n222_), .A2(new_n224_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n221_), .A2(KEYINPUT11), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n226_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT70), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n219_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT6), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n218_), .B(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT70), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G99gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n237_), .A2(new_n211_), .A3(KEYINPUT67), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n239_), .B1(G99gat), .B2(G106gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT7), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n238_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n237_), .A2(new_n211_), .ZN(new_n244_));
  AOI21_X1  g043(.A(new_n243_), .B1(new_n244_), .B2(KEYINPUT7), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n238_), .A2(new_n240_), .A3(new_n243_), .A4(new_n241_), .ZN(new_n248_));
  AND3_X1   g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n247_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n236_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n213_), .B(KEYINPUT69), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n230_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(G99gat), .A2(G106gat), .ZN(new_n254_));
  OAI21_X1  g053(.A(KEYINPUT68), .B1(new_n254_), .B2(new_n241_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT7), .B1(new_n244_), .B2(new_n239_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n255_), .B1(new_n256_), .B2(new_n238_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n248_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n219_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(new_n230_), .A3(new_n252_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n220_), .B(new_n229_), .C1(new_n253_), .C2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G230gat), .A2(G233gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n262_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n220_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n232_), .A2(new_n235_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT71), .B1(new_n257_), .B2(new_n258_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n269_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n252_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT8), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n268_), .B1(new_n274_), .B2(new_n260_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT12), .B1(new_n275_), .B2(new_n229_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n220_), .B1(new_n253_), .B2(new_n261_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT12), .ZN(new_n278_));
  INV_X1    g077(.A(new_n229_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n277_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n267_), .B1(new_n276_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n279_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n266_), .B1(new_n282_), .B2(new_n262_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n206_), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT73), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n276_), .A2(new_n280_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n267_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n282_), .A2(new_n262_), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n286_), .A2(new_n287_), .B1(new_n288_), .B2(new_n265_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n205_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n285_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NOR4_X1   g090(.A1(new_n281_), .A2(new_n283_), .A3(KEYINPUT73), .A4(new_n205_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n284_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT13), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  OAI211_X1 g094(.A(KEYINPUT13), .B(new_n284_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n298_), .A2(KEYINPUT74), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(KEYINPUT74), .ZN(new_n300_));
  AND2_X1   g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT98), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n304_), .A2(KEYINPUT1), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n304_), .B1(new_n306_), .B2(KEYINPUT1), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT87), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n305_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n309_), .B1(new_n308_), .B2(new_n307_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT88), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT88), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n310_), .A2(new_n317_), .A3(new_n314_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n306_), .ZN(new_n320_));
  XOR2_X1   g119(.A(new_n313_), .B(KEYINPUT3), .Z(new_n321_));
  XOR2_X1   g120(.A(new_n311_), .B(KEYINPUT2), .Z(new_n322_));
  OAI211_X1 g121(.A(new_n304_), .B(new_n320_), .C1(new_n321_), .C2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G127gat), .B(G134gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G113gat), .B(G120gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  OR2_X1    g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(new_n327_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(KEYINPUT4), .A3(new_n329_), .ZN(new_n330_));
  OR2_X1    g129(.A1(new_n329_), .A2(KEYINPUT4), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G1gat), .B(G29gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G85gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT0), .B(G57gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n334_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n335_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n333_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n339_), .B1(new_n344_), .B2(new_n341_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT97), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G183gat), .A2(G190gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT23), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n350_), .B1(G183gat), .B2(G190gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G169gat), .A2(G176gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(KEYINPUT22), .B(G169gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n353_), .A2(KEYINPUT84), .ZN(new_n354_));
  INV_X1    g153(.A(G176gat), .ZN(new_n355_));
  INV_X1    g154(.A(G169gat), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n356_), .A2(KEYINPUT22), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT84), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n355_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n351_), .B(new_n352_), .C1(new_n354_), .C2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT25), .B(G183gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT26), .B(G190gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n356_), .A2(new_n355_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n364_), .A2(KEYINPUT24), .A3(new_n352_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT83), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n363_), .A2(KEYINPUT82), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(KEYINPUT82), .B2(new_n363_), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n364_), .A2(KEYINPUT24), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n350_), .A2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n370_), .B1(new_n366_), .B2(new_n365_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n360_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G197gat), .B(G204gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT89), .ZN(new_n374_));
  INV_X1    g173(.A(G197gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(G204gat), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n374_), .B(KEYINPUT21), .C1(KEYINPUT89), .C2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT21), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n373_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G211gat), .B(G218gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n377_), .A2(new_n379_), .A3(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(KEYINPUT90), .ZN(new_n382_));
  INV_X1    g181(.A(new_n373_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(KEYINPUT21), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n381_), .A2(new_n384_), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n372_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n353_), .A2(new_n355_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n351_), .A2(new_n352_), .A3(new_n387_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n388_), .A2(KEYINPUT93), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(KEYINPUT93), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n365_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n392_), .A2(KEYINPUT92), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n370_), .B1(new_n392_), .B2(KEYINPUT92), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n391_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n385_), .ZN(new_n397_));
  OAI211_X1 g196(.A(KEYINPUT20), .B(new_n386_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G226gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n399_), .B(KEYINPUT19), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(G8gat), .B(G36gat), .Z(new_n402_));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n396_), .A2(new_n397_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n400_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT20), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n409_), .B1(new_n372_), .B2(new_n385_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n407_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n401_), .A2(new_n406_), .A3(new_n411_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n412_), .A2(KEYINPUT27), .ZN(new_n413_));
  OAI21_X1  g212(.A(KEYINPUT96), .B1(new_n398_), .B2(new_n400_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n395_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(new_n390_), .A3(new_n389_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n409_), .B1(new_n416_), .B2(new_n385_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT96), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(new_n408_), .A4(new_n386_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n415_), .A2(new_n397_), .A3(new_n388_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n410_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n400_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n414_), .A2(new_n419_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n406_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n408_), .B1(new_n417_), .B2(new_n386_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n407_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n424_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n412_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT27), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n413_), .A2(new_n425_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n343_), .A2(KEYINPUT97), .A3(new_n345_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n348_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT86), .B(KEYINPUT31), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n327_), .B(new_n435_), .Z(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  XOR2_X1   g236(.A(G71gat), .B(G99gat), .Z(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(G43gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G227gat), .A2(G233gat), .ZN(new_n440_));
  INV_X1    g239(.A(G15gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n439_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT85), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT30), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n372_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n372_), .A2(new_n445_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n444_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n446_), .A2(new_n444_), .A3(new_n447_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n443_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n450_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n443_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n437_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n453_), .B1(new_n452_), .B2(new_n448_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n456_), .B(new_n436_), .C1(new_n452_), .C2(new_n453_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G78gat), .B(G106gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n461_), .A2(KEYINPUT91), .ZN(new_n462_));
  INV_X1    g261(.A(new_n324_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT28), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT29), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT28), .B1(new_n324_), .B2(KEYINPUT29), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G22gat), .B(G50gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n466_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n469_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n462_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n385_), .B1(new_n463_), .B2(new_n465_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G228gat), .A2(G233gat), .ZN(new_n475_));
  XOR2_X1   g274(.A(new_n474_), .B(new_n475_), .Z(new_n476_));
  NAND2_X1  g275(.A1(new_n466_), .A2(new_n467_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(new_n468_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n478_), .A2(new_n461_), .A3(new_n470_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n473_), .A2(new_n476_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n476_), .B1(new_n473_), .B2(new_n479_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n459_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n474_), .B(new_n475_), .ZN(new_n484_));
  NOR3_X1   g283(.A1(new_n471_), .A2(new_n460_), .A3(new_n472_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n462_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n486_), .B1(new_n478_), .B2(new_n470_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n484_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n488_), .A2(new_n458_), .A3(new_n480_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n483_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n406_), .A2(KEYINPUT32), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n401_), .A2(new_n411_), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n491_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n423_), .A2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n346_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(KEYINPUT95), .A2(KEYINPUT33), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n345_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n496_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n339_), .B(new_n498_), .C1(new_n344_), .C2(new_n341_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n328_), .A2(new_n329_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n339_), .B1(new_n500_), .B2(new_n334_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n501_), .B1(new_n334_), .B2(new_n332_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n499_), .A2(new_n502_), .A3(new_n412_), .A4(new_n428_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n495_), .B1(new_n497_), .B2(new_n503_), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n481_), .A2(new_n482_), .A3(new_n458_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n434_), .A2(new_n490_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G29gat), .B(G36gat), .Z(new_n507_));
  XOR2_X1   g306(.A(G43gat), .B(G50gat), .Z(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  XOR2_X1   g308(.A(new_n509_), .B(KEYINPUT15), .Z(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT78), .B(G1gat), .ZN(new_n511_));
  INV_X1    g310(.A(G8gat), .ZN(new_n512_));
  OAI21_X1  g311(.A(KEYINPUT14), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G1gat), .B(G8gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n515_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(new_n514_), .A3(new_n516_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n510_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n509_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n520_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G229gat), .A2(G233gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n522_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n521_), .A2(new_n509_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n524_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n528_), .B(KEYINPUT81), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n526_), .B1(new_n529_), .B2(new_n525_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G113gat), .B(G141gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G169gat), .B(G197gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n526_), .B(new_n533_), .C1(new_n529_), .C2(new_n525_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n303_), .B1(new_n506_), .B2(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n503_), .A2(new_n497_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n494_), .A2(new_n492_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n505_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n489_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n458_), .B1(new_n488_), .B2(new_n480_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n543_), .B1(new_n546_), .B2(new_n433_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n547_), .A2(KEYINPUT98), .A3(new_n537_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n539_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G190gat), .B(G218gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G134gat), .B(G162gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n552_), .B(KEYINPUT36), .Z(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n509_), .B(new_n220_), .C1(new_n253_), .C2(new_n261_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n555_), .B1(new_n275_), .B2(new_n510_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT75), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XOR2_X1   g358(.A(new_n559_), .B(KEYINPUT34), .Z(new_n560_));
  NAND2_X1  g359(.A1(new_n558_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n560_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n556_), .A2(new_n557_), .A3(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(KEYINPUT35), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT35), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n556_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n510_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n277_), .A2(new_n568_), .ZN(new_n569_));
  AOI211_X1 g368(.A(KEYINPUT75), .B(new_n560_), .C1(new_n569_), .C2(new_n555_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n562_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n567_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n554_), .B1(new_n564_), .B2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT37), .B1(new_n573_), .B2(KEYINPUT76), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n552_), .A2(KEYINPUT36), .ZN(new_n575_));
  AND3_X1   g374(.A1(new_n564_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n576_), .A2(new_n573_), .A3(KEYINPUT77), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT77), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n570_), .A2(new_n571_), .A3(new_n565_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n566_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n553_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n564_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n578_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n574_), .B1(new_n577_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT37), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT76), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n585_), .B1(new_n581_), .B2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT77), .B1(new_n576_), .B2(new_n573_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n581_), .A2(new_n578_), .A3(new_n582_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n584_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT79), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n520_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(new_n229_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G127gat), .B(G155gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT16), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G183gat), .B(G211gat), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n598_), .B(new_n599_), .Z(new_n600_));
  INV_X1    g399(.A(KEYINPUT17), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n596_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n596_), .A2(KEYINPUT80), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n600_), .A2(new_n601_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n605_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n603_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n592_), .A2(new_n609_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n302_), .A2(new_n549_), .A3(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n348_), .A2(new_n432_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT38), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT99), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n611_), .A2(new_n613_), .A3(new_n511_), .A4(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n614_), .A2(KEYINPUT99), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n609_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n298_), .A2(new_n537_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n576_), .A2(new_n573_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n506_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n620_), .A2(new_n621_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n622_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n626_), .B2(new_n612_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n618_), .A2(new_n627_), .ZN(G1324gat));
  INV_X1    g427(.A(new_n431_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n611_), .A2(new_n512_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT39), .ZN(new_n631_));
  INV_X1    g430(.A(new_n626_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(new_n629_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n631_), .B1(new_n633_), .B2(G8gat), .ZN(new_n634_));
  AOI211_X1 g433(.A(KEYINPUT39), .B(new_n512_), .C1(new_n632_), .C2(new_n629_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n630_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n636_), .B(new_n637_), .Z(G1325gat));
  NAND3_X1  g437(.A1(new_n611_), .A2(new_n441_), .A3(new_n458_), .ZN(new_n639_));
  OAI21_X1  g438(.A(G15gat), .B1(new_n626_), .B2(new_n459_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT41), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n640_), .A2(new_n641_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n639_), .B1(new_n642_), .B2(new_n643_), .ZN(G1326gat));
  NOR2_X1   g443(.A1(new_n481_), .A2(new_n482_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT102), .Z(new_n646_));
  NOR2_X1   g445(.A1(new_n646_), .A2(G22gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT103), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n611_), .A2(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G22gat), .B1(new_n626_), .B2(new_n646_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n650_), .A2(KEYINPUT42), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(KEYINPUT42), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n649_), .B1(new_n651_), .B2(new_n652_), .ZN(G1327gat));
  INV_X1    g452(.A(new_n623_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(new_n619_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n298_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n656_), .B1(new_n539_), .B2(new_n548_), .ZN(new_n657_));
  INV_X1    g456(.A(G29gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(new_n658_), .A3(new_n613_), .ZN(new_n659_));
  OAI21_X1  g458(.A(KEYINPUT43), .B1(new_n591_), .B2(new_n506_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n547_), .A2(new_n661_), .A3(new_n590_), .A4(new_n584_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n297_), .A2(new_n538_), .A3(new_n619_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n663_), .A2(new_n664_), .A3(KEYINPUT44), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n669_), .A2(new_n613_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n659_), .B1(new_n670_), .B2(new_n658_), .ZN(G1328gat));
  NAND3_X1  g470(.A1(new_n667_), .A2(new_n629_), .A3(new_n668_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n667_), .A2(KEYINPUT104), .A3(new_n629_), .A4(new_n668_), .ZN(new_n675_));
  NAND4_X1  g474(.A1(new_n674_), .A2(KEYINPUT106), .A3(G36gat), .A4(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT45), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n431_), .A2(G36gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n657_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n678_), .B1(new_n657_), .B2(new_n679_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n677_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n682_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n684_), .A2(KEYINPUT45), .A3(new_n680_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n683_), .A2(new_n685_), .A3(KEYINPUT106), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT46), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n676_), .A2(new_n686_), .A3(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n687_), .B1(new_n676_), .B2(new_n686_), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1329gat));
  NAND2_X1  g489(.A1(new_n669_), .A2(new_n458_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n459_), .A2(G43gat), .ZN(new_n692_));
  AOI22_X1  g491(.A1(new_n691_), .A2(G43gat), .B1(new_n657_), .B2(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(G1330gat));
  INV_X1    g494(.A(new_n646_), .ZN(new_n696_));
  AOI21_X1  g495(.A(G50gat), .B1(new_n657_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n645_), .ZN(new_n698_));
  AND2_X1   g497(.A1(new_n698_), .A2(G50gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n697_), .B1(new_n669_), .B2(new_n699_), .ZN(G1331gat));
  NOR2_X1   g499(.A1(new_n609_), .A2(new_n537_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n506_), .A2(new_n623_), .A3(new_n702_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n301_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(G57gat), .B1(new_n705_), .B2(new_n612_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n506_), .A2(new_n537_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n610_), .A2(new_n297_), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(G57gat), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n613_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n706_), .A2(new_n710_), .ZN(G1332gat));
  INV_X1    g510(.A(G64gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n704_), .B2(new_n629_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT48), .Z(new_n714_));
  NAND3_X1  g513(.A1(new_n708_), .A2(new_n712_), .A3(new_n629_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1333gat));
  INV_X1    g515(.A(G71gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n717_), .B1(new_n704_), .B2(new_n458_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT108), .B(KEYINPUT49), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n708_), .A2(new_n717_), .A3(new_n458_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1334gat));
  INV_X1    g521(.A(G78gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n708_), .A2(new_n723_), .A3(new_n696_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n704_), .A2(new_n696_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(G78gat), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(KEYINPUT50), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(KEYINPUT50), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n724_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT109), .ZN(G1335gat));
  AND2_X1   g529(.A1(new_n707_), .A2(new_n655_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n731_), .A2(new_n301_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n613_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n297_), .A2(new_n538_), .A3(new_n609_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n613_), .A2(G85gat), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT110), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n734_), .B1(new_n736_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT111), .ZN(G1336gat));
  AND2_X1   g539(.A1(new_n736_), .A2(new_n629_), .ZN(new_n741_));
  INV_X1    g540(.A(G92gat), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n629_), .A2(new_n742_), .ZN(new_n743_));
  OAI22_X1  g542(.A1(new_n741_), .A2(new_n742_), .B1(new_n732_), .B2(new_n743_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT112), .Z(G1337gat));
  AOI21_X1  g544(.A(new_n237_), .B1(new_n736_), .B2(new_n458_), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n732_), .A2(new_n209_), .A3(new_n459_), .ZN(new_n747_));
  AOI211_X1 g546(.A(new_n746_), .B(new_n747_), .C1(KEYINPUT113), .C2(KEYINPUT51), .ZN(new_n748_));
  NOR2_X1   g547(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n748_), .B(new_n749_), .ZN(G1338gat));
  NAND3_X1  g549(.A1(new_n733_), .A2(new_n211_), .A3(new_n698_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT52), .ZN(new_n752_));
  OAI21_X1  g551(.A(G106gat), .B1(new_n752_), .B2(KEYINPUT114), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n736_), .B2(new_n698_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(KEYINPUT114), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT53), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n757_), .B(new_n758_), .ZN(G1339gat));
  NOR3_X1   g558(.A1(new_n612_), .A2(new_n489_), .A3(new_n629_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n295_), .A2(new_n296_), .A3(new_n701_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n762_), .B1(new_n591_), .B2(new_n764_), .ZN(new_n765_));
  AOI211_X1 g564(.A(KEYINPUT115), .B(new_n763_), .C1(new_n584_), .C2(new_n590_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n761_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n581_), .A2(new_n586_), .ZN(new_n769_));
  AOI22_X1  g568(.A1(new_n588_), .A2(new_n589_), .B1(new_n769_), .B2(KEYINPUT37), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n764_), .B1(new_n768_), .B2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(KEYINPUT115), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n591_), .A2(new_n762_), .A3(new_n764_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n772_), .A2(KEYINPUT54), .A3(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n767_), .A2(new_n774_), .ZN(new_n775_));
  XOR2_X1   g574(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n776_));
  NOR2_X1   g575(.A1(new_n291_), .A2(new_n292_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(new_n538_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n275_), .A2(KEYINPUT12), .A3(new_n229_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n278_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n287_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT116), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT116), .B1(new_n281_), .B2(KEYINPUT55), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n281_), .A2(KEYINPUT55), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n262_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n265_), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n784_), .A2(new_n785_), .A3(new_n786_), .A4(new_n788_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n206_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT56), .B1(new_n789_), .B2(new_n206_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n778_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n525_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n522_), .A2(new_n524_), .A3(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n534_), .B(new_n794_), .C1(new_n529_), .C2(new_n793_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n536_), .A2(new_n795_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT117), .Z(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n293_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n792_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n776_), .B1(new_n799_), .B2(new_n654_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n801_));
  AOI211_X1 g600(.A(new_n801_), .B(new_n623_), .C1(new_n792_), .C2(new_n798_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n800_), .A2(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n790_), .A2(new_n791_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n796_), .B(KEYINPUT117), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n805_), .A2(new_n777_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  OR3_X1    g606(.A1(new_n804_), .A2(new_n806_), .A3(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n807_), .B1(new_n804_), .B2(new_n806_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n592_), .A2(new_n808_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n619_), .B1(new_n803_), .B2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n760_), .B1(new_n775_), .B2(new_n811_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n812_), .A2(G113gat), .A3(new_n538_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT59), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n812_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT59), .B(new_n760_), .C1(new_n775_), .C2(new_n811_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n538_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(G113gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n814_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(KEYINPUT119), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n822_), .B(new_n814_), .C1(new_n818_), .C2(new_n819_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1340gat));
  INV_X1    g623(.A(new_n812_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n298_), .A2(KEYINPUT60), .ZN(new_n826_));
  INV_X1    g625(.A(G120gat), .ZN(new_n827_));
  MUX2_X1   g626(.A(KEYINPUT60), .B(new_n826_), .S(new_n827_), .Z(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n302_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n827_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT120), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n829_), .B(new_n833_), .C1(new_n830_), .C2(new_n827_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(G1341gat));
  INV_X1    g634(.A(G127gat), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n825_), .A2(new_n836_), .A3(new_n619_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n609_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n837_), .B1(new_n838_), .B2(new_n836_), .ZN(G1342gat));
  INV_X1    g638(.A(G134gat), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n825_), .A2(new_n840_), .A3(new_n623_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n591_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n840_), .ZN(G1343gat));
  NOR2_X1   g642(.A1(new_n612_), .A2(new_n629_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n545_), .B(new_n844_), .C1(new_n775_), .C2(new_n811_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n845_), .B(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(new_n537_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G141gat), .ZN(new_n849_));
  INV_X1    g648(.A(G141gat), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n847_), .A2(new_n850_), .A3(new_n537_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1344gat));
  NAND2_X1  g651(.A1(new_n847_), .A2(new_n301_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(G148gat), .ZN(new_n854_));
  INV_X1    g653(.A(G148gat), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n847_), .A2(new_n855_), .A3(new_n301_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n856_), .ZN(G1345gat));
  NAND2_X1  g656(.A1(new_n847_), .A2(new_n619_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(KEYINPUT61), .B(G155gat), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n859_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n847_), .A2(new_n619_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1346gat));
  INV_X1    g662(.A(G162gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n847_), .A2(new_n864_), .A3(new_n623_), .ZN(new_n865_));
  OR2_X1    g664(.A1(new_n845_), .A2(new_n846_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n845_), .A2(new_n846_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n591_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n865_), .B1(new_n864_), .B2(new_n868_), .ZN(G1347gat));
  NOR2_X1   g668(.A1(new_n613_), .A2(new_n431_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n458_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n537_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(KEYINPUT122), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n874_), .A2(new_n696_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n775_), .A2(new_n811_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n356_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT62), .ZN(new_n878_));
  AND2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n877_), .A2(new_n878_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n871_), .A2(new_n696_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n876_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(KEYINPUT123), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT123), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n876_), .A2(new_n884_), .A3(new_n881_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n537_), .A2(new_n353_), .ZN(new_n887_));
  OAI22_X1  g686(.A1(new_n879_), .A2(new_n880_), .B1(new_n886_), .B2(new_n887_), .ZN(G1348gat));
  NAND2_X1  g687(.A1(new_n876_), .A2(new_n645_), .ZN(new_n889_));
  NOR4_X1   g688(.A1(new_n889_), .A2(new_n355_), .A3(new_n302_), .A4(new_n871_), .ZN(new_n890_));
  INV_X1    g689(.A(new_n885_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n884_), .B1(new_n876_), .B2(new_n881_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n297_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n890_), .B1(new_n894_), .B2(new_n355_), .ZN(G1349gat));
  NOR2_X1   g694(.A1(new_n609_), .A2(new_n361_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n876_), .A2(new_n619_), .A3(new_n645_), .A4(new_n872_), .ZN(new_n897_));
  OR2_X1    g696(.A1(new_n897_), .A2(KEYINPUT124), .ZN(new_n898_));
  AOI21_X1  g697(.A(G183gat), .B1(new_n897_), .B2(KEYINPUT124), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n893_), .A2(new_n896_), .B1(new_n898_), .B2(new_n899_), .ZN(G1350gat));
  NAND3_X1  g699(.A1(new_n893_), .A2(new_n623_), .A3(new_n362_), .ZN(new_n901_));
  OAI21_X1  g700(.A(G190gat), .B1(new_n886_), .B2(new_n591_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(G1351gat));
  AND2_X1   g702(.A1(new_n876_), .A2(new_n545_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n904_), .A2(new_n537_), .A3(new_n870_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g705(.A1(new_n904_), .A2(new_n301_), .A3(new_n870_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g707(.A(new_n609_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n876_), .A2(new_n545_), .A3(new_n870_), .A4(new_n909_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n910_), .A2(KEYINPUT125), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(KEYINPUT125), .ZN(new_n912_));
  OAI22_X1  g711(.A1(new_n911_), .A2(new_n912_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n910_), .A2(KEYINPUT125), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n910_), .A2(KEYINPUT125), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n913_), .A2(new_n917_), .ZN(G1354gat));
  NAND4_X1  g717(.A1(new_n876_), .A2(new_n623_), .A3(new_n545_), .A4(new_n870_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(KEYINPUT126), .ZN(new_n920_));
  XOR2_X1   g719(.A(KEYINPUT127), .B(G218gat), .Z(new_n921_));
  AND2_X1   g720(.A1(new_n904_), .A2(new_n870_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n591_), .A2(new_n921_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n920_), .A2(new_n921_), .B1(new_n922_), .B2(new_n923_), .ZN(G1355gat));
endmodule


