//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n861_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT21), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  OR2_X1    g003(.A1(G197gat), .A2(G204gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n205_), .A2(KEYINPUT21), .A3(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n204_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n207_), .A2(new_n208_), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G233gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(KEYINPUT93), .A2(G228gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n213_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G155gat), .A2(G162gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G141gat), .ZN(new_n224_));
  INV_X1    g023(.A(G148gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(KEYINPUT3), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n227_), .B1(G141gat), .B2(G148gat), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n226_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G141gat), .A2(G148gat), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT2), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT92), .B1(new_n229_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n226_), .A2(new_n228_), .ZN(new_n236_));
  AND3_X1   g035(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT92), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n236_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n223_), .B1(new_n235_), .B2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n221_), .B1(KEYINPUT1), .B2(new_n219_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n243_), .B1(KEYINPUT1), .B2(new_n219_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(G141gat), .A2(G148gat), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n244_), .A2(new_n246_), .A3(new_n230_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n242_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT29), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n212_), .B(new_n218_), .C1(new_n248_), .C2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(new_n242_), .B2(new_n247_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(new_n212_), .ZN(new_n253_));
  AOI21_X1  g052(.A(KEYINPUT95), .B1(new_n253_), .B2(new_n217_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT95), .ZN(new_n255_));
  AOI211_X1 g054(.A(new_n255_), .B(new_n218_), .C1(new_n252_), .C2(new_n212_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n250_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G78gat), .B(G106gat), .Z(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n258_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n260_), .B(new_n250_), .C1(new_n254_), .C2(new_n256_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT28), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n248_), .A2(new_n263_), .A3(new_n249_), .ZN(new_n264_));
  AND3_X1   g063(.A1(new_n236_), .A2(new_n239_), .A3(new_n240_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n240_), .B1(new_n236_), .B2(new_n239_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n222_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n244_), .A2(new_n246_), .A3(new_n230_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT28), .B1(new_n269_), .B2(KEYINPUT29), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G22gat), .B(G50gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n264_), .A2(new_n270_), .A3(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n272_), .B1(new_n264_), .B2(new_n270_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n262_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n259_), .A2(new_n275_), .A3(new_n261_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT27), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G226gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT19), .ZN(new_n283_));
  INV_X1    g082(.A(G169gat), .ZN(new_n284_));
  INV_X1    g083(.A(G176gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT84), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(KEYINPUT24), .A4(new_n288_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n286_), .A2(KEYINPUT24), .A3(new_n288_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT84), .B1(new_n286_), .B2(KEYINPUT24), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(KEYINPUT83), .A2(G190gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT26), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT25), .ZN(new_n296_));
  OR2_X1    g095(.A1(KEYINPUT82), .A2(G183gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(KEYINPUT82), .A2(G183gat), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n296_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n295_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(G183gat), .A2(G190gat), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT85), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT85), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT23), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n302_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT86), .ZN(new_n308_));
  INV_X1    g107(.A(new_n302_), .ZN(new_n309_));
  OAI22_X1  g108(.A1(new_n307_), .A2(new_n308_), .B1(KEYINPUT23), .B2(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT85), .B(KEYINPUT23), .ZN(new_n311_));
  NOR3_X1   g110(.A1(new_n311_), .A2(KEYINPUT86), .A3(new_n302_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n292_), .B(new_n301_), .C1(new_n310_), .C2(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(KEYINPUT87), .A2(G169gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(KEYINPUT87), .A2(G169gat), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT22), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT88), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT88), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n318_), .B(KEYINPUT22), .C1(new_n314_), .C2(new_n315_), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT89), .B1(new_n284_), .B2(KEYINPUT22), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT89), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT22), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(new_n322_), .A3(G169gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(G176gat), .B1(new_n320_), .B2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n317_), .A2(new_n319_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n309_), .A2(new_n303_), .ZN(new_n326_));
  INV_X1    g125(.A(G190gat), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n297_), .A2(new_n327_), .A3(new_n298_), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n326_), .B(new_n328_), .C1(new_n309_), .C2(new_n311_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n325_), .A2(new_n288_), .A3(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n313_), .A2(new_n330_), .A3(new_n211_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT96), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(KEYINPUT20), .ZN(new_n333_));
  XOR2_X1   g132(.A(KEYINPUT22), .B(G169gat), .Z(new_n334_));
  OAI21_X1  g133(.A(new_n288_), .B1(new_n334_), .B2(G176gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n307_), .A2(new_n308_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT86), .B1(new_n311_), .B2(new_n302_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n336_), .B(new_n337_), .C1(KEYINPUT23), .C2(new_n309_), .ZN(new_n338_));
  OR2_X1    g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n335_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n302_), .A2(KEYINPUT23), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n304_), .A2(new_n306_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n341_), .B1(new_n342_), .B2(new_n302_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n286_), .A2(new_n288_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT97), .B(KEYINPUT24), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT25), .B(G183gat), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT26), .B(G190gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NOR2_X1   g148(.A1(G169gat), .A2(G176gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n345_), .A2(new_n350_), .ZN(new_n351_));
  AND4_X1   g150(.A1(new_n343_), .A2(new_n346_), .A3(new_n349_), .A4(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n212_), .B1(new_n340_), .B2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n333_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n332_), .B1(new_n331_), .B2(KEYINPUT20), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n283_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n340_), .A2(new_n212_), .A3(new_n352_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n283_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n313_), .A2(new_n330_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n212_), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n358_), .A2(KEYINPUT20), .A3(new_n359_), .A4(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G8gat), .B(G36gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT18), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G64gat), .B(G92gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n363_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n356_), .A2(new_n367_), .A3(new_n362_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n370_), .A2(KEYINPUT27), .ZN(new_n372_));
  XOR2_X1   g171(.A(KEYINPUT102), .B(KEYINPUT20), .Z(new_n373_));
  INV_X1    g172(.A(new_n300_), .ZN(new_n374_));
  AND2_X1   g173(.A1(new_n297_), .A2(new_n298_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n374_), .B1(new_n375_), .B2(new_n296_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT24), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n287_), .B1(new_n350_), .B2(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n378_), .B1(new_n344_), .B2(new_n377_), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n376_), .A2(new_n295_), .B1(new_n379_), .B2(new_n289_), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n343_), .A2(new_n328_), .B1(G169gat), .B2(G176gat), .ZN(new_n381_));
  AOI22_X1  g180(.A1(new_n380_), .A2(new_n338_), .B1(new_n381_), .B2(new_n325_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n373_), .B1(new_n382_), .B2(new_n211_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n283_), .B1(new_n383_), .B2(new_n357_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT103), .ZN(new_n385_));
  INV_X1    g184(.A(new_n355_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n386_), .A2(new_n359_), .A3(new_n353_), .A4(new_n333_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT103), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n388_), .B(new_n283_), .C1(new_n383_), .C2(new_n357_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n385_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n368_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n281_), .A2(new_n371_), .B1(new_n372_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n280_), .A2(new_n392_), .ZN(new_n393_));
  XOR2_X1   g192(.A(G127gat), .B(G134gat), .Z(new_n394_));
  XOR2_X1   g193(.A(G113gat), .B(G120gat), .Z(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n397_), .B1(new_n242_), .B2(new_n247_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT98), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n267_), .A2(new_n396_), .A3(new_n268_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n398_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n269_), .A2(KEYINPUT98), .A3(new_n397_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT4), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n269_), .A2(new_n405_), .A3(new_n397_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G225gat), .A2(G233gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  AND2_X1   g207(.A1(new_n406_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n404_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT100), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n411_), .B1(new_n403_), .B2(new_n407_), .ZN(new_n412_));
  AOI211_X1 g211(.A(KEYINPUT100), .B(new_n408_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n410_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G57gat), .B(G85gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n414_), .A2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n410_), .B(new_n419_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G227gat), .A2(G233gat), .ZN(new_n424_));
  INV_X1    g223(.A(G71gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(G99gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n360_), .B(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(new_n397_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G15gat), .B(G43gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT90), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT30), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(KEYINPUT31), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n429_), .B(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n393_), .A2(new_n423_), .A3(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n434_), .B(KEYINPUT91), .ZN(new_n437_));
  AND3_X1   g236(.A1(new_n259_), .A2(new_n275_), .A3(new_n261_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n275_), .B1(new_n259_), .B2(new_n261_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n421_), .B(new_n422_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n372_), .A2(new_n391_), .ZN(new_n441_));
  AND3_X1   g240(.A1(new_n356_), .A2(new_n367_), .A3(new_n362_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n367_), .B1(new_n356_), .B2(new_n362_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n281_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT105), .B1(new_n440_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n423_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT105), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n392_), .A2(new_n447_), .A3(new_n448_), .A4(new_n279_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n367_), .A2(KEYINPUT32), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n356_), .A2(new_n362_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n450_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n452_), .B2(new_n390_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n423_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n422_), .A2(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n442_), .A2(new_n443_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n404_), .A2(KEYINPUT101), .A3(new_n407_), .A4(new_n406_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT101), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n405_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n406_), .A2(new_n407_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n459_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n419_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n458_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n420_), .A2(new_n455_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n410_), .B(new_n465_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n466_));
  NAND4_X1  g265(.A1(new_n456_), .A2(new_n457_), .A3(new_n464_), .A4(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n279_), .B1(new_n454_), .B2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT104), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n446_), .B(new_n449_), .C1(new_n468_), .C2(new_n469_), .ZN(new_n470_));
  AND4_X1   g269(.A1(new_n464_), .A2(new_n466_), .A3(new_n370_), .A4(new_n369_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n471_), .A2(new_n456_), .B1(new_n423_), .B2(new_n453_), .ZN(new_n472_));
  NOR3_X1   g271(.A1(new_n472_), .A2(KEYINPUT104), .A3(new_n279_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n437_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT106), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OAI211_X1 g275(.A(KEYINPUT106), .B(new_n437_), .C1(new_n470_), .C2(new_n473_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n436_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G29gat), .B(G36gat), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n479_), .A2(KEYINPUT75), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(KEYINPUT75), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G43gat), .B(G50gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(new_n484_), .B(KEYINPUT15), .Z(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT76), .B(G15gat), .ZN(new_n486_));
  INV_X1    g285(.A(G22gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT77), .B(G8gat), .ZN(new_n489_));
  INV_X1    g288(.A(G1gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT14), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G1gat), .B(G8gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT78), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n492_), .A2(new_n494_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n485_), .A2(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n497_), .A2(new_n484_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G229gat), .A2(G233gat), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n497_), .A2(new_n484_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n500_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(G113gat), .B(G141gat), .Z(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT81), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G169gat), .B(G197gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n506_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n501_), .A2(new_n505_), .A3(new_n510_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G230gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT64), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT7), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT67), .ZN(new_n519_));
  NOR2_X1   g318(.A1(G99gat), .A2(G106gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G99gat), .A2(G106gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT6), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n521_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT8), .ZN(new_n525_));
  XOR2_X1   g324(.A(G85gat), .B(G92gat), .Z(new_n526_));
  NAND3_X1  g325(.A1(new_n524_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT6), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT68), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT68), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT6), .ZN(new_n531_));
  AND3_X1   g330(.A1(new_n529_), .A2(new_n531_), .A3(new_n522_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n522_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT69), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n522_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n530_), .A2(KEYINPUT6), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n528_), .A2(KEYINPUT68), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n535_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT69), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n529_), .A2(new_n531_), .A3(new_n522_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n534_), .A2(new_n541_), .A3(new_n521_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT70), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n526_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT8), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n543_), .B1(new_n542_), .B2(new_n526_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n527_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  XOR2_X1   g346(.A(KEYINPUT10), .B(G99gat), .Z(new_n548_));
  INV_X1    g347(.A(G106gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT65), .ZN(new_n551_));
  XOR2_X1   g350(.A(KEYINPUT66), .B(G85gat), .Z(new_n552_));
  INV_X1    g351(.A(G92gat), .ZN(new_n553_));
  OR3_X1    g352(.A1(new_n552_), .A2(KEYINPUT9), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n526_), .A2(KEYINPUT9), .ZN(new_n555_));
  NAND4_X1  g354(.A1(new_n551_), .A2(new_n523_), .A3(new_n554_), .A4(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n557_), .A2(KEYINPUT11), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(KEYINPUT11), .ZN(new_n559_));
  XOR2_X1   g358(.A(G71gat), .B(G78gat), .Z(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n559_), .A2(new_n560_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n547_), .A2(new_n556_), .A3(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n547_), .B2(new_n556_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT71), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n565_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n566_), .A2(KEYINPUT71), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n517_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n517_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n567_), .A2(KEYINPUT12), .A3(new_n564_), .ZN(new_n573_));
  AOI211_X1 g372(.A(KEYINPUT12), .B(new_n563_), .C1(new_n547_), .C2(new_n556_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n572_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n571_), .A2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G120gat), .B(G148gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(G176gat), .B(G204gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n580_), .B(new_n581_), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n577_), .A2(new_n583_), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n571_), .A2(new_n576_), .A3(new_n582_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT13), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT13), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n588_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n547_), .A2(new_n556_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n591_), .A2(new_n484_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n485_), .A2(new_n591_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G232gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(KEYINPUT74), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  OR2_X1    g396(.A1(new_n597_), .A2(KEYINPUT35), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n592_), .A2(new_n593_), .A3(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(KEYINPUT35), .A3(new_n597_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n597_), .A2(KEYINPUT35), .ZN(new_n601_));
  NAND4_X1  g400(.A1(new_n592_), .A2(new_n601_), .A3(new_n593_), .A4(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT36), .Z(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n606_), .A2(KEYINPUT36), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n600_), .A2(new_n609_), .A3(new_n602_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n611_), .A2(KEYINPUT37), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT37), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n608_), .A2(new_n613_), .A3(new_n610_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n497_), .A2(G231gat), .A3(G233gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n495_), .A2(new_n496_), .A3(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n563_), .B(KEYINPUT79), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n616_), .A2(new_n620_), .A3(new_n618_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G127gat), .B(G155gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT16), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G183gat), .B(G211gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT17), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n628_), .A2(KEYINPUT17), .ZN(new_n631_));
  OR3_X1    g430(.A1(new_n624_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT80), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n624_), .B2(new_n630_), .ZN(new_n634_));
  AOI211_X1 g433(.A(KEYINPUT80), .B(new_n629_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n632_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n615_), .A2(new_n637_), .ZN(new_n638_));
  NOR4_X1   g437(.A1(new_n478_), .A2(new_n515_), .A3(new_n590_), .A4(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n490_), .A3(new_n423_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT38), .Z(new_n641_));
  INV_X1    g440(.A(new_n590_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n514_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(new_n636_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n611_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT107), .B1(new_n478_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n436_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n477_), .ZN(new_n649_));
  OAI21_X1  g448(.A(KEYINPUT104), .B1(new_n472_), .B2(new_n279_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n468_), .A2(new_n469_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n650_), .A2(new_n651_), .A3(new_n446_), .A4(new_n449_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT106), .B1(new_n652_), .B2(new_n437_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n648_), .B1(new_n649_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n655_), .A3(new_n611_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n645_), .B1(new_n647_), .B2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n490_), .B1(new_n657_), .B2(new_n423_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n641_), .A2(new_n658_), .ZN(G1324gat));
  XNOR2_X1  g458(.A(KEYINPUT109), .B(KEYINPUT40), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n647_), .A2(new_n656_), .ZN(new_n661_));
  NAND4_X1  g460(.A1(new_n661_), .A2(KEYINPUT108), .A3(new_n445_), .A4(new_n644_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G8gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(KEYINPUT108), .B1(new_n657_), .B2(new_n445_), .ZN(new_n664_));
  OAI21_X1  g463(.A(KEYINPUT39), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n661_), .A2(new_n445_), .A3(new_n644_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  NAND4_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(G8gat), .A4(new_n662_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n665_), .A2(new_n670_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n639_), .A2(new_n445_), .A3(new_n489_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n660_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n660_), .ZN(new_n675_));
  AOI211_X1 g474(.A(new_n672_), .B(new_n675_), .C1(new_n665_), .C2(new_n670_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1325gat));
  INV_X1    g476(.A(G15gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n437_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n639_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n657_), .A2(new_n679_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n681_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT41), .B1(new_n681_), .B2(G15gat), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(G1326gat));
  NAND3_X1  g483(.A1(new_n639_), .A2(new_n487_), .A3(new_n279_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n657_), .ZN(new_n686_));
  OAI21_X1  g485(.A(G22gat), .B1(new_n686_), .B2(new_n280_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n687_), .A2(KEYINPUT42), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(KEYINPUT42), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n685_), .B1(new_n688_), .B2(new_n689_), .ZN(G1327gat));
  NOR2_X1   g489(.A1(new_n478_), .A2(new_n515_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n646_), .A2(new_n636_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n590_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G29gat), .B1(new_n695_), .B2(new_n423_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n615_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n654_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n637_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n643_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n654_), .A2(KEYINPUT43), .A3(new_n697_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n700_), .A2(new_n701_), .A3(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n700_), .A2(KEYINPUT44), .A3(new_n701_), .A4(new_n702_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  AND2_X1   g506(.A1(new_n423_), .A2(G29gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n696_), .B1(new_n707_), .B2(new_n708_), .ZN(G1328gat));
  NAND3_X1  g508(.A1(new_n705_), .A2(new_n445_), .A3(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G36gat), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n392_), .B(KEYINPUT110), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n694_), .A2(G36gat), .A3(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT45), .Z(new_n714_));
  NAND2_X1  g513(.A1(new_n711_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT46), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n711_), .A2(new_n714_), .A3(KEYINPUT46), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1329gat));
  NAND4_X1  g518(.A1(new_n705_), .A2(G43gat), .A3(new_n434_), .A4(new_n706_), .ZN(new_n720_));
  INV_X1    g519(.A(G43gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n721_), .B1(new_n694_), .B2(new_n437_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g523(.A1(new_n694_), .A2(G50gat), .A3(new_n280_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n705_), .A2(new_n279_), .A3(new_n706_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(KEYINPUT111), .ZN(new_n727_));
  OAI21_X1  g526(.A(G50gat), .B1(new_n726_), .B2(KEYINPUT111), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n725_), .B1(new_n727_), .B2(new_n728_), .ZN(G1331gat));
  NOR3_X1   g528(.A1(new_n642_), .A2(new_n514_), .A3(new_n636_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n661_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(G57gat), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n447_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n478_), .A2(new_n514_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n642_), .A2(new_n638_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n737_), .A2(KEYINPUT112), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(KEYINPUT112), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n738_), .A2(new_n423_), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n733_), .B1(new_n740_), .B2(new_n732_), .ZN(G1332gat));
  OR3_X1    g540(.A1(new_n736_), .A2(G64gat), .A3(new_n712_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G64gat), .B1(new_n731_), .B2(new_n712_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n743_), .A2(KEYINPUT48), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n743_), .A2(KEYINPUT48), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n742_), .B1(new_n744_), .B2(new_n745_), .ZN(G1333gat));
  NAND3_X1  g545(.A1(new_n737_), .A2(new_n425_), .A3(new_n679_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G71gat), .B1(new_n731_), .B2(new_n437_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(KEYINPUT49), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(KEYINPUT49), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n747_), .B1(new_n749_), .B2(new_n750_), .ZN(G1334gat));
  OR3_X1    g550(.A1(new_n736_), .A2(G78gat), .A3(new_n280_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n661_), .A2(new_n279_), .A3(new_n730_), .ZN(new_n753_));
  XOR2_X1   g552(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n754_));
  AND3_X1   g553(.A1(new_n753_), .A2(G78gat), .A3(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n753_), .B2(G78gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT114), .ZN(G1335gat));
  NAND2_X1  g557(.A1(new_n698_), .A2(new_n699_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n642_), .A2(new_n514_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n759_), .A2(new_n636_), .A3(new_n702_), .A4(new_n760_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n761_), .A2(new_n447_), .A3(new_n552_), .ZN(new_n762_));
  NOR4_X1   g561(.A1(new_n478_), .A2(new_n514_), .A3(new_n642_), .A4(new_n692_), .ZN(new_n763_));
  AOI21_X1  g562(.A(G85gat), .B1(new_n763_), .B2(new_n423_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1336gat));
  OAI21_X1  g564(.A(G92gat), .B1(new_n761_), .B2(new_n712_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n763_), .A2(new_n553_), .A3(new_n445_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1337gat));
  OAI21_X1  g567(.A(G99gat), .B1(new_n761_), .B2(new_n437_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n763_), .A2(new_n548_), .A3(new_n434_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n769_), .A2(new_n770_), .B1(KEYINPUT115), .B2(new_n771_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(KEYINPUT115), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n772_), .B(new_n773_), .ZN(G1338gat));
  NAND3_X1  g573(.A1(new_n763_), .A2(new_n549_), .A3(new_n279_), .ZN(new_n775_));
  OAI21_X1  g574(.A(G106gat), .B1(new_n761_), .B2(new_n280_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n776_), .A2(KEYINPUT52), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT52), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(G106gat), .C1(new_n761_), .C2(new_n280_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n775_), .B1(new_n777_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT53), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n783_), .B(new_n775_), .C1(new_n777_), .C2(new_n780_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1339gat));
  NAND2_X1  g584(.A1(new_n564_), .A2(KEYINPUT12), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n786_), .A2(new_n566_), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT55), .B(new_n517_), .C1(new_n787_), .C2(new_n574_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n573_), .A2(new_n572_), .A3(new_n575_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n573_), .A2(new_n575_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT55), .B1(new_n791_), .B2(new_n517_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n582_), .B1(new_n790_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT56), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  OAI211_X1 g594(.A(KEYINPUT56), .B(new_n582_), .C1(new_n790_), .C2(new_n792_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(KEYINPUT121), .A3(new_n796_), .ZN(new_n797_));
  OR3_X1    g596(.A1(new_n793_), .A2(KEYINPUT121), .A3(new_n794_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n498_), .A2(new_n499_), .A3(new_n504_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT119), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n504_), .B1(new_n499_), .B2(new_n502_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(new_n510_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n801_), .A2(new_n800_), .A3(new_n510_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n799_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT120), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n807_), .B(new_n799_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n806_), .A2(new_n513_), .A3(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n585_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n797_), .A2(new_n798_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n797_), .A2(new_n798_), .A3(KEYINPUT58), .A4(new_n810_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n697_), .A3(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n515_), .A2(new_n585_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n793_), .A2(new_n817_), .A3(new_n794_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n796_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n817_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n816_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n586_), .A2(new_n809_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AND2_X1   g622(.A1(new_n611_), .A2(KEYINPUT57), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n646_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n826_));
  OAI211_X1 g625(.A(new_n815_), .B(new_n825_), .C1(KEYINPUT57), .C2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n636_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n637_), .A2(KEYINPUT116), .A3(new_n515_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT116), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n636_), .B2(new_n514_), .ZN(new_n831_));
  AOI22_X1  g630(.A1(new_n829_), .A2(new_n831_), .B1(KEYINPUT117), .B2(KEYINPUT54), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n832_), .A2(new_n615_), .A3(new_n587_), .A4(new_n589_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(KEYINPUT117), .A2(KEYINPUT54), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n833_), .B(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n828_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n393_), .A2(new_n447_), .A3(new_n435_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n828_), .B2(new_n836_), .ZN(new_n842_));
  AOI211_X1 g641(.A(KEYINPUT122), .B(new_n835_), .C1(new_n827_), .C2(new_n636_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n839_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n840_), .B1(new_n844_), .B2(KEYINPUT59), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n845_), .A2(new_n514_), .ZN(new_n846_));
  INV_X1    g645(.A(G113gat), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n514_), .A2(new_n847_), .ZN(new_n848_));
  OAI22_X1  g647(.A1(new_n846_), .A2(new_n847_), .B1(new_n844_), .B2(new_n848_), .ZN(G1340gat));
  INV_X1    g648(.A(new_n844_), .ZN(new_n850_));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n642_), .B2(KEYINPUT60), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n850_), .B(new_n852_), .C1(KEYINPUT60), .C2(new_n851_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n845_), .A2(new_n590_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n851_), .ZN(G1341gat));
  AOI21_X1  g654(.A(G127gat), .B1(new_n850_), .B2(new_n637_), .ZN(new_n856_));
  INV_X1    g655(.A(G127gat), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n636_), .A2(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT123), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n856_), .B1(new_n845_), .B2(new_n859_), .ZN(G1342gat));
  INV_X1    g659(.A(G134gat), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n850_), .A2(new_n861_), .A3(new_n646_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n845_), .A2(new_n697_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(new_n861_), .ZN(G1343gat));
  OR2_X1    g663(.A1(new_n842_), .A2(new_n843_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n712_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n437_), .A2(new_n279_), .ZN(new_n867_));
  NOR3_X1   g666(.A1(new_n866_), .A2(new_n867_), .A3(new_n447_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n865_), .A2(new_n514_), .A3(new_n868_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g669(.A1(new_n865_), .A2(new_n590_), .A3(new_n868_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g671(.A1(new_n865_), .A2(new_n637_), .A3(new_n868_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  INV_X1    g674(.A(G162gat), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n865_), .A2(new_n876_), .A3(new_n646_), .A4(new_n868_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n865_), .A2(new_n697_), .A3(new_n868_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n877_), .B1(new_n879_), .B2(new_n876_), .ZN(G1347gat));
  NAND3_X1  g679(.A1(new_n866_), .A2(new_n447_), .A3(new_n679_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n881_), .A2(new_n279_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n837_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n284_), .B1(new_n884_), .B2(new_n514_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n885_), .A2(KEYINPUT62), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(KEYINPUT62), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n884_), .A2(new_n514_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n886_), .B(new_n887_), .C1(new_n334_), .C2(new_n888_), .ZN(G1348gat));
  NOR3_X1   g688(.A1(new_n642_), .A2(new_n881_), .A3(new_n285_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n865_), .A2(new_n280_), .A3(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n883_), .A2(new_n642_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n891_), .B1(G176gat), .B2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(KEYINPUT124), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT124), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n891_), .B(new_n895_), .C1(G176gat), .C2(new_n892_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n896_), .ZN(G1349gat));
  NOR3_X1   g696(.A1(new_n883_), .A2(new_n347_), .A3(new_n636_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n881_), .A2(new_n636_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n865_), .A2(new_n280_), .A3(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n898_), .B1(new_n900_), .B2(new_n375_), .ZN(G1350gat));
  OAI21_X1  g700(.A(G190gat), .B1(new_n883_), .B2(new_n615_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n646_), .A2(new_n348_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n883_), .B2(new_n903_), .ZN(G1351gat));
  NOR3_X1   g703(.A1(new_n712_), .A2(new_n867_), .A3(new_n423_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n905_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  OAI211_X1 g707(.A(KEYINPUT125), .B(new_n905_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(G197gat), .B1(new_n910_), .B2(new_n514_), .ZN(new_n911_));
  INV_X1    g710(.A(G197gat), .ZN(new_n912_));
  AOI211_X1 g711(.A(new_n912_), .B(new_n515_), .C1(new_n908_), .C2(new_n909_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n911_), .A2(new_n913_), .ZN(G1352gat));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n915_), .A2(G204gat), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n642_), .B1(new_n915_), .B2(G204gat), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n910_), .B2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n918_), .ZN(new_n920_));
  AOI211_X1 g719(.A(new_n920_), .B(new_n916_), .C1(new_n908_), .C2(new_n909_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n919_), .A2(new_n921_), .ZN(G1353gat));
  NOR2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(KEYINPUT127), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n636_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n924_), .B1(new_n910_), .B2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n925_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n924_), .ZN(new_n928_));
  AOI211_X1 g727(.A(new_n927_), .B(new_n928_), .C1(new_n908_), .C2(new_n909_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n926_), .A2(new_n929_), .ZN(G1354gat));
  INV_X1    g729(.A(G218gat), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n910_), .A2(new_n931_), .A3(new_n646_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n615_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n931_), .B2(new_n933_), .ZN(G1355gat));
endmodule


