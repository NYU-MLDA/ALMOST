//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n945_, new_n946_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_, new_n973_, new_n975_, new_n976_, new_n977_,
    new_n978_, new_n979_, new_n981_, new_n982_, new_n984_, new_n985_,
    new_n986_, new_n987_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n1000_,
    new_n1001_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT19), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT20), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT24), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n211_), .B1(G169gat), .B2(G176gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT82), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n212_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(KEYINPUT25), .B(G183gat), .Z(new_n218_));
  XOR2_X1   g017(.A(KEYINPUT26), .B(G190gat), .Z(new_n219_));
  OAI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G183gat), .ZN(new_n221_));
  INV_X1    g020(.A(G190gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT23), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(G183gat), .A3(G190gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(KEYINPUT83), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT83), .ZN(new_n227_));
  OAI211_X1 g026(.A(new_n227_), .B(KEYINPUT23), .C1(new_n221_), .C2(new_n222_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n213_), .A2(new_n211_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n226_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT94), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT94), .ZN(new_n232_));
  NAND4_X1  g031(.A1(new_n226_), .A2(new_n232_), .A3(new_n228_), .A4(new_n229_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n220_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  AOI22_X1  g033(.A1(new_n223_), .A2(new_n225_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n235_), .A2(KEYINPUT95), .ZN(new_n236_));
  NOR2_X1   g035(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(G169gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n238_), .B1(new_n235_), .B2(KEYINPUT95), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n236_), .A2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n234_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G204gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(G197gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT91), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT91), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n245_), .A2(new_n242_), .A3(G197gat), .ZN(new_n246_));
  INV_X1    g045(.A(G197gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G204gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n244_), .A2(new_n246_), .A3(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT21), .ZN(new_n250_));
  INV_X1    g049(.A(G218gat), .ZN(new_n251_));
  OR2_X1    g050(.A1(new_n251_), .A2(G211gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(G211gat), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n250_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n249_), .A2(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n250_), .B1(new_n243_), .B2(new_n248_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT90), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n244_), .A2(new_n246_), .A3(new_n250_), .A4(new_n248_), .ZN(new_n259_));
  AND2_X1   g058(.A1(new_n252_), .A2(new_n253_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n255_), .B1(new_n258_), .B2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n210_), .B1(new_n241_), .B2(new_n262_), .ZN(new_n263_));
  OR2_X1    g062(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n264_));
  OR2_X1    g063(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(KEYINPUT81), .A2(G190gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(KEYINPUT80), .A2(G183gat), .ZN(new_n267_));
  NAND4_X1  g066(.A1(new_n264_), .A2(new_n265_), .A3(new_n266_), .A4(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n226_), .A2(new_n268_), .A3(new_n228_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT84), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n226_), .A2(new_n268_), .A3(KEYINPUT84), .A4(new_n228_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(new_n238_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n223_), .A2(new_n225_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n217_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n215_), .A2(new_n216_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(new_n211_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n264_), .A2(new_n266_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n278_), .B1(new_n279_), .B2(KEYINPUT26), .ZN(new_n280_));
  NOR2_X1   g079(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n265_), .A2(new_n267_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n281_), .B1(new_n282_), .B2(KEYINPUT25), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n275_), .B(new_n277_), .C1(new_n280_), .C2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n273_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n249_), .A2(new_n254_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n256_), .B(KEYINPUT90), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n259_), .A2(new_n260_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n286_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n209_), .B1(new_n263_), .B2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n234_), .B2(new_n240_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n262_), .A2(new_n273_), .A3(new_n284_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n292_), .A2(KEYINPUT20), .A3(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n208_), .B(KEYINPUT93), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n206_), .B1(new_n291_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT27), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n295_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT96), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n263_), .A2(new_n209_), .A3(new_n290_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT96), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n294_), .A2(new_n302_), .A3(new_n295_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n300_), .A2(new_n205_), .A3(new_n301_), .A4(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT99), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n303_), .A2(new_n301_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT99), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(new_n205_), .A4(new_n300_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n298_), .B1(new_n305_), .B2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n303_), .A2(new_n301_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n302_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n206_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT27), .B1(new_n312_), .B2(new_n304_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n309_), .A2(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(G22gat), .B(G50gat), .Z(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n317_));
  NOR2_X1   g116(.A1(G141gat), .A2(G148gat), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT3), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G141gat), .A2(G148gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT2), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n320_), .A2(new_n323_), .A3(new_n324_), .A4(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G155gat), .B(G162gat), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  AND2_X1   g128(.A1(G141gat), .A2(G148gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n330_), .A2(new_n318_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n332_));
  OAI211_X1 g131(.A(new_n331_), .B(new_n332_), .C1(new_n327_), .C2(KEYINPUT1), .ZN(new_n333_));
  AND3_X1   g132(.A1(new_n329_), .A2(KEYINPUT88), .A3(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(KEYINPUT88), .B1(new_n329_), .B2(new_n333_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n317_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT28), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n329_), .A2(new_n333_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT88), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n329_), .A2(KEYINPUT88), .A3(new_n333_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT28), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(new_n343_), .A3(new_n317_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT89), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n337_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n345_), .B1(new_n337_), .B2(new_n344_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n316_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n337_), .A2(new_n344_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT89), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(new_n315_), .A3(new_n346_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n349_), .A2(new_n352_), .A3(KEYINPUT92), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n340_), .A2(KEYINPUT29), .A3(new_n341_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G228gat), .A2(G233gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n289_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n317_), .B1(new_n329_), .B2(new_n333_), .ZN(new_n357_));
  OAI211_X1 g156(.A(G228gat), .B(G233gat), .C1(new_n262_), .C2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G78gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n356_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n359_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n362_));
  OAI21_X1  g161(.A(G106gat), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n356_), .A2(new_n358_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(G78gat), .ZN(new_n365_));
  INV_X1    g164(.A(G106gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(new_n360_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n363_), .A2(new_n367_), .ZN(new_n368_));
  OR2_X1    g167(.A1(new_n353_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT92), .ZN(new_n370_));
  NOR3_X1   g169(.A1(new_n347_), .A2(new_n348_), .A3(new_n316_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n315_), .B1(new_n351_), .B2(new_n346_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n373_), .A2(new_n353_), .A3(new_n368_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n369_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n285_), .A2(KEYINPUT30), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n273_), .A2(new_n284_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G227gat), .A2(G233gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT85), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G15gat), .B(G43gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n380_), .B(KEYINPUT85), .ZN(new_n385_));
  INV_X1    g184(.A(new_n383_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n384_), .A2(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G71gat), .B(G99gat), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n384_), .A2(new_n387_), .A3(new_n389_), .ZN(new_n392_));
  AOI21_X1  g191(.A(KEYINPUT86), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n379_), .A2(new_n393_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n391_), .A2(KEYINPUT86), .A3(new_n392_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n395_), .A2(new_n393_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(new_n378_), .A3(new_n376_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT87), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n394_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT31), .ZN(new_n400_));
  XOR2_X1   g199(.A(G127gat), .B(G134gat), .Z(new_n401_));
  INV_X1    g200(.A(G120gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(G113gat), .ZN(new_n403_));
  INV_X1    g202(.A(G113gat), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(G120gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G127gat), .B(G134gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n408_), .A2(new_n403_), .A3(new_n405_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT31), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n394_), .A2(new_n397_), .A3(new_n398_), .A4(new_n412_), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n400_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(G85gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT0), .B(G57gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G225gat), .A2(G233gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n340_), .A2(new_n341_), .A3(new_n411_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(new_n421_), .B2(KEYINPUT4), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n410_), .A2(new_n333_), .A3(new_n329_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT97), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n410_), .A2(KEYINPUT97), .A3(new_n333_), .A4(new_n329_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n421_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT4), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT98), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n334_), .A2(new_n335_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n431_), .A2(new_n411_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT98), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(KEYINPUT4), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n422_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n428_), .A2(new_n420_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n418_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n422_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n433_), .B1(new_n432_), .B2(KEYINPUT4), .ZN(new_n439_));
  AND4_X1   g238(.A1(new_n433_), .A2(new_n427_), .A3(KEYINPUT4), .A4(new_n421_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n438_), .B1(new_n439_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n418_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n436_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n437_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n411_), .B1(new_n400_), .B2(new_n413_), .ZN(new_n446_));
  NOR3_X1   g245(.A1(new_n414_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n314_), .A2(new_n375_), .A3(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n418_), .B1(new_n428_), .B2(new_n419_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n430_), .A2(new_n434_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n421_), .A2(KEYINPUT4), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n451_), .A2(new_n420_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n449_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n444_), .A2(KEYINPUT33), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT33), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n441_), .A2(new_n455_), .A3(new_n442_), .A4(new_n443_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n453_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n312_), .A2(new_n304_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n306_), .A2(new_n300_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n460_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n291_), .A2(new_n296_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n437_), .A2(new_n444_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n457_), .A2(new_n459_), .B1(new_n461_), .B2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n369_), .A2(new_n374_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT27), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n458_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n445_), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n468_), .A2(new_n369_), .A3(new_n469_), .A4(new_n374_), .ZN(new_n470_));
  OAI22_X1  g269(.A1(new_n465_), .A2(new_n466_), .B1(new_n470_), .B2(new_n309_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n414_), .A2(new_n446_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n448_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(G190gat), .B(G218gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT72), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G134gat), .B(G162gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT36), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G232gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT34), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT35), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G85gat), .A2(G92gat), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n487_), .A2(KEYINPUT9), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G99gat), .A2(G106gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT6), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT6), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(G99gat), .A3(G106gat), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n488_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n493_));
  OR2_X1    g292(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n494_), .A2(new_n366_), .A3(new_n495_), .ZN(new_n496_));
  OR2_X1    g295(.A1(G85gat), .A2(G92gat), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(KEYINPUT9), .A3(new_n487_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n493_), .A2(new_n496_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT67), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n493_), .A2(KEYINPUT67), .A3(new_n496_), .A4(new_n498_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT65), .ZN(new_n503_));
  INV_X1    g302(.A(G99gat), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n503_), .A2(new_n504_), .A3(new_n366_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT7), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n490_), .A2(new_n492_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT7), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n503_), .A2(new_n508_), .A3(new_n504_), .A4(new_n366_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n506_), .A2(new_n507_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT8), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n497_), .A2(new_n487_), .ZN(new_n512_));
  AND3_X1   g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n511_), .B1(new_n510_), .B2(new_n512_), .ZN(new_n514_));
  OAI211_X1 g313(.A(new_n501_), .B(new_n502_), .C1(new_n513_), .C2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G29gat), .B(G36gat), .Z(new_n516_));
  INV_X1    g315(.A(G50gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(G43gat), .ZN(new_n518_));
  INV_X1    g317(.A(G43gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(G50gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n518_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G29gat), .B(G36gat), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n523_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n522_), .A2(KEYINPUT15), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT15), .B1(new_n522_), .B2(new_n524_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n515_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(KEYINPUT71), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT71), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n515_), .A2(new_n530_), .A3(new_n527_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n499_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n510_), .A2(new_n512_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT8), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n533_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n522_), .A2(new_n524_), .ZN(new_n538_));
  AOI22_X1  g337(.A1(new_n537_), .A2(new_n538_), .B1(new_n484_), .B2(new_n483_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n486_), .B1(new_n532_), .B2(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n515_), .A2(new_n530_), .A3(new_n527_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n530_), .B1(new_n515_), .B2(new_n527_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n486_), .B(new_n539_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n480_), .B1(new_n540_), .B2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT74), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n539_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n485_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n478_), .A2(KEYINPUT36), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n543_), .A3(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n479_), .B1(new_n548_), .B2(new_n543_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT74), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n546_), .A2(new_n550_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n474_), .A2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n499_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n557_));
  INV_X1    g356(.A(G64gat), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(G57gat), .ZN(new_n559_));
  INV_X1    g358(.A(G57gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(G64gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT66), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n559_), .A2(new_n561_), .A3(KEYINPUT66), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G71gat), .B(G78gat), .Z(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(KEYINPUT11), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n565_), .ZN(new_n570_));
  AOI21_X1  g369(.A(KEYINPUT66), .B1(new_n559_), .B2(new_n561_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT11), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT11), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n564_), .A2(new_n573_), .A3(new_n565_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n572_), .A2(new_n574_), .A3(new_n567_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n557_), .A2(new_n569_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n569_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n537_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G230gat), .A2(G233gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT64), .Z(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n583_), .B1(new_n537_), .B2(new_n577_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n581_), .B1(new_n537_), .B2(new_n577_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n575_), .A2(KEYINPUT12), .A3(new_n569_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n515_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n584_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G120gat), .B(G148gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G176gat), .B(G204gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n582_), .A2(new_n588_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n593_), .B1(new_n582_), .B2(new_n588_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT13), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT13), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n598_), .A2(new_n599_), .A3(new_n594_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n597_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G113gat), .B(G141gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G169gat), .B(G197gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n603_), .B(new_n604_), .Z(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT76), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT14), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT75), .B(G8gat), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(G1gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(G15gat), .B(G22gat), .Z(new_n611_));
  OAI21_X1  g410(.A(new_n607_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(KEYINPUT75), .A2(G8gat), .ZN(new_n613_));
  NOR2_X1   g412(.A1(KEYINPUT75), .A2(G8gat), .ZN(new_n614_));
  OAI21_X1  g413(.A(G1gat), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(KEYINPUT14), .ZN(new_n616_));
  INV_X1    g415(.A(new_n611_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(new_n617_), .A3(KEYINPUT76), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G1gat), .B(G8gat), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n612_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n619_), .B1(new_n612_), .B2(new_n618_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n538_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G229gat), .A2(G233gat), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n619_), .ZN(new_n625_));
  NOR3_X1   g424(.A1(new_n610_), .A2(new_n607_), .A3(new_n611_), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT76), .B1(new_n616_), .B2(new_n617_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n625_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n612_), .A2(new_n618_), .A3(new_n619_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n628_), .A2(new_n527_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT78), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT78), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n628_), .A2(new_n527_), .A3(new_n632_), .A4(new_n629_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n624_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n538_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n628_), .A2(new_n635_), .A3(new_n629_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n623_), .B1(new_n622_), .B2(new_n636_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n606_), .B1(new_n634_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n637_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n631_), .A2(new_n633_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n639_), .B(new_n605_), .C1(new_n640_), .C2(new_n624_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(KEYINPUT79), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT79), .ZN(new_n643_));
  OAI211_X1 g442(.A(new_n643_), .B(new_n606_), .C1(new_n634_), .C2(new_n637_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  AND2_X1   g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n577_), .B(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n628_), .A2(new_n629_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(G127gat), .B(G155gat), .Z(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT16), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G183gat), .B(G211gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT17), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n649_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n654_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n649_), .A2(new_n655_), .A3(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n656_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n602_), .A2(new_n645_), .A3(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n556_), .A2(new_n445_), .A3(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G1gat), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT38), .ZN(new_n664_));
  INV_X1    g463(.A(new_n474_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n550_), .B1(new_n551_), .B2(KEYINPUT73), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT73), .ZN(new_n667_));
  AOI211_X1 g466(.A(new_n667_), .B(new_n479_), .C1(new_n548_), .C2(new_n543_), .ZN(new_n668_));
  OAI21_X1  g467(.A(KEYINPUT37), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT37), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n546_), .A2(new_n553_), .A3(new_n670_), .A4(new_n550_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n659_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT77), .ZN(new_n674_));
  INV_X1    g473(.A(new_n645_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n601_), .B(KEYINPUT70), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n665_), .A2(new_n674_), .A3(new_n675_), .A4(new_n676_), .ZN(new_n677_));
  OR3_X1    g476(.A1(new_n677_), .A2(G1gat), .A3(new_n469_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n678_), .A2(KEYINPUT100), .A3(new_n664_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT100), .B1(new_n678_), .B2(new_n664_), .ZN(new_n680_));
  OAI221_X1 g479(.A(new_n663_), .B1(new_n664_), .B2(new_n678_), .C1(new_n679_), .C2(new_n680_), .ZN(G1324gat));
  INV_X1    g480(.A(new_n314_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n556_), .A2(new_n682_), .A3(new_n661_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT39), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n683_), .A2(new_n684_), .A3(G8gat), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(new_n683_), .B2(G8gat), .ZN(new_n687_));
  OR2_X1    g486(.A1(new_n314_), .A2(new_n609_), .ZN(new_n688_));
  OAI22_X1  g487(.A1(new_n686_), .A2(new_n687_), .B1(new_n677_), .B2(new_n688_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g489(.A1(new_n556_), .A2(new_n472_), .A3(new_n661_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(KEYINPUT41), .B1(new_n691_), .B2(G15gat), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n473_), .A2(G15gat), .ZN(new_n695_));
  OAI22_X1  g494(.A1(new_n693_), .A2(new_n694_), .B1(new_n677_), .B2(new_n695_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT101), .ZN(G1326gat));
  NAND3_X1  g496(.A1(new_n556_), .A2(new_n466_), .A3(new_n661_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G22gat), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n700_));
  XNOR2_X1  g499(.A(new_n699_), .B(new_n700_), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n375_), .A2(G22gat), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n701_), .B1(new_n677_), .B2(new_n702_), .ZN(G1327gat));
  NAND2_X1  g502(.A1(new_n555_), .A2(new_n660_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n704_), .A2(new_n602_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n464_), .A2(new_n461_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n453_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n436_), .B1(new_n450_), .B2(new_n438_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n455_), .B1(new_n708_), .B2(new_n442_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n456_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n707_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n706_), .B1(new_n711_), .B2(new_n458_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(new_n375_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n309_), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n466_), .A2(new_n469_), .A3(new_n714_), .A4(new_n468_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n472_), .B1(new_n713_), .B2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(new_n675_), .B(new_n705_), .C1(new_n716_), .C2(new_n448_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT103), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT103), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n665_), .A2(new_n719_), .A3(new_n675_), .A4(new_n705_), .ZN(new_n720_));
  INV_X1    g519(.A(G29gat), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n445_), .A2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT104), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n718_), .A2(new_n720_), .A3(new_n723_), .ZN(new_n724_));
  OAI21_X1  g523(.A(KEYINPUT43), .B1(new_n474_), .B2(new_n672_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT43), .ZN(new_n726_));
  INV_X1    g525(.A(new_n672_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n726_), .B(new_n727_), .C1(new_n716_), .C2(new_n448_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n602_), .A2(new_n645_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n660_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT44), .B1(new_n729_), .B2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT44), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n734_), .B(new_n731_), .C1(new_n725_), .C2(new_n728_), .ZN(new_n735_));
  NOR3_X1   g534(.A1(new_n733_), .A2(new_n735_), .A3(new_n469_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n724_), .B1(new_n736_), .B2(new_n721_), .ZN(G1328gat));
  INV_X1    g536(.A(KEYINPUT46), .ZN(new_n738_));
  INV_X1    g537(.A(G36gat), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n733_), .A2(new_n735_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(new_n682_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n718_), .A2(new_n720_), .A3(new_n739_), .A4(new_n682_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n738_), .B1(new_n741_), .B2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n742_), .B(KEYINPUT45), .ZN(new_n746_));
  NOR3_X1   g545(.A1(new_n733_), .A2(new_n735_), .A3(new_n314_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n746_), .B(KEYINPUT46), .C1(new_n739_), .C2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n745_), .A2(new_n748_), .ZN(G1329gat));
  NOR2_X1   g548(.A1(new_n473_), .A2(new_n519_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n740_), .A2(new_n750_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n718_), .A2(new_n720_), .A3(new_n472_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n752_), .A2(new_n519_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT47), .B1(new_n751_), .B2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n740_), .B2(new_n750_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT47), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n754_), .A2(new_n757_), .ZN(G1330gat));
  NOR2_X1   g557(.A1(new_n375_), .A2(new_n517_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n718_), .A2(new_n720_), .A3(new_n466_), .ZN(new_n760_));
  AOI22_X1  g559(.A1(new_n740_), .A2(new_n759_), .B1(new_n517_), .B2(new_n760_), .ZN(G1331gat));
  AND2_X1   g560(.A1(new_n674_), .A2(new_n602_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT105), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n474_), .A2(new_n675_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(KEYINPUT105), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n763_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(new_n560_), .A3(new_n445_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n676_), .A2(new_n675_), .A3(new_n660_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n556_), .A2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G57gat), .B1(new_n769_), .B2(new_n469_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(new_n770_), .ZN(G1332gat));
  NOR2_X1   g570(.A1(new_n314_), .A2(G64gat), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n763_), .A2(new_n764_), .A3(new_n765_), .A4(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n556_), .A2(new_n682_), .A3(new_n768_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(G64gat), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n775_), .B1(new_n774_), .B2(G64gat), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n773_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT106), .ZN(G1333gat));
  INV_X1    g579(.A(G71gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n766_), .A2(new_n781_), .A3(new_n472_), .ZN(new_n782_));
  OAI21_X1  g581(.A(G71gat), .B1(new_n769_), .B2(new_n473_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT49), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1334gat));
  NAND3_X1  g584(.A1(new_n766_), .A2(new_n359_), .A3(new_n466_), .ZN(new_n786_));
  OAI21_X1  g585(.A(G78gat), .B1(new_n769_), .B2(new_n375_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n787_), .B(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(G1335gat));
  INV_X1    g589(.A(new_n729_), .ZN(new_n791_));
  NOR3_X1   g590(.A1(new_n675_), .A2(new_n659_), .A3(new_n601_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n791_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(G85gat), .A3(new_n445_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n676_), .A2(new_n704_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n764_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n445_), .ZN(new_n799_));
  INV_X1    g598(.A(G85gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT108), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT108), .B(new_n800_), .C1(new_n797_), .C2(new_n469_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n795_), .B1(new_n801_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT109), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n795_), .B(new_n806_), .C1(new_n801_), .C2(new_n803_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1336gat));
  AOI21_X1  g607(.A(G92gat), .B1(new_n798_), .B2(new_n682_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n682_), .A2(G92gat), .ZN(new_n810_));
  XOR2_X1   g609(.A(new_n810_), .B(KEYINPUT110), .Z(new_n811_));
  AOI21_X1  g610(.A(new_n809_), .B1(new_n794_), .B2(new_n811_), .ZN(G1337gat));
  AOI21_X1  g611(.A(new_n504_), .B1(new_n794_), .B2(new_n472_), .ZN(new_n813_));
  AND4_X1   g612(.A1(new_n472_), .A2(new_n798_), .A3(new_n494_), .A4(new_n495_), .ZN(new_n814_));
  OR3_X1    g613(.A1(new_n813_), .A2(KEYINPUT51), .A3(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT51), .B1(new_n813_), .B2(new_n814_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(G1338gat));
  NAND3_X1  g616(.A1(new_n798_), .A2(new_n366_), .A3(new_n466_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n729_), .A2(new_n466_), .A3(new_n792_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n819_), .A2(new_n820_), .A3(G106gat), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n820_), .B1(new_n819_), .B2(G106gat), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n818_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT53), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n825_), .B(new_n818_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1339gat));
  NOR2_X1   g626(.A1(new_n473_), .A2(new_n469_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n828_), .A2(new_n829_), .A3(new_n375_), .A4(new_n314_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n314_), .A2(new_n445_), .A3(new_n375_), .A4(new_n472_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT114), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT112), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n622_), .A2(G229gat), .A3(G233gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n620_), .A2(new_n621_), .A3(new_n538_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n635_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n623_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n840_), .A2(new_n606_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n835_), .B1(new_n837_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n622_), .A2(new_n636_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n605_), .B1(new_n843_), .B2(new_n623_), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n844_), .B(KEYINPUT112), .C1(new_n640_), .C2(new_n836_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n842_), .A2(new_n641_), .A3(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n595_), .A2(new_n596_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n642_), .A2(new_n644_), .A3(new_n594_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n588_), .A2(KEYINPUT55), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n584_), .A2(new_n585_), .A3(new_n587_), .A4(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n850_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n584_), .A2(new_n587_), .A3(new_n578_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n581_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n593_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n856_));
  XOR2_X1   g655(.A(KEYINPUT111), .B(KEYINPUT56), .Z(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n850_), .A2(new_n852_), .B1(new_n581_), .B2(new_n854_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n593_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  OAI22_X1  g661(.A1(new_n856_), .A2(new_n858_), .B1(new_n859_), .B2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n848_), .B1(new_n849_), .B2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n834_), .B1(new_n864_), .B2(new_n555_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n598_), .A2(new_n594_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n866_), .A2(new_n641_), .A3(new_n842_), .A4(new_n845_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n862_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n576_), .A2(new_n583_), .B1(new_n515_), .B2(new_n586_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n851_), .B1(new_n869_), .B2(new_n585_), .ZN(new_n870_));
  AND4_X1   g669(.A1(new_n851_), .A2(new_n584_), .A3(new_n585_), .A4(new_n587_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n855_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n593_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n868_), .B1(new_n874_), .B2(new_n857_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n642_), .A2(new_n644_), .A3(new_n594_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n867_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(KEYINPUT57), .A3(new_n554_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n865_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT113), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n859_), .B2(new_n862_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n860_), .B1(new_n859_), .B2(new_n593_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n872_), .A2(KEYINPUT113), .A3(new_n861_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n881_), .A2(new_n882_), .A3(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n846_), .A2(new_n595_), .ZN(new_n885_));
  AND3_X1   g684(.A1(new_n884_), .A2(KEYINPUT58), .A3(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(KEYINPUT58), .B1(new_n884_), .B2(new_n885_), .ZN(new_n887_));
  NOR3_X1   g686(.A1(new_n886_), .A2(new_n887_), .A3(new_n672_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n660_), .B1(new_n879_), .B2(new_n888_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n659_), .A2(new_n601_), .A3(new_n645_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n672_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT54), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n833_), .B1(new_n889_), .B2(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(G113gat), .B1(new_n893_), .B2(new_n675_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(KEYINPUT115), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n896_));
  INV_X1    g695(.A(new_n833_), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n877_), .A2(KEYINPUT57), .A3(new_n554_), .ZN(new_n898_));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n877_), .B2(new_n554_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  OR3_X1    g699(.A1(new_n886_), .A2(new_n887_), .A3(new_n672_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n659_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n891_), .B(new_n903_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n896_), .B(new_n897_), .C1(new_n902_), .C2(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n905_), .A2(KEYINPUT116), .A3(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT118), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n889_), .A2(new_n892_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT116), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n909_), .A2(new_n910_), .A3(new_n897_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(KEYINPUT59), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n910_), .B1(new_n893_), .B2(new_n896_), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n907_), .B(new_n908_), .C1(new_n912_), .C2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  AOI211_X1 g714(.A(KEYINPUT117), .B(new_n833_), .C1(new_n889_), .C2(new_n892_), .ZN(new_n916_));
  OAI211_X1 g715(.A(KEYINPUT59), .B(new_n911_), .C1(new_n916_), .C2(new_n910_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n908_), .B1(new_n917_), .B2(new_n907_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n915_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n645_), .A2(new_n404_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n895_), .B1(new_n919_), .B2(new_n920_), .ZN(G1340gat));
  OAI21_X1  g720(.A(new_n402_), .B1(new_n601_), .B2(KEYINPUT60), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n893_), .B(new_n922_), .C1(KEYINPUT60), .C2(new_n402_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n676_), .B1(new_n917_), .B2(new_n907_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n923_), .B1(new_n924_), .B2(new_n402_), .ZN(G1341gat));
  AOI21_X1  g724(.A(G127gat), .B1(new_n893_), .B2(new_n659_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n659_), .A2(G127gat), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n927_), .B(KEYINPUT119), .Z(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n919_), .B2(new_n928_), .ZN(G1342gat));
  AOI21_X1  g728(.A(G134gat), .B1(new_n893_), .B2(new_n555_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n727_), .A2(G134gat), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(new_n919_), .B2(new_n931_), .ZN(G1343gat));
  AOI21_X1  g731(.A(new_n472_), .B1(new_n889_), .B2(new_n892_), .ZN(new_n933_));
  AND4_X1   g732(.A1(new_n445_), .A2(new_n933_), .A3(new_n466_), .A4(new_n314_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n675_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(KEYINPUT120), .B(G141gat), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n935_), .B(new_n936_), .ZN(G1344gat));
  INV_X1    g736(.A(new_n676_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n934_), .A2(new_n938_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT121), .B(G148gat), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n939_), .B(new_n940_), .ZN(G1345gat));
  NAND2_X1  g740(.A1(new_n934_), .A2(new_n659_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(KEYINPUT61), .B(G155gat), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1346gat));
  INV_X1    g743(.A(G162gat), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n934_), .A2(new_n945_), .A3(new_n555_), .ZN(new_n946_));
  AND2_X1   g745(.A1(new_n934_), .A2(new_n727_), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n947_), .B2(new_n945_), .ZN(G1347gat));
  AND3_X1   g747(.A1(new_n682_), .A2(new_n375_), .A3(new_n447_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(new_n675_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n950_), .B1(new_n889_), .B2(new_n892_), .ZN(new_n951_));
  INV_X1    g750(.A(G169gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(KEYINPUT62), .B1(new_n951_), .B2(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n953_), .A2(KEYINPUT123), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT123), .ZN(new_n955_));
  OAI211_X1 g754(.A(new_n955_), .B(KEYINPUT62), .C1(new_n951_), .C2(new_n952_), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT122), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n952_), .A2(KEYINPUT62), .ZN(new_n958_));
  INV_X1    g757(.A(new_n958_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n957_), .B1(new_n951_), .B2(new_n959_), .ZN(new_n960_));
  INV_X1    g759(.A(new_n951_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n961_), .A2(KEYINPUT122), .A3(new_n958_), .ZN(new_n962_));
  NAND4_X1  g761(.A1(new_n954_), .A2(new_n956_), .A3(new_n960_), .A4(new_n962_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(KEYINPUT22), .B(G169gat), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n951_), .A2(new_n964_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n963_), .A2(new_n965_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n966_), .A2(KEYINPUT124), .ZN(new_n967_));
  INV_X1    g766(.A(KEYINPUT124), .ZN(new_n968_));
  NAND3_X1  g767(.A1(new_n963_), .A2(new_n968_), .A3(new_n965_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n967_), .A2(new_n969_), .ZN(G1348gat));
  NAND2_X1  g769(.A1(new_n909_), .A2(new_n949_), .ZN(new_n971_));
  OAI21_X1  g770(.A(G176gat), .B1(new_n971_), .B2(new_n676_), .ZN(new_n972_));
  OR2_X1    g771(.A1(new_n601_), .A2(G176gat), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n972_), .B1(new_n971_), .B2(new_n973_), .ZN(G1349gat));
  NOR2_X1   g773(.A1(new_n971_), .A2(new_n660_), .ZN(new_n975_));
  INV_X1    g774(.A(new_n282_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n218_), .B1(new_n976_), .B2(KEYINPUT125), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n975_), .A2(new_n977_), .ZN(new_n978_));
  NOR2_X1   g777(.A1(new_n282_), .A2(KEYINPUT125), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n978_), .B1(new_n975_), .B2(new_n979_), .ZN(G1350gat));
  OAI21_X1  g779(.A(G190gat), .B1(new_n971_), .B2(new_n672_), .ZN(new_n981_));
  OR2_X1    g780(.A1(new_n554_), .A2(new_n219_), .ZN(new_n982_));
  OAI21_X1  g781(.A(new_n981_), .B1(new_n971_), .B2(new_n982_), .ZN(G1351gat));
  NOR3_X1   g782(.A1(new_n314_), .A2(new_n445_), .A3(new_n375_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n933_), .A2(new_n984_), .ZN(new_n985_));
  NOR2_X1   g784(.A1(new_n985_), .A2(new_n645_), .ZN(new_n986_));
  XNOR2_X1  g785(.A(KEYINPUT126), .B(G197gat), .ZN(new_n987_));
  XNOR2_X1  g786(.A(new_n986_), .B(new_n987_), .ZN(G1352gat));
  NOR2_X1   g787(.A1(new_n985_), .A2(new_n676_), .ZN(new_n989_));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n989_), .B1(new_n990_), .B2(new_n242_), .ZN(new_n991_));
  XOR2_X1   g790(.A(KEYINPUT127), .B(G204gat), .Z(new_n992_));
  OAI21_X1  g791(.A(new_n991_), .B1(new_n989_), .B2(new_n992_), .ZN(G1353gat));
  INV_X1    g792(.A(new_n985_), .ZN(new_n994_));
  NAND2_X1  g793(.A1(new_n994_), .A2(new_n659_), .ZN(new_n995_));
  NOR2_X1   g794(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n996_));
  AND2_X1   g795(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n997_));
  NOR3_X1   g796(.A1(new_n995_), .A2(new_n996_), .A3(new_n997_), .ZN(new_n998_));
  AOI21_X1  g797(.A(new_n998_), .B1(new_n995_), .B2(new_n996_), .ZN(G1354gat));
  OAI21_X1  g798(.A(G218gat), .B1(new_n985_), .B2(new_n672_), .ZN(new_n1000_));
  NAND2_X1  g799(.A1(new_n555_), .A2(new_n251_), .ZN(new_n1001_));
  OAI21_X1  g800(.A(new_n1000_), .B1(new_n985_), .B2(new_n1001_), .ZN(G1355gat));
endmodule


