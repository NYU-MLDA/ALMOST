//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n737_, new_n738_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n781_, new_n782_, new_n784_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n913_, new_n914_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n927_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n947_,
    new_n948_, new_n949_, new_n951_, new_n952_, new_n953_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n961_,
    new_n963_, new_n964_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(G155gat), .ZN(new_n203_));
  INV_X1    g002(.A(G162gat), .ZN(new_n204_));
  OR3_X1    g003(.A1(new_n203_), .A2(new_n204_), .A3(KEYINPUT1), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT1), .B1(new_n203_), .B2(new_n204_), .ZN(new_n206_));
  OAI211_X1 g005(.A(new_n205_), .B(new_n206_), .C1(G155gat), .C2(G162gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G141gat), .A2(G148gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n207_), .A2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT3), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n208_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n214_), .A2(new_n216_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(G155gat), .B(G162gat), .Z(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(KEYINPUT86), .A3(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT86), .B1(new_n219_), .B2(new_n220_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n212_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G127gat), .ZN(new_n225_));
  INV_X1    g024(.A(G134gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT85), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G127gat), .A2(G134gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n228_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n232_));
  OAI21_X1  g031(.A(G113gat), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(new_n229_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT85), .ZN(new_n235_));
  INV_X1    g034(.A(G113gat), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n230_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n233_), .A2(G120gat), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  AOI21_X1  g038(.A(G120gat), .B1(new_n233_), .B2(new_n237_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n224_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n219_), .A2(new_n220_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT86), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  AOI22_X1  g043(.A1(new_n244_), .A2(new_n221_), .B1(new_n207_), .B2(new_n211_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n233_), .A2(new_n237_), .ZN(new_n246_));
  INV_X1    g045(.A(G120gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n245_), .A2(new_n248_), .A3(new_n238_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n241_), .A2(new_n249_), .A3(KEYINPUT4), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G225gat), .A2(G233gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n238_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(new_n224_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n250_), .A2(new_n252_), .A3(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(KEYINPUT93), .B(KEYINPUT0), .Z(new_n257_));
  XNOR2_X1  g056(.A(G1gat), .B(G29gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G57gat), .B(G85gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n241_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n256_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n262_), .B1(new_n256_), .B2(new_n263_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT94), .ZN(new_n267_));
  INV_X1    g066(.A(G197gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n268_), .A2(G204gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(KEYINPUT87), .B(G197gat), .Z(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n270_), .B2(G204gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT21), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G211gat), .B(G218gat), .ZN(new_n273_));
  OR3_X1    g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G197gat), .A2(G204gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT87), .B(G197gat), .ZN(new_n277_));
  OAI211_X1 g076(.A(KEYINPUT21), .B(new_n276_), .C1(new_n277_), .C2(G204gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n269_), .ZN(new_n279_));
  INV_X1    g078(.A(G204gat), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n272_), .B(new_n279_), .C1(new_n277_), .C2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n278_), .A2(new_n281_), .A3(new_n273_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT88), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  OR2_X1    g083(.A1(new_n282_), .A2(new_n283_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n275_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G169gat), .ZN(new_n287_));
  INV_X1    g086(.A(G176gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(KEYINPUT24), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT82), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT25), .B(G183gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(G190gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n289_), .A2(KEYINPUT82), .A3(KEYINPUT24), .A4(new_n290_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT83), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT23), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n289_), .A2(KEYINPUT24), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n293_), .A2(new_n296_), .A3(KEYINPUT83), .A4(new_n297_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n300_), .A2(new_n302_), .A3(new_n303_), .A4(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n302_), .B1(G183gat), .B2(G190gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G169gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n305_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n286_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n282_), .B(new_n283_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n274_), .ZN(new_n313_));
  XOR2_X1   g112(.A(KEYINPUT90), .B(KEYINPUT24), .Z(new_n314_));
  NAND3_X1  g113(.A1(new_n314_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n296_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT91), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  OR2_X1    g117(.A1(new_n314_), .A2(new_n289_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(KEYINPUT91), .A3(new_n296_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n318_), .A2(new_n302_), .A3(new_n319_), .A4(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n309_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n313_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT19), .ZN(new_n325_));
  AND4_X1   g124(.A1(KEYINPUT20), .A2(new_n311_), .A3(new_n323_), .A4(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT20), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n305_), .A2(new_n309_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n327_), .B1(new_n313_), .B2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n286_), .A2(new_n309_), .A3(new_n321_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n325_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n267_), .B1(new_n326_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n325_), .ZN(new_n333_));
  AND4_X1   g132(.A1(KEYINPUT20), .A2(new_n311_), .A3(new_n323_), .A4(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n322_), .A2(KEYINPUT95), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT95), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n321_), .A2(new_n336_), .A3(new_n309_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n286_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n333_), .B1(new_n338_), .B2(new_n329_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n334_), .A2(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G64gat), .B(G92gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT32), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n332_), .A2(new_n340_), .A3(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(KEYINPUT94), .B1(new_n326_), .B2(new_n331_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(new_n347_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n266_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n346_), .B1(new_n326_), .B2(new_n331_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT20), .B1(new_n286_), .B2(new_n310_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n313_), .A2(new_n322_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n333_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n311_), .A2(new_n323_), .A3(KEYINPUT20), .A4(new_n325_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n356_), .A2(new_n357_), .A3(new_n345_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n353_), .A2(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n264_), .A2(KEYINPUT33), .ZN(new_n360_));
  AND2_X1   g159(.A1(new_n256_), .A2(new_n263_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n250_), .A2(new_n251_), .A3(new_n255_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n241_), .A2(new_n249_), .A3(new_n252_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n261_), .A3(new_n363_), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n361_), .A2(new_n262_), .B1(new_n364_), .B2(KEYINPUT33), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n359_), .A2(new_n360_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n313_), .B1(new_n367_), .B2(new_n245_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G228gat), .A2(G233gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(G22gat), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT28), .B1(new_n224_), .B2(KEYINPUT29), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT28), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n245_), .A2(new_n374_), .A3(new_n367_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n372_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n373_), .A2(new_n375_), .A3(new_n372_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(G50gat), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(G50gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n378_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n380_), .B1(new_n381_), .B2(new_n376_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n379_), .A2(new_n382_), .A3(KEYINPUT89), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G78gat), .B(G106gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n384_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n379_), .A2(new_n382_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n371_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n385_), .A2(new_n371_), .A3(new_n387_), .ZN(new_n389_));
  OAI22_X1  g188(.A1(new_n352_), .A2(new_n366_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT96), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT97), .B(KEYINPUT27), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n359_), .A2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n353_), .B(KEYINPUT27), .C1(new_n340_), .C2(new_n346_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n394_), .A2(new_n266_), .A3(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n389_), .A2(new_n388_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n385_), .A2(new_n387_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n370_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n385_), .A2(new_n371_), .A3(new_n387_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n402_), .B(KEYINPUT96), .C1(new_n352_), .C2(new_n366_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n392_), .A2(new_n398_), .A3(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT84), .B(G43gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT31), .B(G15gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT30), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n328_), .B(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n253_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n411_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G71gat), .B(G99gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G227gat), .A2(G233gat), .ZN(new_n415_));
  XOR2_X1   g214(.A(new_n414_), .B(new_n415_), .Z(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n412_), .A2(new_n413_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n417_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n408_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n420_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n422_), .A2(new_n407_), .A3(new_n418_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n421_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n402_), .A2(new_n424_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n396_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT98), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT98), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n396_), .A2(new_n402_), .A3(new_n424_), .A4(new_n429_), .ZN(new_n430_));
  AOI22_X1  g229(.A1(new_n404_), .A2(new_n425_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G113gat), .B(G141gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n432_), .B(new_n287_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(new_n268_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT81), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT80), .ZN(new_n437_));
  NOR2_X1   g236(.A1(G29gat), .A2(G36gat), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT73), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G29gat), .A2(G36gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n439_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT73), .B1(new_n443_), .B2(new_n438_), .ZN(new_n444_));
  INV_X1    g243(.A(G43gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n442_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n445_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n380_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n440_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(new_n443_), .A2(new_n438_), .A3(KEYINPUT73), .ZN(new_n451_));
  OAI21_X1  g250(.A(G43gat), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n452_), .A2(G50gat), .A3(new_n446_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n449_), .A2(new_n453_), .ZN(new_n454_));
  OR2_X1    g253(.A1(G15gat), .A2(G22gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G15gat), .A2(G22gat), .ZN(new_n456_));
  INV_X1    g255(.A(G8gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT77), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT77), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G8gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n460_), .A3(G1gat), .ZN(new_n461_));
  AOI221_X4 g260(.A(KEYINPUT78), .B1(new_n455_), .B2(new_n456_), .C1(new_n461_), .C2(KEYINPUT14), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT78), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(KEYINPUT14), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n455_), .A2(new_n456_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(G1gat), .B1(new_n462_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT14), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT77), .B(G8gat), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n468_), .B1(new_n469_), .B2(G1gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n465_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT78), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n464_), .A2(new_n463_), .A3(new_n465_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n202_), .A3(new_n473_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n467_), .A2(G8gat), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(G8gat), .B1(new_n467_), .B2(new_n474_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n454_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  AND3_X1   g276(.A1(new_n472_), .A2(new_n202_), .A3(new_n473_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n202_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n457_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n467_), .A2(G8gat), .A3(new_n474_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT15), .ZN(new_n482_));
  NOR3_X1   g281(.A1(new_n447_), .A2(new_n448_), .A3(new_n380_), .ZN(new_n483_));
  AOI21_X1  g282(.A(G50gat), .B1(new_n452_), .B2(new_n446_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n482_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n449_), .A2(new_n453_), .A3(KEYINPUT15), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n480_), .A2(new_n481_), .A3(new_n485_), .A4(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n437_), .B1(new_n477_), .B2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n475_), .A2(new_n476_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n485_), .A2(new_n486_), .ZN(new_n490_));
  AOI21_X1  g289(.A(KEYINPUT80), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G229gat), .A2(G233gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NOR3_X1   g292(.A1(new_n488_), .A2(new_n491_), .A3(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n489_), .A2(new_n453_), .A3(new_n449_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n492_), .B1(new_n495_), .B2(new_n477_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n436_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n477_), .A2(new_n487_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT80), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n487_), .A2(new_n437_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n492_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n495_), .A2(new_n477_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n493_), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n501_), .A2(new_n435_), .A3(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n497_), .A2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G120gat), .B(G148gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT5), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(G176gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(new_n280_), .ZN(new_n509_));
  XNOR2_X1  g308(.A(KEYINPUT68), .B(KEYINPUT12), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT10), .B(G99gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT64), .B(G106gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(G85gat), .ZN(new_n515_));
  INV_X1    g314(.A(G92gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(KEYINPUT9), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G99gat), .A2(G106gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT6), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT6), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(G99gat), .A3(G106gat), .ZN(new_n523_));
  AND2_X1   g322(.A1(G85gat), .A2(G92gat), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT9), .ZN(new_n525_));
  AOI22_X1  g324(.A1(new_n521_), .A2(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n514_), .A2(new_n519_), .A3(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT66), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT67), .ZN(new_n530_));
  NOR2_X1   g329(.A1(G85gat), .A2(G92gat), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n530_), .B1(new_n524_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n517_), .A2(KEYINPUT67), .A3(new_n518_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n529_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(G99gat), .ZN(new_n535_));
  INV_X1    g334(.A(G106gat), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n536_), .A3(KEYINPUT65), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT7), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n521_), .A2(new_n523_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT7), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n540_), .A2(new_n535_), .A3(new_n536_), .A4(KEYINPUT65), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n538_), .A2(new_n539_), .A3(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n534_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT8), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT8), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n534_), .A2(new_n545_), .A3(new_n542_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n528_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G71gat), .B(G78gat), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G57gat), .B(G64gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(KEYINPUT11), .A3(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n548_), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n550_), .A2(KEYINPUT11), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n551_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n511_), .B1(new_n547_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(G230gat), .ZN(new_n558_));
  INV_X1    g357(.A(G233gat), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n545_), .B1(new_n534_), .B2(new_n542_), .ZN(new_n562_));
  AND3_X1   g361(.A1(new_n534_), .A2(new_n545_), .A3(new_n542_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n556_), .B(new_n527_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n527_), .B1(new_n563_), .B2(new_n562_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n566_), .A2(KEYINPUT68), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n555_), .A3(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n557_), .A2(new_n561_), .A3(new_n564_), .A4(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n564_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n544_), .A2(new_n546_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n556_), .B1(new_n571_), .B2(new_n527_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n560_), .B1(new_n570_), .B2(new_n572_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n569_), .A2(new_n573_), .A3(KEYINPUT69), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT69), .B1(new_n569_), .B2(new_n573_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n509_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT70), .ZN(new_n577_));
  INV_X1    g376(.A(new_n509_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(new_n569_), .A3(new_n573_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT70), .ZN(new_n580_));
  OAI211_X1 g379(.A(new_n580_), .B(new_n509_), .C1(new_n574_), .C2(new_n575_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n577_), .A2(new_n579_), .A3(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT13), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT13), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n577_), .A2(new_n584_), .A3(new_n579_), .A4(new_n581_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n583_), .A2(KEYINPUT71), .A3(new_n585_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT71), .B1(new_n583_), .B2(new_n585_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n505_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT76), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n485_), .A2(new_n486_), .A3(new_n565_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G232gat), .A2(G233gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT34), .Z(new_n592_));
  XOR2_X1   g391(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n547_), .A2(new_n454_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n590_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n592_), .A2(new_n593_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n596_), .A2(new_n597_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n589_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n596_), .A2(new_n597_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(KEYINPUT76), .A3(new_n598_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT74), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n605_), .A2(new_n226_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n226_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(G162gat), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  AOI21_X1  g408(.A(G162gat), .B1(new_n606_), .B2(new_n607_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT36), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n610_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n608_), .A3(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n601_), .A2(new_n603_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n614_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n602_), .A2(new_n617_), .A3(new_n598_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n619_), .A2(KEYINPUT100), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n555_), .B(new_n624_), .Z(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT79), .Z(new_n626_));
  INV_X1    g425(.A(new_n489_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G127gat), .B(G155gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT16), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(G183gat), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(G211gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT17), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n626_), .A2(new_n627_), .ZN(new_n634_));
  AND3_X1   g433(.A1(new_n628_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT17), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n632_), .A2(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n637_), .B1(new_n628_), .B2(new_n634_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n635_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n623_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n431_), .A2(new_n588_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n266_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n202_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT101), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n431_), .A2(new_n588_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT37), .B1(new_n616_), .B2(new_n618_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n611_), .A2(new_n614_), .A3(KEYINPUT75), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT75), .B1(new_n611_), .B2(new_n614_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n651_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n652_), .A2(KEYINPUT37), .A3(new_n618_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n648_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n640_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n647_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n647_), .A2(KEYINPUT99), .A3(new_n656_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n659_), .A2(new_n202_), .A3(new_n644_), .A4(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n661_), .A2(KEYINPUT38), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(KEYINPUT38), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n646_), .B1(new_n662_), .B2(new_n663_), .ZN(G1324gat));
  INV_X1    g463(.A(KEYINPUT39), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n394_), .A2(new_n395_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n643_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n665_), .B1(new_n668_), .B2(G8gat), .ZN(new_n669_));
  AOI211_X1 g468(.A(KEYINPUT39), .B(new_n457_), .C1(new_n643_), .C2(new_n667_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n659_), .A2(new_n660_), .ZN(new_n671_));
  OR2_X1    g470(.A1(new_n666_), .A2(new_n469_), .ZN(new_n672_));
  OAI22_X1  g471(.A1(new_n669_), .A2(new_n670_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g473(.A1(new_n643_), .A2(new_n424_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(G15gat), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT41), .ZN(new_n677_));
  NOR3_X1   g476(.A1(new_n671_), .A2(G15gat), .A3(new_n425_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n677_), .A2(new_n678_), .ZN(G1326gat));
  NAND2_X1  g478(.A1(new_n643_), .A2(new_n397_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G22gat), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n681_), .A2(KEYINPUT102), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(KEYINPUT102), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(KEYINPUT42), .A3(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT42), .B1(new_n682_), .B2(new_n683_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n402_), .A2(G22gat), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT103), .ZN(new_n687_));
  OAI22_X1  g486(.A1(new_n684_), .A2(new_n685_), .B1(new_n671_), .B2(new_n687_), .ZN(G1327gat));
  NAND2_X1  g487(.A1(new_n404_), .A2(new_n425_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n428_), .A2(new_n430_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(new_n692_), .A3(new_n655_), .ZN(new_n693_));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n431_), .B2(new_n654_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n588_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT44), .B1(new_n695_), .B2(new_n640_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n693_), .A2(new_n694_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n588_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n698_), .A2(KEYINPUT44), .A3(new_n699_), .A4(new_n640_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n697_), .A2(new_n644_), .A3(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(G29gat), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT104), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n623_), .B2(new_n640_), .ZN(new_n704_));
  NOR4_X1   g503(.A1(new_n620_), .A2(new_n639_), .A3(new_n622_), .A4(KEYINPUT104), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n647_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n644_), .A2(new_n702_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT105), .ZN(new_n710_));
  OAI22_X1  g509(.A1(new_n701_), .A2(new_n702_), .B1(new_n708_), .B2(new_n710_), .ZN(G1328gat));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n712_), .A2(KEYINPUT46), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n714_));
  NOR4_X1   g513(.A1(new_n431_), .A2(new_n706_), .A3(G36gat), .A4(new_n588_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(new_n667_), .ZN(new_n716_));
  INV_X1    g515(.A(G36gat), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n691_), .A2(new_n717_), .A3(new_n699_), .A4(new_n707_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n718_), .A2(KEYINPUT106), .A3(new_n666_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT45), .B1(new_n716_), .B2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n715_), .A2(new_n714_), .A3(new_n667_), .ZN(new_n721_));
  OAI21_X1  g520(.A(KEYINPUT106), .B1(new_n718_), .B2(new_n666_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT45), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n721_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n713_), .B1(new_n720_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n700_), .A2(new_n667_), .ZN(new_n726_));
  OAI21_X1  g525(.A(G36gat), .B1(new_n726_), .B2(new_n696_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n712_), .A2(KEYINPUT46), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n725_), .A2(new_n727_), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n725_), .B2(new_n727_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1329gat));
  OAI21_X1  g530(.A(new_n445_), .B1(new_n708_), .B2(new_n425_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n700_), .A2(G43gat), .A3(new_n424_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n696_), .ZN(new_n734_));
  XOR2_X1   g533(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(G1330gat));
  NAND4_X1  g535(.A1(new_n697_), .A2(G50gat), .A3(new_n397_), .A4(new_n700_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n380_), .B1(new_n708_), .B2(new_n402_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n737_), .A2(new_n738_), .ZN(G1331gat));
  NOR2_X1   g538(.A1(new_n586_), .A2(new_n587_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n741_), .A2(new_n505_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n691_), .A2(new_n742_), .ZN(new_n743_));
  NOR3_X1   g542(.A1(new_n743_), .A2(new_n640_), .A3(new_n655_), .ZN(new_n744_));
  AOI21_X1  g543(.A(G57gat), .B1(new_n744_), .B2(new_n644_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n743_), .A2(new_n642_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n644_), .A2(G57gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n745_), .B1(new_n746_), .B2(new_n747_), .ZN(G1332gat));
  INV_X1    g547(.A(G64gat), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n667_), .A2(new_n749_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT109), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n744_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT48), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n746_), .A2(new_n667_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n754_), .B2(G64gat), .ZN(new_n755_));
  AOI211_X1 g554(.A(KEYINPUT48), .B(new_n749_), .C1(new_n746_), .C2(new_n667_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n752_), .B1(new_n755_), .B2(new_n756_), .ZN(G1333gat));
  INV_X1    g556(.A(G71gat), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n744_), .A2(new_n758_), .A3(new_n424_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT49), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n746_), .A2(new_n424_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(G71gat), .ZN(new_n762_));
  AOI211_X1 g561(.A(KEYINPUT49), .B(new_n758_), .C1(new_n746_), .C2(new_n424_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(G1334gat));
  INV_X1    g563(.A(G78gat), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n744_), .A2(new_n765_), .A3(new_n397_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n746_), .A2(new_n397_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(G78gat), .ZN(new_n769_));
  AOI211_X1 g568(.A(KEYINPUT50), .B(new_n765_), .C1(new_n746_), .C2(new_n397_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(G1335gat));
  INV_X1    g570(.A(KEYINPUT110), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n698_), .A2(new_n772_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n741_), .A2(new_n505_), .A3(new_n639_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n693_), .A2(new_n694_), .A3(KEYINPUT110), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n773_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  NOR3_X1   g575(.A1(new_n776_), .A2(new_n515_), .A3(new_n266_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n743_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n644_), .A3(new_n707_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n777_), .B1(new_n515_), .B2(new_n779_), .ZN(G1336gat));
  NOR3_X1   g579(.A1(new_n776_), .A2(new_n516_), .A3(new_n666_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n778_), .A2(new_n667_), .A3(new_n707_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n516_), .B2(new_n782_), .ZN(G1337gat));
  OAI21_X1  g582(.A(G99gat), .B1(new_n776_), .B2(new_n425_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n778_), .A2(new_n707_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n424_), .A2(new_n512_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n784_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n784_), .B(new_n788_), .C1(new_n785_), .C2(new_n786_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(G1338gat));
  NAND4_X1  g591(.A1(new_n778_), .A2(new_n513_), .A3(new_n397_), .A4(new_n707_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n698_), .A2(new_n397_), .A3(new_n774_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n795_));
  AND3_X1   g594(.A1(new_n794_), .A2(new_n795_), .A3(G106gat), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n795_), .B1(new_n794_), .B2(G106gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n793_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g598(.A1(new_n667_), .A2(new_n266_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n426_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT57), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n560_), .A2(KEYINPUT114), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n557_), .A2(new_n564_), .A3(new_n568_), .A4(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n568_), .A2(new_n564_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n510_), .B1(new_n565_), .B2(new_n555_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n805_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(KEYINPUT55), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n809_), .B1(new_n813_), .B2(new_n569_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT115), .B1(new_n814_), .B2(new_n578_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT56), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n568_), .B(new_n564_), .C1(new_n572_), .C2(new_n510_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n806_), .B1(new_n817_), .B2(new_n805_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n569_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n808_), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT115), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n820_), .A2(new_n821_), .A3(new_n509_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n815_), .A2(new_n816_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n820_), .A2(KEYINPUT56), .A3(new_n509_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n815_), .A2(KEYINPUT116), .A3(new_n816_), .A4(new_n822_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n505_), .B2(new_n579_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n579_), .ZN(new_n831_));
  AOI211_X1 g630(.A(KEYINPUT113), .B(new_n831_), .C1(new_n497_), .C2(new_n504_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n494_), .A2(new_n434_), .A3(new_n496_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n434_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n493_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n495_), .A2(new_n492_), .A3(new_n477_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n835_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n834_), .A2(new_n838_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n828_), .A2(new_n833_), .B1(new_n582_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n803_), .B1(new_n840_), .B2(new_n623_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n828_), .A2(new_n833_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n839_), .A2(new_n582_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n623_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(KEYINPUT57), .A3(new_n845_), .ZN(new_n846_));
  AND3_X1   g645(.A1(new_n820_), .A2(KEYINPUT56), .A3(new_n509_), .ZN(new_n847_));
  AOI21_X1  g646(.A(KEYINPUT56), .B1(new_n820_), .B2(new_n509_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n501_), .A2(new_n835_), .A3(new_n503_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n836_), .A2(new_n837_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n835_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n849_), .A2(new_n852_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n853_), .A2(KEYINPUT117), .A3(KEYINPUT58), .A4(new_n579_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n816_), .B1(new_n814_), .B2(new_n578_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n826_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n839_), .A2(new_n856_), .A3(KEYINPUT58), .A4(new_n579_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n854_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n839_), .A2(new_n856_), .A3(new_n579_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n654_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  AND3_X1   g663(.A1(new_n860_), .A2(new_n861_), .A3(new_n864_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n861_), .B1(new_n860_), .B2(new_n864_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n841_), .B(new_n846_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n640_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n583_), .A2(new_n585_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n505_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(new_n639_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT112), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n869_), .A2(KEYINPUT112), .A3(new_n870_), .A4(new_n639_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n655_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n875_), .B(new_n876_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n802_), .B1(new_n868_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT59), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n802_), .A2(KEYINPUT59), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n623_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n882_), .A2(KEYINPUT57), .B1(new_n864_), .B2(new_n860_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n639_), .B1(new_n883_), .B2(new_n841_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n873_), .A2(new_n874_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n876_), .B1(new_n885_), .B2(new_n654_), .ZN(new_n886_));
  AOI211_X1 g685(.A(KEYINPUT54), .B(new_n655_), .C1(new_n873_), .C2(new_n874_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n881_), .B1(new_n884_), .B2(new_n888_), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n880_), .A2(G113gat), .A3(new_n505_), .A4(new_n889_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n236_), .B1(new_n879_), .B2(new_n870_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1340gat));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n740_), .B(new_n889_), .C1(new_n878_), .C2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(G120gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n247_), .B1(new_n741_), .B2(KEYINPUT60), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n878_), .B(new_n896_), .C1(KEYINPUT60), .C2(new_n247_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n895_), .A2(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT119), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n895_), .A2(KEYINPUT119), .A3(new_n897_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1341gat));
  NAND4_X1  g701(.A1(new_n880_), .A2(G127gat), .A3(new_n639_), .A4(new_n889_), .ZN(new_n903_));
  AOI21_X1  g702(.A(G127gat), .B1(new_n878_), .B2(new_n639_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n904_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(new_n905_), .ZN(new_n907_));
  AND3_X1   g706(.A1(new_n903_), .A2(new_n906_), .A3(new_n907_), .ZN(G1342gat));
  XNOR2_X1  g707(.A(KEYINPUT121), .B(G134gat), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n880_), .A2(new_n655_), .A3(new_n889_), .A4(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n226_), .B1(new_n879_), .B2(new_n845_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1343gat));
  AOI21_X1  g711(.A(new_n888_), .B1(new_n640_), .B2(new_n867_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n913_), .A2(new_n424_), .A3(new_n402_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n914_), .A2(new_n505_), .A3(new_n800_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT122), .B(G141gat), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(G1344gat));
  NAND3_X1  g716(.A1(new_n914_), .A2(new_n740_), .A3(new_n800_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT123), .B(G148gat), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(G1345gat));
  NAND3_X1  g719(.A1(new_n914_), .A2(new_n639_), .A3(new_n800_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(KEYINPUT61), .B(G155gat), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(KEYINPUT124), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n921_), .B(new_n923_), .ZN(G1346gat));
  AND2_X1   g723(.A1(new_n914_), .A2(new_n800_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n654_), .A2(new_n204_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n914_), .A2(new_n623_), .A3(new_n800_), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n925_), .A2(new_n926_), .B1(new_n927_), .B2(new_n204_), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n884_), .A2(new_n888_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n666_), .A2(new_n644_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n801_), .A2(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n929_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(KEYINPUT125), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n934_), .B1(new_n929_), .B2(new_n931_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(KEYINPUT22), .B(G169gat), .ZN(new_n936_));
  NAND4_X1  g735(.A1(new_n933_), .A2(new_n505_), .A3(new_n935_), .A4(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT62), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n932_), .A2(new_n505_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n938_), .B1(new_n939_), .B2(G169gat), .ZN(new_n940_));
  AOI211_X1 g739(.A(KEYINPUT62), .B(new_n287_), .C1(new_n932_), .C2(new_n505_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n937_), .B1(new_n940_), .B2(new_n941_), .ZN(G1348gat));
  NAND3_X1  g741(.A1(new_n933_), .A2(new_n740_), .A3(new_n935_), .ZN(new_n943_));
  NOR2_X1   g742(.A1(new_n913_), .A2(new_n931_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n741_), .A2(new_n288_), .ZN(new_n945_));
  AOI22_X1  g744(.A1(new_n943_), .A2(new_n288_), .B1(new_n944_), .B2(new_n945_), .ZN(G1349gat));
  AOI21_X1  g745(.A(G183gat), .B1(new_n944_), .B2(new_n639_), .ZN(new_n947_));
  AND2_X1   g746(.A1(new_n933_), .A2(new_n935_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n640_), .A2(new_n294_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n947_), .B1(new_n948_), .B2(new_n949_), .ZN(G1350gat));
  NAND3_X1  g749(.A1(new_n948_), .A2(new_n295_), .A3(new_n623_), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n933_), .A2(new_n655_), .A3(new_n935_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(G190gat), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n951_), .A2(new_n953_), .ZN(G1351gat));
  AOI21_X1  g753(.A(new_n424_), .B1(new_n868_), .B2(new_n877_), .ZN(new_n955_));
  AND3_X1   g754(.A1(new_n955_), .A2(new_n397_), .A3(new_n930_), .ZN(new_n956_));
  NAND4_X1  g755(.A1(new_n956_), .A2(KEYINPUT126), .A3(G197gat), .A4(new_n505_), .ZN(new_n957_));
  NAND4_X1  g756(.A1(new_n955_), .A2(new_n505_), .A3(new_n397_), .A4(new_n930_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n958_), .A2(new_n268_), .ZN(new_n959_));
  INV_X1    g758(.A(KEYINPUT126), .ZN(new_n960_));
  OAI21_X1  g759(.A(new_n960_), .B1(new_n958_), .B2(new_n268_), .ZN(new_n961_));
  AND3_X1   g760(.A1(new_n957_), .A2(new_n959_), .A3(new_n961_), .ZN(G1352gat));
  NAND2_X1  g761(.A1(new_n956_), .A2(new_n740_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(KEYINPUT127), .B(G204gat), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n963_), .B(new_n964_), .ZN(G1353gat));
  XOR2_X1   g764(.A(KEYINPUT63), .B(G211gat), .Z(new_n966_));
  AND3_X1   g765(.A1(new_n956_), .A2(new_n639_), .A3(new_n966_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n956_), .A2(new_n639_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n967_), .B1(new_n968_), .B2(new_n969_), .ZN(G1354gat));
  AOI21_X1  g769(.A(G218gat), .B1(new_n956_), .B2(new_n623_), .ZN(new_n971_));
  AND2_X1   g770(.A1(new_n655_), .A2(G218gat), .ZN(new_n972_));
  AOI21_X1  g771(.A(new_n971_), .B1(new_n956_), .B2(new_n972_), .ZN(G1355gat));
endmodule


