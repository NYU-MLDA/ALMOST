//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n662_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n866_, new_n867_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_, new_n907_, new_n908_;
  XOR2_X1   g000(.A(KEYINPUT25), .B(G183gat), .Z(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT81), .ZN(new_n203_));
  INV_X1    g002(.A(G190gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT26), .ZN(new_n205_));
  OR2_X1    g004(.A1(new_n204_), .A2(KEYINPUT26), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT81), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT25), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n207_), .B1(new_n208_), .B2(G183gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n203_), .A2(new_n205_), .A3(new_n206_), .A4(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n213_), .A2(KEYINPUT24), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(KEYINPUT24), .A3(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n210_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G183gat), .ZN(new_n220_));
  OR3_X1    g019(.A1(new_n220_), .A2(new_n204_), .A3(KEYINPUT23), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT23), .B1(new_n220_), .B2(new_n204_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n222_), .A2(KEYINPUT82), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(KEYINPUT82), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n221_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n221_), .A2(new_n222_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G183gat), .A2(G190gat), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(new_n211_), .ZN(new_n231_));
  OAI22_X1  g030(.A1(new_n219_), .A2(new_n226_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G227gat), .A2(G233gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(G15gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(new_n234_), .B(KEYINPUT30), .Z(new_n235_));
  XNOR2_X1  g034(.A(new_n232_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G127gat), .B(G134gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(G113gat), .B(G120gat), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n238_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT83), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(KEYINPUT83), .A3(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n236_), .B(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G71gat), .B(G99gat), .ZN(new_n247_));
  INV_X1    g046(.A(G43gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(KEYINPUT31), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n246_), .B(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G197gat), .A2(G204gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT87), .B(G197gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n253_), .B1(new_n254_), .B2(G204gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G211gat), .B(G218gat), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT21), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT88), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT88), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n255_), .A2(new_n261_), .A3(new_n258_), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n255_), .A2(KEYINPUT21), .ZN(new_n263_));
  INV_X1    g062(.A(new_n256_), .ZN(new_n264_));
  OR2_X1    g063(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n265_));
  INV_X1    g064(.A(G204gat), .ZN(new_n266_));
  NAND2_X1  g065(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n257_), .B1(G197gat), .B2(G204gat), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n264_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n260_), .A2(new_n262_), .B1(new_n263_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT89), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n270_), .B1(KEYINPUT21), .B2(new_n255_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n262_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n261_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n274_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(KEYINPUT89), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G228gat), .A2(G233gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT86), .ZN(new_n280_));
  OR3_X1    g079(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G141gat), .A2(G148gat), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT2), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n281_), .A2(new_n284_), .A3(new_n285_), .A4(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288_));
  OR2_X1    g087(.A1(G155gat), .A2(G162gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G141gat), .ZN(new_n291_));
  INV_X1    g090(.A(G148gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n288_), .A2(KEYINPUT1), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n289_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n288_), .A2(KEYINPUT1), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n282_), .B(new_n293_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n290_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT29), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n273_), .A2(new_n278_), .A3(new_n280_), .A4(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G78gat), .B(G106gat), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n277_), .A2(new_n299_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n280_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n300_), .A2(new_n302_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT90), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n300_), .A2(KEYINPUT90), .A3(new_n302_), .A4(new_n305_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n300_), .A2(new_n305_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(new_n301_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n308_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n298_), .A2(KEYINPUT29), .ZN(new_n313_));
  XOR2_X1   g112(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(G22gat), .B(G50gat), .Z(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n313_), .A2(new_n315_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n317_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n319_), .B1(new_n317_), .B2(new_n320_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(KEYINPUT85), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT85), .ZN(new_n325_));
  INV_X1    g124(.A(new_n320_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n318_), .B1(new_n326_), .B2(new_n316_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n325_), .B1(new_n327_), .B2(new_n321_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n324_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n312_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT91), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n312_), .A2(new_n329_), .A3(KEYINPUT91), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n311_), .B(new_n306_), .C1(new_n321_), .C2(new_n327_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  XOR2_X1   g135(.A(G8gat), .B(G36gat), .Z(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT96), .ZN(new_n338_));
  XOR2_X1   g137(.A(G64gat), .B(G92gat), .Z(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n273_), .A2(new_n278_), .A3(new_n232_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT94), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n273_), .A2(new_n278_), .A3(KEYINPUT94), .A4(new_n232_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n228_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n225_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(KEYINPUT22), .B(G169gat), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT93), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n212_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(new_n353_), .A3(new_n215_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n221_), .A2(new_n222_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n206_), .A2(new_n205_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n218_), .B(new_n355_), .C1(new_n202_), .C2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n271_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT92), .B(KEYINPUT19), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G226gat), .A2(G233gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n358_), .A2(KEYINPUT20), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n347_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n232_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n271_), .A2(new_n272_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n277_), .A2(KEYINPUT89), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT20), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n354_), .A2(new_n357_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n370_), .B1(new_n371_), .B2(new_n277_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n362_), .B1(new_n369_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n342_), .B1(new_n365_), .B2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n363_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n342_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n376_), .A2(new_n373_), .A3(new_n377_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n243_), .A2(new_n298_), .A3(new_n244_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n241_), .A2(new_n297_), .A3(new_n290_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(KEYINPUT4), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G225gat), .A2(G233gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(KEYINPUT97), .B(KEYINPUT4), .Z(new_n385_));
  NAND4_X1  g184(.A1(new_n243_), .A2(new_n298_), .A3(new_n244_), .A4(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n382_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT98), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n380_), .A2(new_n381_), .A3(new_n383_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT98), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n382_), .A2(new_n390_), .A3(new_n384_), .A4(new_n386_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(G1gat), .B(G29gat), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G85gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT0), .B(G57gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n393_), .B(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT33), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n388_), .A2(new_n389_), .A3(new_n391_), .A4(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT99), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n391_), .A2(new_n389_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n402_), .A2(KEYINPUT99), .A3(new_n388_), .A4(new_n397_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n395_), .ZN(new_n405_));
  AND3_X1   g204(.A1(new_n380_), .A2(new_n381_), .A3(new_n384_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n386_), .A2(new_n383_), .ZN(new_n407_));
  AOI211_X1 g206(.A(new_n405_), .B(new_n406_), .C1(new_n382_), .C2(new_n407_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n388_), .A2(new_n389_), .A3(new_n391_), .A4(new_n405_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n409_), .B2(new_n396_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n379_), .A2(KEYINPUT100), .A3(new_n404_), .A4(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n365_), .A2(new_n374_), .A3(new_n342_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n377_), .B1(new_n376_), .B2(new_n373_), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n404_), .A2(new_n412_), .A3(new_n413_), .A4(new_n410_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT100), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n416_), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n342_), .A2(KEYINPUT32), .ZN(new_n418_));
  OR3_X1    g217(.A1(new_n376_), .A2(new_n418_), .A3(new_n373_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n388_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n395_), .B1(new_n420_), .B2(new_n401_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT104), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n421_), .A2(new_n422_), .A3(new_n409_), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT104), .B(new_n395_), .C1(new_n420_), .C2(new_n401_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n419_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT101), .B(KEYINPUT20), .Z(new_n426_));
  AND3_X1   g225(.A1(new_n358_), .A2(KEYINPUT102), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT102), .B1(new_n358_), .B2(new_n426_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n347_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT103), .B1(new_n430_), .B2(new_n362_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n362_), .B1(new_n347_), .B2(new_n429_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT103), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n369_), .A2(new_n362_), .A3(new_n372_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n431_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n425_), .B1(new_n436_), .B2(new_n418_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n336_), .B1(new_n417_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n423_), .A2(new_n424_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n440_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT27), .B1(new_n412_), .B2(new_n413_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n435_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n443_));
  AOI211_X1 g242(.A(KEYINPUT103), .B(new_n362_), .C1(new_n347_), .C2(new_n429_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n377_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n412_), .A2(KEYINPUT27), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n442_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n441_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n252_), .B1(new_n438_), .B2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n440_), .A2(new_n251_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n336_), .A2(new_n447_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n449_), .A2(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G15gat), .B(G22gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT75), .B(G8gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(G1gat), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n454_), .B1(new_n456_), .B2(KEYINPUT14), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT76), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G1gat), .B(G8gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT76), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n457_), .B(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n459_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n460_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G43gat), .B(G50gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G29gat), .B(G36gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT71), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n468_), .A2(KEYINPUT71), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n467_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G29gat), .B(G36gat), .Z(new_n473_));
  INV_X1    g272(.A(KEYINPUT71), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(new_n469_), .A3(new_n466_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n472_), .A2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n465_), .A2(KEYINPUT78), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(KEYINPUT78), .B1(new_n465_), .B2(new_n478_), .ZN(new_n481_));
  OAI22_X1  g280(.A1(new_n480_), .A2(new_n481_), .B1(new_n478_), .B2(new_n465_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G229gat), .A2(G233gat), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n481_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n479_), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n483_), .B(KEYINPUT79), .Z(new_n488_));
  INV_X1    g287(.A(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n465_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT15), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n470_), .A2(new_n471_), .A3(new_n467_), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n466_), .B1(new_n475_), .B2(new_n469_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n491_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n472_), .A2(KEYINPUT15), .A3(new_n476_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n489_), .B1(new_n490_), .B2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n487_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n485_), .A2(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G113gat), .B(G141gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT80), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G169gat), .B(G197gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n501_), .B(new_n502_), .Z(new_n503_));
  NAND2_X1  g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n482_), .A2(new_n484_), .B1(new_n487_), .B2(new_n497_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n503_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n453_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(G85gat), .ZN(new_n511_));
  INV_X1    g310(.A(G92gat), .ZN(new_n512_));
  NOR3_X1   g311(.A1(new_n511_), .A2(new_n512_), .A3(KEYINPUT9), .ZN(new_n513_));
  XOR2_X1   g312(.A(G85gat), .B(G92gat), .Z(new_n514_));
  AOI21_X1  g313(.A(new_n513_), .B1(new_n514_), .B2(KEYINPUT9), .ZN(new_n515_));
  XNOR2_X1  g314(.A(KEYINPUT10), .B(G99gat), .ZN(new_n516_));
  OR2_X1    g315(.A1(new_n516_), .A2(G106gat), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT6), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT65), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT65), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT6), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n519_), .A2(new_n521_), .A3(G99gat), .A4(G106gat), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G99gat), .A2(G106gat), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n520_), .A2(KEYINPUT6), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n518_), .A2(KEYINPUT65), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n515_), .A2(new_n517_), .A3(new_n522_), .A4(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT66), .ZN(new_n528_));
  INV_X1    g327(.A(G99gat), .ZN(new_n529_));
  INV_X1    g328(.A(G106gat), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT7), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT7), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n528_), .A2(new_n533_), .A3(new_n529_), .A4(new_n530_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n526_), .A2(new_n522_), .A3(new_n532_), .A4(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT8), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n514_), .A2(KEYINPUT67), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n535_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n536_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n527_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G57gat), .B(G64gat), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n543_));
  XOR2_X1   g342(.A(G71gat), .B(G78gat), .Z(new_n544_));
  NAND3_X1  g343(.A1(new_n542_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  OR2_X1    g344(.A1(new_n543_), .A2(new_n544_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n540_), .A2(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n547_), .B(new_n527_), .C1(new_n538_), .C2(new_n539_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(KEYINPUT12), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT12), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n540_), .A2(new_n552_), .A3(new_n548_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT64), .ZN(new_n556_));
  AOI21_X1  g355(.A(KEYINPUT68), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT68), .ZN(new_n558_));
  INV_X1    g357(.A(new_n556_), .ZN(new_n559_));
  AOI211_X1 g358(.A(new_n558_), .B(new_n559_), .C1(new_n551_), .C2(new_n553_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n549_), .A2(new_n550_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n559_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G120gat), .B(G148gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT5), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G176gat), .B(G204gat), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n561_), .A2(new_n563_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n570_));
  OAI22_X1  g369(.A1(new_n569_), .A2(new_n570_), .B1(KEYINPUT69), .B2(KEYINPUT13), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n569_), .A2(new_n570_), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n573_));
  OAI21_X1  g372(.A(new_n571_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(G231gat), .A2(G233gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n465_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(new_n548_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G127gat), .B(G155gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT16), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G183gat), .B(G211gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n579_), .B(new_n580_), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  OR2_X1    g381(.A1(new_n582_), .A2(KEYINPUT17), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(KEYINPUT17), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n577_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n585_), .A2(KEYINPUT77), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT77), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n587_), .B1(new_n577_), .B2(new_n584_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n586_), .B1(new_n585_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G232gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT35), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n496_), .A2(new_n540_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT72), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT72), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n496_), .A2(new_n540_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  OAI22_X1  g401(.A1(new_n540_), .A2(new_n477_), .B1(KEYINPUT35), .B2(new_n593_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n597_), .B1(new_n602_), .B2(new_n604_), .ZN(new_n605_));
  AOI211_X1 g404(.A(new_n596_), .B(new_n603_), .C1(new_n599_), .C2(new_n601_), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT74), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G190gat), .B(G218gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT73), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(G134gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(G162gat), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n613_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n612_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n607_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n615_), .ZN(new_n617_));
  OAI221_X1 g416(.A(KEYINPUT74), .B1(new_n617_), .B2(new_n613_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT37), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n616_), .A2(KEYINPUT37), .A3(new_n618_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n590_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n510_), .A2(new_n574_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(G1gat), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(new_n627_), .A3(new_n440_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT38), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n628_), .B1(KEYINPUT106), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT106), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n630_), .B1(new_n631_), .B2(KEYINPUT38), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n628_), .A2(KEYINPUT106), .A3(new_n629_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n453_), .A2(new_n619_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n574_), .A2(new_n508_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n635_), .A2(new_n590_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT105), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n639_), .A2(new_n440_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n632_), .B(new_n633_), .C1(new_n640_), .C2(new_n627_), .ZN(G1324gat));
  INV_X1    g440(.A(new_n447_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n634_), .A2(new_n642_), .A3(new_n636_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT107), .B1(new_n643_), .B2(G8gat), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(KEYINPUT107), .A3(G8gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n645_), .A2(KEYINPUT39), .A3(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n625_), .A2(new_n447_), .A3(new_n455_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT39), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n648_), .B1(new_n644_), .B2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n647_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n647_), .B2(new_n650_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1325gat));
  INV_X1    g453(.A(G15gat), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n626_), .A2(new_n655_), .A3(new_n252_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n639_), .A2(new_n252_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT41), .B1(new_n657_), .B2(G15gat), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n659_));
  AOI211_X1 g458(.A(new_n659_), .B(new_n655_), .C1(new_n639_), .C2(new_n252_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n656_), .B1(new_n658_), .B2(new_n660_), .ZN(G1326gat));
  INV_X1    g460(.A(G22gat), .ZN(new_n662_));
  INV_X1    g461(.A(new_n336_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n626_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT42), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n639_), .A2(new_n663_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n666_), .B2(G22gat), .ZN(new_n667_));
  AOI211_X1 g466(.A(KEYINPUT42), .B(new_n662_), .C1(new_n639_), .C2(new_n663_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(G1327gat));
  NOR2_X1   g468(.A1(new_n635_), .A2(new_n589_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n671_), .B(new_n623_), .C1(new_n449_), .C2(new_n452_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n418_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n419_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n676_), .A2(new_n416_), .A3(new_n411_), .ZN(new_n677_));
  AOI22_X1  g476(.A1(new_n677_), .A2(new_n336_), .B1(new_n441_), .B2(new_n447_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n451_), .B1(new_n678_), .B2(new_n252_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n671_), .B1(new_n679_), .B2(new_n623_), .ZN(new_n680_));
  OAI211_X1 g479(.A(KEYINPUT44), .B(new_n670_), .C1(new_n673_), .C2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(G29gat), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n439_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n670_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n680_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(new_n672_), .ZN(new_n686_));
  XOR2_X1   g485(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n687_));
  OAI211_X1 g486(.A(new_n681_), .B(new_n683_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n590_), .A2(new_n619_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n574_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n510_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n682_), .B1(new_n692_), .B2(new_n439_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n688_), .A2(new_n693_), .ZN(G1328gat));
  OAI211_X1 g493(.A(new_n642_), .B(new_n681_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G36gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n447_), .A2(G36gat), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n510_), .A2(new_n691_), .A3(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT45), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT46), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n696_), .A2(KEYINPUT46), .A3(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1329gat));
  OAI21_X1  g503(.A(new_n248_), .B1(new_n692_), .B2(new_n251_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n681_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n252_), .A2(G43gat), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n705_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g508(.A1(new_n692_), .A2(G50gat), .A3(new_n336_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n663_), .B(new_n681_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G50gat), .B1(new_n711_), .B2(new_n712_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n710_), .B1(new_n713_), .B2(new_n714_), .ZN(G1331gat));
  INV_X1    g514(.A(G57gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n453_), .A2(new_n508_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(new_n690_), .A3(new_n624_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n718_), .B2(new_n439_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT111), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n590_), .A2(new_n508_), .A3(new_n574_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n634_), .A2(new_n721_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n722_), .A2(new_n716_), .A3(new_n439_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n720_), .A2(new_n723_), .ZN(G1332gat));
  OAI21_X1  g523(.A(G64gat), .B1(new_n722_), .B2(new_n447_), .ZN(new_n725_));
  XOR2_X1   g524(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n726_));
  XNOR2_X1  g525(.A(new_n725_), .B(new_n726_), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n447_), .A2(G64gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n718_), .B2(new_n728_), .ZN(G1333gat));
  OAI21_X1  g528(.A(G71gat), .B1(new_n722_), .B2(new_n251_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT49), .ZN(new_n731_));
  OR2_X1    g530(.A1(new_n251_), .A2(G71gat), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n718_), .B2(new_n732_), .ZN(G1334gat));
  OR3_X1    g532(.A1(new_n718_), .A2(G78gat), .A3(new_n336_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G78gat), .B1(new_n722_), .B2(new_n336_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(KEYINPUT50), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(KEYINPUT50), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n734_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  OAI211_X1 g539(.A(KEYINPUT113), .B(new_n734_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1335gat));
  NOR2_X1   g541(.A1(new_n689_), .A2(new_n574_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n717_), .A2(new_n743_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT114), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n717_), .A2(new_n746_), .A3(new_n743_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G85gat), .B1(new_n748_), .B2(new_n440_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n685_), .A2(new_n672_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n574_), .A2(new_n589_), .A3(new_n508_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n440_), .A2(G85gat), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT115), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n749_), .B1(new_n752_), .B2(new_n754_), .ZN(G1336gat));
  NAND3_X1  g554(.A1(new_n748_), .A2(new_n512_), .A3(new_n642_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n752_), .A2(new_n642_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n757_), .B2(new_n512_), .ZN(G1337gat));
  AOI21_X1  g557(.A(new_n529_), .B1(new_n752_), .B2(new_n252_), .ZN(new_n759_));
  AOI211_X1 g558(.A(new_n251_), .B(new_n516_), .C1(new_n745_), .C2(new_n747_), .ZN(new_n760_));
  OR3_X1    g559(.A1(new_n759_), .A2(new_n760_), .A3(KEYINPUT51), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT51), .B1(new_n759_), .B2(new_n760_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(G1338gat));
  XNOR2_X1  g562(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n663_), .B(new_n751_), .C1(new_n673_), .C2(new_n680_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n766_), .A2(new_n767_), .A3(G106gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n766_), .B2(G106gat), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n768_), .A2(new_n769_), .A3(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n766_), .A2(G106gat), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n772_), .A2(KEYINPUT116), .A3(new_n770_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n336_), .A2(G106gat), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n748_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n765_), .B1(new_n771_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n772_), .A2(KEYINPUT116), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n766_), .A2(new_n767_), .A3(G106gat), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(KEYINPUT52), .A3(new_n779_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n780_), .A2(new_n773_), .A3(new_n775_), .A4(new_n764_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n777_), .A2(new_n781_), .ZN(G1339gat));
  NAND2_X1  g581(.A1(new_n621_), .A2(new_n622_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n574_), .A2(new_n589_), .A3(new_n509_), .A4(new_n783_), .ZN(new_n784_));
  XOR2_X1   g583(.A(KEYINPUT118), .B(KEYINPUT54), .Z(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n784_), .B(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n554_), .A2(KEYINPUT55), .A3(new_n556_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n551_), .A2(new_n559_), .A3(new_n553_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n561_), .B2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT56), .B1(new_n792_), .B2(new_n568_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n569_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT56), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n557_), .A2(new_n560_), .A3(KEYINPUT55), .ZN(new_n796_));
  OAI211_X1 g595(.A(new_n795_), .B(new_n567_), .C1(new_n796_), .C2(new_n790_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n508_), .A2(new_n793_), .A3(new_n794_), .A4(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n488_), .B1(new_n490_), .B2(new_n496_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n506_), .B1(new_n487_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n482_), .A2(new_n488_), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n505_), .A2(new_n506_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n572_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n798_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n619_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n619_), .B1(new_n798_), .B2(new_n803_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT57), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n793_), .A2(new_n794_), .A3(new_n802_), .A4(new_n797_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT58), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT119), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n814_), .A3(new_n623_), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n811_), .A2(new_n812_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n814_), .B1(new_n813_), .B2(new_n623_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n808_), .B(new_n810_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n787_), .B1(new_n819_), .B2(new_n590_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n336_), .A2(new_n447_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n821_), .A2(new_n439_), .A3(new_n251_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n820_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(G113gat), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n824_), .A2(new_n825_), .A3(new_n508_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n820_), .B2(new_n823_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n809_), .B(new_n807_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n813_), .A2(new_n623_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT119), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(new_n816_), .A3(new_n815_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n589_), .B1(new_n829_), .B2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT59), .B(new_n822_), .C1(new_n833_), .C2(new_n787_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n509_), .B1(new_n828_), .B2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n826_), .B1(new_n835_), .B2(new_n825_), .ZN(G1340gat));
  INV_X1    g635(.A(G120gat), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n837_), .B1(new_n574_), .B2(KEYINPUT60), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n839_), .B1(new_n837_), .B2(KEYINPUT60), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n824_), .B(new_n841_), .C1(KEYINPUT120), .C2(new_n838_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n574_), .B1(new_n828_), .B2(new_n834_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(new_n837_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT121), .B(new_n842_), .C1(new_n843_), .C2(new_n837_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(G1341gat));
  INV_X1    g647(.A(G127gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n824_), .A2(new_n849_), .A3(new_n589_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n590_), .B1(new_n828_), .B2(new_n834_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n849_), .ZN(G1342gat));
  AOI21_X1  g651(.A(G134gat), .B1(new_n824_), .B2(new_n619_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n828_), .A2(new_n834_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT122), .B(G134gat), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n783_), .A2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n853_), .B1(new_n854_), .B2(new_n856_), .ZN(G1343gat));
  NAND4_X1  g656(.A1(new_n663_), .A2(new_n440_), .A3(new_n447_), .A4(new_n251_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT123), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n820_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n508_), .ZN(new_n861_));
  XOR2_X1   g660(.A(KEYINPUT124), .B(G141gat), .Z(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1344gat));
  NAND2_X1  g662(.A1(new_n860_), .A2(new_n690_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(new_n864_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g664(.A1(new_n860_), .A2(new_n589_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(KEYINPUT61), .B(G155gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n866_), .B(new_n867_), .ZN(G1346gat));
  INV_X1    g667(.A(G162gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n860_), .A2(new_n869_), .A3(new_n619_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n860_), .A2(new_n623_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n870_), .B1(new_n872_), .B2(new_n869_), .ZN(G1347gat));
  NAND2_X1  g672(.A1(new_n336_), .A2(new_n450_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n642_), .B(new_n875_), .C1(new_n833_), .C2(new_n787_), .ZN(new_n876_));
  OAI21_X1  g675(.A(G169gat), .B1(new_n876_), .B2(new_n509_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT62), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n820_), .A2(new_n447_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n508_), .A2(new_n352_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(KEYINPUT125), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n879_), .A2(new_n875_), .A3(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n878_), .A2(new_n882_), .ZN(G1348gat));
  NOR2_X1   g682(.A1(new_n876_), .A2(new_n574_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(new_n212_), .ZN(G1349gat));
  NAND4_X1  g684(.A1(new_n879_), .A2(new_n202_), .A3(new_n589_), .A4(new_n875_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n220_), .B1(new_n876_), .B2(new_n590_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1350gat));
  OAI21_X1  g687(.A(G190gat), .B1(new_n876_), .B2(new_n783_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n619_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n876_), .B2(new_n890_), .ZN(G1351gat));
  AND2_X1   g690(.A1(new_n441_), .A2(new_n251_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n642_), .B(new_n892_), .C1(new_n833_), .C2(new_n787_), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n508_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g695(.A1(new_n894_), .A2(new_n690_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT126), .B(G204gat), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1353gat));
  NOR2_X1   g698(.A1(new_n893_), .A2(new_n590_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n901_));
  AND2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n900_), .B2(new_n901_), .ZN(G1354gat));
  AND3_X1   g703(.A1(new_n894_), .A2(G218gat), .A3(new_n623_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n893_), .A2(new_n805_), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n906_), .A2(KEYINPUT127), .ZN(new_n907_));
  AOI21_X1  g706(.A(G218gat), .B1(new_n906_), .B2(KEYINPUT127), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n905_), .B1(new_n907_), .B2(new_n908_), .ZN(G1355gat));
endmodule


