//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 0 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT90), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT88), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT89), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT88), .ZN(new_n207_));
  INV_X1    g006(.A(G204gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n207_), .A2(new_n208_), .A3(G197gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n205_), .A2(new_n206_), .A3(KEYINPUT21), .A4(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(G211gat), .B(G218gat), .Z(new_n211_));
  INV_X1    g010(.A(KEYINPUT21), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n211_), .B1(new_n212_), .B2(new_n204_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n210_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n209_), .A2(KEYINPUT21), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n215_), .B1(KEYINPUT88), .B2(new_n204_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(new_n206_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n203_), .B1(new_n214_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n205_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT89), .B1(new_n219_), .B2(new_n215_), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n220_), .A2(KEYINPUT90), .A3(new_n210_), .A4(new_n213_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n218_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n204_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(new_n211_), .A3(KEYINPUT21), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(G169gat), .ZN(new_n227_));
  INV_X1    g026(.A(G183gat), .ZN(new_n228_));
  INV_X1    g027(.A(G190gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT23), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT23), .ZN(new_n231_));
  NAND3_X1  g030(.A1(new_n231_), .A2(G183gat), .A3(G190gat), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n227_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT25), .B(G183gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT75), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT26), .B1(new_n237_), .B2(new_n229_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n229_), .A2(KEYINPUT26), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n236_), .B(new_n238_), .C1(new_n239_), .C2(new_n237_), .ZN(new_n240_));
  OR3_X1    g039(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(G169gat), .ZN(new_n244_));
  INV_X1    g043(.A(G176gat), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n243_), .B(KEYINPUT76), .C1(new_n244_), .C2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT76), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n244_), .A2(new_n245_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n247_), .B1(new_n248_), .B2(new_n242_), .ZN(new_n249_));
  NAND4_X1  g048(.A1(new_n240_), .A2(new_n241_), .A3(new_n246_), .A4(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n232_), .B(KEYINPUT77), .ZN(new_n251_));
  INV_X1    g050(.A(new_n230_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n235_), .B1(new_n250_), .B2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT78), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT78), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n256_), .B(new_n235_), .C1(new_n250_), .C2(new_n253_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n202_), .B1(new_n225_), .B2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G226gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT19), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT26), .B(G190gat), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n233_), .B1(new_n236_), .B2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n263_), .A2(new_n241_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n227_), .B1(new_n253_), .B2(new_n234_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT96), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(KEYINPUT96), .B(new_n227_), .C1(new_n253_), .C2(new_n234_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n266_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n224_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n272_), .B1(new_n218_), .B2(new_n221_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n261_), .B1(new_n271_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n259_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(KEYINPUT97), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n261_), .B(KEYINPUT95), .Z(new_n277_));
  OAI21_X1  g076(.A(KEYINPUT20), .B1(new_n271_), .B2(new_n273_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n225_), .A2(new_n258_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n277_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT97), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n259_), .A2(new_n274_), .A3(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n276_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G8gat), .B(G36gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n284_), .B(KEYINPUT18), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G64gat), .B(G92gat), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n285_), .B(new_n286_), .Z(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n283_), .A2(new_n288_), .ZN(new_n289_));
  NAND4_X1  g088(.A1(new_n276_), .A2(new_n287_), .A3(new_n280_), .A4(new_n282_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT27), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NOR3_X1   g090(.A1(new_n278_), .A2(new_n279_), .A3(new_n277_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n261_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n273_), .A2(new_n265_), .A3(new_n267_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n293_), .B1(new_n259_), .B2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n288_), .B1(new_n292_), .B2(new_n295_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n290_), .A2(KEYINPUT27), .A3(new_n296_), .ZN(new_n297_));
  NOR2_X1   g096(.A1(new_n291_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n255_), .A2(KEYINPUT30), .A3(new_n257_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT30), .B1(new_n255_), .B2(new_n257_), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT79), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT30), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n258_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT79), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n305_), .A3(new_n299_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G71gat), .B(G99gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(G43gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G227gat), .A2(G233gat), .ZN(new_n309_));
  INV_X1    g108(.A(G15gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n308_), .B(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n302_), .A2(new_n306_), .A3(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(KEYINPUT79), .B(new_n312_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT83), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G127gat), .B(G134gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G113gat), .B(G120gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n320_), .A2(new_n321_), .ZN(new_n323_));
  NOR2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT83), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n314_), .A2(new_n328_), .A3(new_n315_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n317_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  INV_X1    g130(.A(G141gat), .ZN(new_n332_));
  INV_X1    g131(.A(G148gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(G155gat), .A2(G162gat), .ZN(new_n335_));
  XOR2_X1   g134(.A(new_n335_), .B(KEYINPUT84), .Z(new_n336_));
  NAND2_X1  g135(.A1(G155gat), .A2(G162gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n336_), .B1(KEYINPUT1), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(KEYINPUT1), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT85), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n331_), .B(new_n334_), .C1(new_n338_), .C2(new_n340_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n334_), .A2(KEYINPUT3), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n334_), .A2(KEYINPUT3), .ZN(new_n343_));
  AOI22_X1  g142(.A1(KEYINPUT86), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n344_));
  NOR2_X1   g143(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n342_), .B(new_n343_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n344_), .A2(new_n345_), .ZN(new_n347_));
  OAI211_X1 g146(.A(new_n336_), .B(new_n337_), .C1(new_n346_), .C2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n341_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n324_), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n341_), .B(new_n348_), .C1(new_n322_), .C2(new_n323_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n351_), .A3(KEYINPUT4), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT4), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(new_n324_), .A3(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n352_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G1gat), .B(G29gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n359_), .B(G85gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(KEYINPUT0), .B(G57gat), .ZN(new_n361_));
  XOR2_X1   g160(.A(new_n360_), .B(new_n361_), .Z(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n357_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n358_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n356_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n362_), .B1(new_n367_), .B2(new_n364_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n316_), .A2(KEYINPUT83), .A3(new_n326_), .ZN(new_n371_));
  AND3_X1   g170(.A1(new_n330_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT94), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n341_), .A2(new_n374_), .A3(new_n348_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n375_), .A2(KEYINPUT28), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(KEYINPUT28), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G22gat), .B(G50gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n376_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n349_), .A2(KEYINPUT29), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G228gat), .A2(G233gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(new_n385_), .B(KEYINPUT87), .Z(new_n386_));
  NAND3_X1  g185(.A1(new_n225_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G78gat), .B(G106gat), .ZN(new_n388_));
  XOR2_X1   g187(.A(new_n388_), .B(KEYINPUT91), .Z(new_n389_));
  INV_X1    g188(.A(new_n386_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n374_), .B1(new_n341_), .B2(new_n348_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n390_), .B1(new_n273_), .B2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n387_), .A2(new_n389_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT92), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n387_), .A2(new_n392_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n389_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT92), .ZN(new_n398_));
  NAND4_X1  g197(.A1(new_n387_), .A2(new_n392_), .A3(new_n398_), .A4(new_n389_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n383_), .A2(new_n394_), .A3(new_n397_), .A4(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n393_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(KEYINPUT93), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT93), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n395_), .A2(new_n403_), .A3(new_n396_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n401_), .B1(new_n402_), .B2(new_n404_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n373_), .B(new_n400_), .C1(new_n405_), .C2(new_n383_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n403_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n408_));
  AOI211_X1 g207(.A(KEYINPUT93), .B(new_n389_), .C1(new_n387_), .C2(new_n392_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n393_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(new_n382_), .A3(new_n381_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n373_), .B1(new_n411_), .B2(new_n400_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n298_), .B(new_n372_), .C1(new_n407_), .C2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n330_), .A2(new_n371_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n407_), .A2(new_n412_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n298_), .A2(new_n370_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n416_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n400_), .B1(new_n405_), .B2(new_n383_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(KEYINPUT94), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n406_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n287_), .A2(KEYINPUT32), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n276_), .A2(new_n280_), .A3(new_n282_), .A4(new_n423_), .ZN(new_n424_));
  OAI211_X1 g223(.A(KEYINPUT32), .B(new_n287_), .C1(new_n292_), .C2(new_n295_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n369_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT99), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n289_), .A2(new_n290_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(KEYINPUT98), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT33), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n368_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n350_), .A2(new_n357_), .A3(new_n351_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n433_), .B(new_n363_), .C1(new_n355_), .C2(new_n357_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n368_), .A2(new_n431_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n432_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT98), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n289_), .A2(new_n437_), .A3(new_n290_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n430_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n422_), .A2(new_n428_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n414_), .B1(new_n419_), .B2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G113gat), .B(G141gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G169gat), .B(G197gat), .ZN(new_n443_));
  XOR2_X1   g242(.A(new_n442_), .B(new_n443_), .Z(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(G15gat), .B(G22gat), .Z(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(G1gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT67), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G1gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n449_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(G8gat), .ZN(new_n453_));
  AOI21_X1  g252(.A(KEYINPUT68), .B1(new_n453_), .B2(KEYINPUT14), .ZN(new_n454_));
  INV_X1    g253(.A(G8gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT68), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT14), .ZN(new_n458_));
  NOR3_X1   g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n447_), .B1(new_n454_), .B2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G1gat), .B(G8gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n457_), .B1(new_n456_), .B2(new_n458_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT67), .B(G1gat), .ZN(new_n465_));
  OAI211_X1 g264(.A(KEYINPUT68), .B(KEYINPUT14), .C1(new_n465_), .C2(new_n455_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n467_), .A2(new_n447_), .A3(new_n461_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G29gat), .B(G36gat), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G43gat), .B(G50gat), .Z(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G43gat), .B(G50gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n469_), .A2(new_n473_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n472_), .A2(KEYINPUT15), .A3(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT15), .B1(new_n472_), .B2(new_n474_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n463_), .A2(new_n468_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n472_), .A2(new_n474_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n461_), .B1(new_n467_), .B2(new_n447_), .ZN(new_n480_));
  AOI211_X1 g279(.A(new_n446_), .B(new_n462_), .C1(new_n464_), .C2(new_n466_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n479_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G229gat), .A2(G233gat), .ZN(new_n483_));
  AND3_X1   g282(.A1(new_n478_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n479_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n463_), .A2(new_n485_), .A3(new_n468_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n483_), .B1(new_n486_), .B2(new_n482_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n445_), .B1(new_n484_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(KEYINPUT72), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT72), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n490_), .B(new_n445_), .C1(new_n484_), .C2(new_n487_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n483_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n485_), .B1(new_n463_), .B2(new_n468_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n480_), .A2(new_n481_), .A3(new_n479_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n493_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n478_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n444_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT73), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n496_), .A2(KEYINPUT73), .A3(new_n497_), .A4(new_n444_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT74), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n492_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n503_), .B1(new_n492_), .B2(new_n502_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  XOR2_X1   g305(.A(KEYINPUT10), .B(G99gat), .Z(new_n507_));
  INV_X1    g306(.A(G106gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT6), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT6), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(G99gat), .A3(G106gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n511_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G85gat), .A2(G92gat), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n515_), .A2(KEYINPUT9), .ZN(new_n516_));
  INV_X1    g315(.A(G85gat), .ZN(new_n517_));
  INV_X1    g316(.A(G92gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(KEYINPUT9), .A3(new_n515_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n509_), .A2(new_n514_), .A3(new_n516_), .A4(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n519_), .A2(new_n515_), .ZN(new_n522_));
  NOR4_X1   g321(.A1(KEYINPUT64), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT64), .ZN(new_n524_));
  NOR2_X1   g323(.A1(G99gat), .A2(G106gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT7), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n524_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(G99gat), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n508_), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n511_), .A2(new_n513_), .B1(new_n530_), .B2(KEYINPUT7), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n522_), .B1(new_n528_), .B2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n521_), .B1(new_n532_), .B2(KEYINPUT8), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT64), .B1(new_n530_), .B2(KEYINPUT7), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n530_), .A2(KEYINPUT7), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n525_), .A2(new_n524_), .A3(new_n526_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n534_), .A2(new_n514_), .A3(new_n535_), .A4(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n522_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT8), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n477_), .B1(new_n533_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G232gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT34), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT35), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n539_), .A2(new_n540_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n532_), .A2(KEYINPUT8), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(new_n479_), .A4(new_n521_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n542_), .A2(new_n547_), .A3(new_n550_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n545_), .A2(new_n546_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G190gat), .B(G218gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G134gat), .B(G162gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n554_), .B(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(KEYINPUT36), .ZN(new_n557_));
  INV_X1    g356(.A(new_n552_), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n542_), .A2(new_n558_), .A3(new_n547_), .A4(new_n550_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n553_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT66), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n556_), .B(KEYINPUT36), .Z(new_n562_));
  INV_X1    g361(.A(new_n553_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n559_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n562_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT37), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n561_), .A2(KEYINPUT37), .A3(new_n565_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G71gat), .B(G78gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G57gat), .B(G64gat), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(KEYINPUT11), .B2(new_n573_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n573_), .A2(KEYINPUT11), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n573_), .A2(new_n572_), .A3(KEYINPUT11), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n533_), .B2(new_n541_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n548_), .A2(new_n549_), .A3(new_n521_), .A4(new_n578_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(KEYINPUT12), .A3(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT12), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n579_), .B(new_n583_), .C1(new_n533_), .C2(new_n541_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G230gat), .A2(G233gat), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n580_), .A2(new_n581_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n586_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  XOR2_X1   g390(.A(G120gat), .B(G148gat), .Z(new_n592_));
  XNOR2_X1  g391(.A(G176gat), .B(G204gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT65), .B(KEYINPUT5), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n591_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n587_), .A2(new_n590_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT13), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n597_), .A2(KEYINPUT13), .A3(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605_));
  XOR2_X1   g404(.A(new_n578_), .B(new_n605_), .Z(new_n606_));
  NAND2_X1  g405(.A1(new_n463_), .A2(new_n468_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(G127gat), .B(G155gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT16), .ZN(new_n611_));
  XOR2_X1   g410(.A(G183gat), .B(G211gat), .Z(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(KEYINPUT71), .B(KEYINPUT17), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n609_), .A2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(KEYINPUT70), .B(KEYINPUT17), .Z(new_n617_));
  AOI211_X1 g416(.A(new_n613_), .B(new_n617_), .C1(new_n608_), .C2(KEYINPUT69), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n608_), .A2(KEYINPUT69), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n616_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n604_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n571_), .A2(new_n622_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n441_), .A2(new_n506_), .A3(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(new_n369_), .A3(new_n465_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT38), .ZN(new_n626_));
  INV_X1    g425(.A(new_n566_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT100), .B1(new_n441_), .B2(new_n627_), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n422_), .A2(new_n428_), .A3(new_n439_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n291_), .A2(new_n297_), .A3(new_n369_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n415_), .B1(new_n422_), .B2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n413_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT100), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n633_), .A3(new_n566_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n506_), .A2(new_n604_), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n628_), .A2(new_n634_), .A3(new_n635_), .A4(new_n620_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G1gat), .B1(new_n636_), .B2(new_n370_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n626_), .A2(new_n637_), .ZN(G1324gat));
  INV_X1    g437(.A(new_n298_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n624_), .A2(new_n455_), .A3(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT101), .B(KEYINPUT39), .ZN(new_n641_));
  OAI211_X1 g440(.A(G8gat), .B(new_n641_), .C1(new_n636_), .C2(new_n298_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n632_), .A2(new_n566_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n621_), .B1(new_n644_), .B2(KEYINPUT100), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n645_), .A2(new_n635_), .A3(new_n639_), .A4(new_n634_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n641_), .B1(new_n646_), .B2(G8gat), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n640_), .B1(new_n643_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(KEYINPUT40), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n651_), .B(new_n640_), .C1(new_n643_), .C2(new_n647_), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n649_), .A2(new_n650_), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n650_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1325gat));
  OAI21_X1  g454(.A(G15gat), .B1(new_n636_), .B2(new_n415_), .ZN(new_n656_));
  XOR2_X1   g455(.A(new_n656_), .B(KEYINPUT41), .Z(new_n657_));
  NAND3_X1  g456(.A1(new_n624_), .A2(new_n310_), .A3(new_n416_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1326gat));
  OAI21_X1  g458(.A(G22gat), .B1(new_n636_), .B2(new_n422_), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT42), .ZN(new_n661_));
  INV_X1    g460(.A(G22gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n624_), .A2(new_n662_), .A3(new_n417_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(G1327gat));
  NOR2_X1   g463(.A1(new_n441_), .A2(new_n506_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n621_), .A2(new_n627_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n666_), .A2(new_n604_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(new_n668_));
  OR3_X1    g467(.A1(new_n668_), .A2(G29gat), .A3(new_n370_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n632_), .A2(new_n570_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n671_));
  OAI21_X1  g470(.A(KEYINPUT43), .B1(new_n571_), .B2(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n620_), .B1(new_n670_), .B2(new_n672_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n632_), .A2(new_n671_), .A3(KEYINPUT43), .A4(new_n570_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n635_), .A3(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT44), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n673_), .A2(KEYINPUT44), .A3(new_n635_), .A4(new_n674_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n369_), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT105), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G29gat), .B1(new_n679_), .B2(new_n680_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n669_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT106), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n685_), .B(new_n669_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1328gat));
  NAND3_X1  g486(.A1(new_n677_), .A2(new_n639_), .A3(new_n678_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G36gat), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n298_), .A2(G36gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n665_), .A2(new_n667_), .A3(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n691_), .B(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n689_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT46), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT108), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n693_), .B1(new_n688_), .B2(G36gat), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n698_), .A2(new_n699_), .A3(KEYINPUT46), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n698_), .A2(KEYINPUT109), .A3(KEYINPUT46), .ZN(new_n701_));
  AOI21_X1  g500(.A(KEYINPUT109), .B1(new_n698_), .B2(KEYINPUT46), .ZN(new_n702_));
  OAI22_X1  g501(.A1(new_n697_), .A2(new_n700_), .B1(new_n701_), .B2(new_n702_), .ZN(G1329gat));
  NAND3_X1  g502(.A1(new_n677_), .A2(new_n416_), .A3(new_n678_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G43gat), .ZN(new_n705_));
  OR3_X1    g504(.A1(new_n668_), .A2(G43gat), .A3(new_n415_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT47), .Z(G1330gat));
  AND2_X1   g507(.A1(new_n677_), .A2(new_n678_), .ZN(new_n709_));
  INV_X1    g508(.A(G50gat), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n422_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n665_), .A2(new_n417_), .A3(new_n667_), .ZN(new_n712_));
  AOI22_X1  g511(.A1(new_n709_), .A2(new_n711_), .B1(new_n710_), .B2(new_n712_), .ZN(G1331gat));
  INV_X1    g512(.A(new_n506_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n604_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n645_), .A2(new_n634_), .A3(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(G57gat), .B1(new_n717_), .B2(new_n370_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n571_), .A2(new_n604_), .A3(new_n620_), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT110), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(new_n506_), .A3(new_n632_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n370_), .A2(G57gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(G1332gat));
  OAI21_X1  g522(.A(G64gat), .B1(new_n717_), .B2(new_n298_), .ZN(new_n724_));
  XOR2_X1   g523(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n298_), .A2(G64gat), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n721_), .B2(new_n727_), .ZN(G1333gat));
  OAI21_X1  g527(.A(G71gat), .B1(new_n717_), .B2(new_n415_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT49), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n415_), .A2(G71gat), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n730_), .B1(new_n721_), .B2(new_n731_), .ZN(G1334gat));
  OAI21_X1  g531(.A(G78gat), .B1(new_n717_), .B2(new_n422_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT50), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n422_), .A2(G78gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n721_), .B2(new_n735_), .ZN(G1335gat));
  AND2_X1   g535(.A1(new_n673_), .A2(new_n674_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n716_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n370_), .ZN(new_n739_));
  NOR4_X1   g538(.A1(new_n441_), .A2(new_n714_), .A3(new_n715_), .A4(new_n666_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(new_n517_), .A3(new_n369_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1336gat));
  OAI21_X1  g541(.A(G92gat), .B1(new_n738_), .B2(new_n298_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n740_), .A2(new_n518_), .A3(new_n639_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT112), .ZN(G1337gat));
  OAI21_X1  g545(.A(G99gat), .B1(new_n738_), .B2(new_n415_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n416_), .A2(new_n507_), .ZN(new_n748_));
  AOI22_X1  g547(.A1(new_n740_), .A2(new_n748_), .B1(KEYINPUT113), .B2(KEYINPUT51), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(KEYINPUT113), .A2(KEYINPUT51), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n750_), .B(new_n751_), .Z(G1338gat));
  NAND3_X1  g551(.A1(new_n740_), .A2(new_n508_), .A3(new_n417_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n737_), .A2(new_n417_), .A3(new_n716_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT52), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n755_), .A3(G106gat), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n755_), .B1(new_n754_), .B2(G106gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n753_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT53), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n753_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1339gat));
  NOR2_X1   g562(.A1(new_n417_), .A2(new_n639_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n415_), .A2(new_n370_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n493_), .B1(new_n486_), .B2(new_n482_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n494_), .A2(new_n483_), .ZN(new_n768_));
  AOI211_X1 g567(.A(new_n444_), .B(new_n767_), .C1(new_n478_), .C2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  AND3_X1   g569(.A1(new_n770_), .A2(new_n502_), .A3(new_n599_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT115), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n587_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n589_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT115), .B1(new_n775_), .B2(KEYINPUT55), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(KEYINPUT55), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n582_), .A2(new_n589_), .A3(new_n584_), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n774_), .A2(new_n776_), .A3(new_n777_), .A4(new_n778_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n596_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT56), .B1(new_n779_), .B2(new_n596_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n771_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT58), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI211_X1 g583(.A(KEYINPUT58), .B(new_n771_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n784_), .A2(new_n570_), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT55), .B1(new_n585_), .B2(new_n586_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n777_), .B(new_n778_), .C1(new_n787_), .C2(new_n772_), .ZN(new_n788_));
  NOR3_X1   g587(.A1(new_n775_), .A2(KEYINPUT115), .A3(KEYINPUT55), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n596_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n779_), .A2(KEYINPUT56), .A3(new_n596_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n599_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n492_), .A2(new_n502_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT74), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n492_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n796_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n779_), .A2(KEYINPUT116), .A3(KEYINPUT56), .A4(new_n596_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n795_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n600_), .A2(new_n502_), .A3(new_n770_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n627_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n786_), .B1(new_n804_), .B2(KEYINPUT57), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n780_), .A2(new_n781_), .A3(KEYINPUT116), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n801_), .B(new_n599_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n803_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n808_), .A2(KEYINPUT57), .A3(new_n566_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(KEYINPUT117), .B1(new_n805_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n808_), .A2(new_n566_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n809_), .A4(new_n786_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n811_), .A2(new_n621_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n571_), .A2(new_n818_), .A3(new_n622_), .A4(new_n506_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT114), .ZN(new_n820_));
  OR2_X1    g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n820_), .ZN(new_n822_));
  OAI21_X1  g621(.A(KEYINPUT54), .B1(new_n623_), .B2(new_n714_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n766_), .B1(new_n817_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(G113gat), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n714_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n825_), .B2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n824_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n814_), .A2(new_n809_), .A3(new_n786_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n620_), .B1(new_n832_), .B2(KEYINPUT117), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n831_), .B1(new_n833_), .B2(new_n816_), .ZN(new_n834_));
  OAI211_X1 g633(.A(KEYINPUT118), .B(KEYINPUT59), .C1(new_n834_), .C2(new_n766_), .ZN(new_n835_));
  AOI21_X1  g634(.A(KEYINPUT57), .B1(new_n808_), .B2(new_n566_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n784_), .A2(new_n570_), .A3(new_n785_), .ZN(new_n837_));
  OAI21_X1  g636(.A(KEYINPUT119), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n839_), .B(new_n786_), .C1(new_n804_), .C2(KEYINPUT57), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n838_), .A2(new_n809_), .A3(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n621_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT120), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT120), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n841_), .A2(new_n844_), .A3(new_n621_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n824_), .A3(new_n845_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n766_), .A2(KEYINPUT59), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n830_), .A2(new_n835_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n848_), .A2(new_n714_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n827_), .B1(new_n849_), .B2(new_n826_), .ZN(G1340gat));
  INV_X1    g649(.A(KEYINPUT121), .ZN(new_n851_));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n848_), .B2(new_n604_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n825_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n852_), .A2(KEYINPUT60), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT60), .ZN(new_n856_));
  AOI21_X1  g655(.A(G120gat), .B1(new_n604_), .B2(new_n856_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n854_), .A2(new_n855_), .A3(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n851_), .B1(new_n853_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n858_), .ZN(new_n860_));
  AOI221_X4 g659(.A(new_n715_), .B1(new_n846_), .B2(new_n847_), .C1(new_n830_), .C2(new_n835_), .ZN(new_n861_));
  OAI211_X1 g660(.A(KEYINPUT121), .B(new_n860_), .C1(new_n861_), .C2(new_n852_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(G1341gat));
  INV_X1    g662(.A(G127gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n825_), .A2(new_n864_), .A3(new_n620_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n848_), .A2(new_n620_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n864_), .ZN(G1342gat));
  AOI21_X1  g666(.A(G134gat), .B1(new_n825_), .B2(new_n627_), .ZN(new_n868_));
  XOR2_X1   g667(.A(new_n868_), .B(KEYINPUT122), .Z(new_n869_));
  AND2_X1   g668(.A1(new_n570_), .A2(G134gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n869_), .B1(new_n848_), .B2(new_n870_), .ZN(G1343gat));
  NAND2_X1  g670(.A1(new_n417_), .A2(new_n415_), .ZN(new_n872_));
  OR4_X1    g671(.A1(new_n370_), .A2(new_n834_), .A3(new_n639_), .A4(new_n872_), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n873_), .A2(new_n506_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(new_n332_), .ZN(G1344gat));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n715_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(new_n333_), .ZN(G1345gat));
  NOR2_X1   g676(.A1(new_n873_), .A2(new_n621_), .ZN(new_n878_));
  XOR2_X1   g677(.A(KEYINPUT61), .B(G155gat), .Z(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1346gat));
  OAI21_X1  g679(.A(G162gat), .B1(new_n873_), .B2(new_n571_), .ZN(new_n881_));
  OR2_X1    g680(.A1(new_n566_), .A2(G162gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n881_), .B1(new_n873_), .B2(new_n882_), .ZN(G1347gat));
  XOR2_X1   g682(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n884_));
  NAND3_X1  g683(.A1(new_n639_), .A2(new_n370_), .A3(new_n416_), .ZN(new_n885_));
  XOR2_X1   g684(.A(new_n885_), .B(KEYINPUT123), .Z(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n417_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n846_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n714_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n884_), .B1(new_n890_), .B2(KEYINPUT22), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(new_n244_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n890_), .A2(new_n884_), .ZN(new_n893_));
  OAI211_X1 g692(.A(G169gat), .B(new_n884_), .C1(new_n890_), .C2(KEYINPUT22), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n892_), .A2(new_n893_), .A3(new_n894_), .ZN(G1348gat));
  AOI21_X1  g694(.A(G176gat), .B1(new_n889_), .B2(new_n604_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n834_), .A2(new_n417_), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n887_), .A2(new_n245_), .A3(new_n715_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n896_), .B1(new_n897_), .B2(new_n898_), .ZN(G1349gat));
  INV_X1    g698(.A(new_n889_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n900_), .A2(new_n236_), .A3(new_n621_), .ZN(new_n901_));
  NOR4_X1   g700(.A1(new_n834_), .A2(new_n417_), .A3(new_n621_), .A4(new_n887_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903_));
  OR2_X1    g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(G183gat), .B1(new_n902_), .B2(new_n903_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n901_), .B1(new_n904_), .B2(new_n905_), .ZN(G1350gat));
  OAI21_X1  g705(.A(G190gat), .B1(new_n900_), .B2(new_n571_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n889_), .A2(new_n262_), .A3(new_n627_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1351gat));
  INV_X1    g708(.A(new_n834_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n872_), .A2(new_n369_), .A3(new_n298_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n714_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g714(.A1(new_n912_), .A2(new_n715_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(KEYINPUT126), .B(G204gat), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n916_), .B(new_n917_), .ZN(G1353gat));
  NAND2_X1  g717(.A1(new_n913_), .A2(new_n620_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  AND2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n919_), .A2(new_n920_), .A3(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n919_), .B2(new_n920_), .ZN(G1354gat));
  AND3_X1   g722(.A1(new_n913_), .A2(G218gat), .A3(new_n570_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n912_), .A2(new_n566_), .ZN(new_n925_));
  OR2_X1    g724(.A1(new_n925_), .A2(KEYINPUT127), .ZN(new_n926_));
  AOI21_X1  g725(.A(G218gat), .B1(new_n925_), .B2(KEYINPUT127), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n924_), .B1(new_n926_), .B2(new_n927_), .ZN(G1355gat));
endmodule


