//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 1 0 1 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n570_, new_n571_, new_n572_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n813_, new_n814_,
    new_n815_, new_n817_, new_n818_, new_n819_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n889_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT23), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(G183gat), .B2(G190gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT22), .B(G169gat), .Z(new_n212_));
  OAI21_X1  g011(.A(new_n211_), .B1(G176gat), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G169gat), .ZN(new_n214_));
  INV_X1    g013(.A(G176gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(KEYINPUT24), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT25), .B(G183gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT26), .B(G190gat), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n216_), .A2(KEYINPUT24), .A3(new_n210_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n208_), .A3(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n213_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G211gat), .B(G218gat), .Z(new_n224_));
  XOR2_X1   g023(.A(KEYINPUT88), .B(G197gat), .Z(new_n225_));
  INV_X1    g024(.A(G204gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT21), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(G197gat), .B2(G204gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n224_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  MUX2_X1   g029(.A(G197gat), .B(new_n225_), .S(G204gat), .Z(new_n231_));
  OAI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(KEYINPUT21), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n231_), .A2(KEYINPUT21), .A3(new_n224_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n223_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT83), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT22), .B1(new_n236_), .B2(new_n214_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n214_), .A2(KEYINPUT22), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n215_), .B(new_n237_), .C1(new_n238_), .C2(new_n236_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n211_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(new_n222_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n235_), .B(KEYINPUT20), .C1(new_n241_), .C2(new_n234_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G226gat), .A2(G233gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT19), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT20), .B1(new_n223_), .B2(new_n234_), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n241_), .A2(new_n234_), .ZN(new_n247_));
  NOR3_X1   g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n244_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n206_), .B1(new_n245_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n248_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n242_), .A2(new_n244_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n250_), .A2(new_n205_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT27), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n246_), .A2(new_n247_), .ZN(new_n256_));
  MUX2_X1   g055(.A(new_n242_), .B(new_n256_), .S(new_n244_), .Z(new_n257_));
  XOR2_X1   g056(.A(new_n205_), .B(KEYINPUT94), .Z(new_n258_));
  OAI211_X1 g057(.A(new_n252_), .B(KEYINPUT27), .C1(new_n257_), .C2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  XOR2_X1   g059(.A(G127gat), .B(G134gat), .Z(new_n261_));
  XOR2_X1   g060(.A(G113gat), .B(G120gat), .Z(new_n262_));
  XOR2_X1   g061(.A(new_n261_), .B(new_n262_), .Z(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT85), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  AND2_X1   g064(.A1(G141gat), .A2(G148gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n267_), .B1(KEYINPUT1), .B2(new_n268_), .ZN(new_n269_));
  OR2_X1    g068(.A1(new_n268_), .A2(KEYINPUT1), .ZN(new_n270_));
  AOI211_X1 g069(.A(new_n265_), .B(new_n266_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT3), .ZN(new_n273_));
  AOI22_X1  g072(.A1(KEYINPUT2), .A2(new_n266_), .B1(new_n265_), .B2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(KEYINPUT2), .B2(new_n266_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT87), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n276_), .B1(new_n265_), .B2(new_n273_), .ZN(new_n277_));
  OAI211_X1 g076(.A(KEYINPUT87), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n275_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n267_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n268_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n272_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n264_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT91), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G225gat), .A2(G233gat), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n282_), .A2(new_n263_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT91), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n264_), .A2(new_n287_), .A3(new_n282_), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .A4(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT92), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n288_), .A2(new_n286_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n292_), .A2(KEYINPUT92), .A3(new_n285_), .A4(new_n284_), .ZN(new_n293_));
  AOI21_X1  g092(.A(KEYINPUT4), .B1(new_n264_), .B2(new_n282_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n284_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n295_), .B2(KEYINPUT4), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n291_), .B(new_n293_), .C1(new_n296_), .C2(new_n285_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G29gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(G85gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT0), .B(G57gat), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n299_), .B(new_n300_), .Z(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n304_), .B1(new_n292_), .B2(new_n284_), .ZN(new_n305_));
  OAI211_X1 g104(.A(G225gat), .B(G233gat), .C1(new_n305_), .C2(new_n294_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n291_), .A2(new_n293_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n306_), .A2(new_n307_), .A3(new_n301_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n303_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT93), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT93), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n303_), .A2(new_n308_), .A3(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n260_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G227gat), .A2(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(G71gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(G99gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n241_), .B(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G15gat), .B(G43gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT84), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(KEYINPUT30), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n264_), .B(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n320_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G22gat), .B(G50gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(KEYINPUT28), .B1(new_n282_), .B2(KEYINPUT29), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NOR3_X1   g127(.A1(new_n282_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n326_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n329_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n326_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n327_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G78gat), .B(G106gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT89), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n282_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n234_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n330_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n337_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G228gat), .A2(G233gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n344_), .B(KEYINPUT90), .Z(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n340_), .B1(new_n337_), .B2(new_n341_), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n343_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n337_), .A2(new_n341_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n340_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n345_), .B1(new_n351_), .B2(new_n342_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n325_), .B1(new_n348_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n346_), .B1(new_n343_), .B2(new_n347_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n325_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n351_), .A2(new_n342_), .A3(new_n345_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n353_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT33), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n308_), .A2(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n285_), .B1(new_n305_), .B2(new_n294_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n295_), .A2(new_n285_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n362_), .A2(new_n301_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n253_), .B1(new_n361_), .B2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n306_), .A2(new_n307_), .A3(KEYINPUT33), .A4(new_n301_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n360_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n250_), .A2(new_n251_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n368_));
  MUX2_X1   g167(.A(new_n257_), .B(new_n367_), .S(new_n368_), .Z(new_n369_));
  NAND2_X1  g168(.A1(new_n309_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n348_), .A2(new_n352_), .A3(new_n355_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n313_), .A2(new_n358_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G113gat), .B(G141gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT81), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G169gat), .B(G197gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G15gat), .B(G22gat), .ZN(new_n379_));
  INV_X1    g178(.A(G1gat), .ZN(new_n380_));
  INV_X1    g179(.A(G8gat), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT14), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G1gat), .B(G8gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n383_), .B(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G29gat), .B(G36gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G43gat), .B(G50gat), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n387_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n385_), .B(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(G229gat), .A3(G233gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(KEYINPUT15), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n389_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT15), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n393_), .A2(new_n396_), .A3(new_n385_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G229gat), .A2(G233gat), .ZN(new_n398_));
  XOR2_X1   g197(.A(new_n398_), .B(KEYINPUT80), .Z(new_n399_));
  OAI211_X1 g198(.A(new_n397_), .B(new_n399_), .C1(new_n390_), .C2(new_n385_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n378_), .B1(new_n392_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n392_), .A2(new_n400_), .A3(new_n378_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(KEYINPUT82), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT82), .ZN(new_n405_));
  INV_X1    g204(.A(new_n403_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n405_), .B1(new_n406_), .B2(new_n401_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n410_));
  XOR2_X1   g209(.A(KEYINPUT10), .B(G99gat), .Z(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT65), .B(G106gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT66), .ZN(new_n414_));
  INV_X1    g213(.A(G85gat), .ZN(new_n415_));
  INV_X1    g214(.A(G92gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT67), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n418_), .A3(KEYINPUT9), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G85gat), .A2(G92gat), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT9), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(KEYINPUT67), .B2(new_n421_), .ZN(new_n422_));
  OR2_X1    g221(.A1(new_n419_), .A2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G99gat), .A2(G106gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(KEYINPUT6), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT6), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n426_), .A2(G99gat), .A3(G106gat), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n419_), .A2(new_n422_), .B1(new_n425_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT66), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n411_), .A2(new_n429_), .A3(new_n412_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n414_), .A2(new_n423_), .A3(new_n428_), .A4(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(G85gat), .A2(G92gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(G85gat), .A2(G92gat), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT69), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT69), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n417_), .A2(new_n436_), .A3(new_n420_), .ZN(new_n437_));
  AOI21_X1  g236(.A(KEYINPUT8), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n425_), .A2(new_n427_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n440_));
  NOR2_X1   g239(.A1(G99gat), .A2(G106gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT7), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n439_), .A2(KEYINPUT68), .A3(new_n440_), .A4(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n438_), .A2(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n443_), .A2(new_n440_), .ZN(new_n446_));
  AOI21_X1  g245(.A(KEYINPUT68), .B1(new_n446_), .B2(new_n439_), .ZN(new_n447_));
  OAI21_X1  g246(.A(KEYINPUT70), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n439_), .A2(new_n440_), .A3(new_n443_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT68), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT70), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n451_), .A2(new_n452_), .A3(new_n444_), .A4(new_n438_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n448_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n435_), .A2(new_n437_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n449_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT8), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n432_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G57gat), .B(G64gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(KEYINPUT71), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n459_), .A2(KEYINPUT11), .ZN(new_n462_));
  XOR2_X1   g261(.A(G71gat), .B(G78gat), .Z(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n461_), .B(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n410_), .B1(new_n458_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G230gat), .A2(G233gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT64), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n468_), .B1(new_n458_), .B2(new_n465_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n464_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n461_), .B(new_n470_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n448_), .A2(new_n453_), .B1(KEYINPUT8), .B2(new_n456_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n471_), .B(KEYINPUT12), .C1(new_n472_), .C2(new_n432_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n466_), .A2(new_n469_), .A3(new_n473_), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n471_), .A2(new_n472_), .A3(new_n432_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n454_), .A2(new_n457_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n465_), .B1(new_n476_), .B2(new_n431_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n468_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(new_n478_), .ZN(new_n479_));
  XOR2_X1   g278(.A(G120gat), .B(G148gat), .Z(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT75), .ZN(new_n481_));
  XOR2_X1   g280(.A(G176gat), .B(G204gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT76), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n481_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n486_), .A2(KEYINPUT73), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n479_), .B(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n488_), .A2(KEYINPUT13), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(KEYINPUT13), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NOR3_X1   g290(.A1(new_n373_), .A2(new_n409_), .A3(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT79), .B(KEYINPUT37), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n458_), .A2(new_n394_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT78), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n393_), .A2(new_n396_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n497_), .B1(new_n472_), .B2(new_n432_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G232gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT34), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT35), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n495_), .A2(new_n496_), .A3(new_n498_), .A4(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT77), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT77), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n495_), .A2(new_n506_), .A3(new_n498_), .A4(new_n503_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n501_), .A2(new_n502_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n505_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n495_), .A2(new_n498_), .A3(new_n503_), .ZN(new_n510_));
  OAI221_X1 g309(.A(KEYINPUT77), .B1(new_n502_), .B2(new_n501_), .C1(new_n510_), .C2(KEYINPUT78), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G190gat), .B(G218gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G134gat), .B(G162gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(new_n514_), .B(KEYINPUT36), .Z(new_n515_));
  AND3_X1   g314(.A1(new_n509_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n514_), .A2(KEYINPUT36), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n518_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n494_), .B1(new_n516_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n509_), .A2(new_n511_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n517_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n509_), .A2(new_n511_), .A3(new_n515_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(new_n493_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G231gat), .A2(G233gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n385_), .B(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(new_n465_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G127gat), .B(G155gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT16), .ZN(new_n531_));
  XOR2_X1   g330(.A(G183gat), .B(G211gat), .Z(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n528_), .A2(new_n529_), .A3(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n533_), .B(KEYINPUT17), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n528_), .A2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n534_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n525_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n492_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n310_), .A2(new_n312_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n540_), .A2(G1gat), .A3(new_n541_), .ZN(new_n542_));
  XOR2_X1   g341(.A(new_n542_), .B(KEYINPUT38), .Z(new_n543_));
  NAND2_X1  g342(.A1(new_n313_), .A2(new_n358_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n371_), .A2(new_n372_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n516_), .A2(new_n519_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n491_), .A2(new_n409_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n546_), .A2(new_n548_), .A3(new_n537_), .A4(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(G1gat), .B1(new_n550_), .B2(new_n541_), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(KEYINPUT95), .Z(new_n552_));
  NAND2_X1  g351(.A1(new_n543_), .A2(new_n552_), .ZN(G1324gat));
  INV_X1    g352(.A(new_n260_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n540_), .A2(G8gat), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(G8gat), .B1(new_n550_), .B2(new_n554_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT39), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n558_), .A2(KEYINPUT96), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(KEYINPUT96), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n557_), .A2(KEYINPUT39), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT97), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n556_), .B1(new_n561_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT40), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  OAI211_X1 g366(.A(KEYINPUT40), .B(new_n556_), .C1(new_n561_), .C2(new_n564_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(G1325gat));
  OAI21_X1  g368(.A(G15gat), .B1(new_n550_), .B2(new_n325_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT41), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n540_), .A2(G15gat), .A3(new_n325_), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n571_), .A2(new_n572_), .ZN(G1326gat));
  NOR2_X1   g372(.A1(new_n348_), .A2(new_n352_), .ZN(new_n574_));
  OAI21_X1  g373(.A(G22gat), .B1(new_n550_), .B2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT42), .ZN(new_n576_));
  OR2_X1    g375(.A1(new_n574_), .A2(G22gat), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n576_), .B1(new_n540_), .B2(new_n577_), .ZN(G1327gat));
  INV_X1    g377(.A(KEYINPUT44), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT43), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n546_), .A2(new_n580_), .A3(new_n525_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT99), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT99), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n546_), .A2(new_n583_), .A3(new_n580_), .A4(new_n525_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n520_), .A2(new_n524_), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT43), .B1(new_n373_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT98), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT98), .B(KEYINPUT43), .C1(new_n373_), .C2(new_n585_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n582_), .A2(new_n584_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n549_), .A2(new_n538_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n579_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n541_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n582_), .A2(new_n584_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n588_), .A2(new_n589_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n591_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(KEYINPUT44), .A3(new_n597_), .ZN(new_n598_));
  AND4_X1   g397(.A1(G29gat), .A2(new_n592_), .A3(new_n593_), .A4(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n548_), .A2(new_n537_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n492_), .A2(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(G29gat), .B1(new_n601_), .B2(new_n593_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n599_), .A2(new_n602_), .ZN(G1328gat));
  NAND3_X1  g402(.A1(new_n592_), .A2(new_n598_), .A3(new_n260_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(G36gat), .ZN(new_n605_));
  INV_X1    g404(.A(G36gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n260_), .B(KEYINPUT100), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n601_), .A2(new_n606_), .A3(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT45), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n605_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT46), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n605_), .A2(KEYINPUT46), .A3(new_n610_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(G1329gat));
  NAND4_X1  g414(.A1(new_n592_), .A2(new_n598_), .A3(G43gat), .A4(new_n355_), .ZN(new_n616_));
  AOI21_X1  g415(.A(G43gat), .B1(new_n601_), .B2(new_n355_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT101), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g419(.A1(new_n574_), .A2(G50gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT103), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n601_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n574_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n592_), .A2(new_n598_), .A3(new_n624_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n625_), .A2(KEYINPUT102), .A3(G50gat), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT102), .B1(new_n625_), .B2(G50gat), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n623_), .B1(new_n626_), .B2(new_n627_), .ZN(G1331gat));
  INV_X1    g427(.A(new_n491_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n629_), .A2(new_n408_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR4_X1   g430(.A1(new_n373_), .A2(new_n631_), .A3(new_n547_), .A4(new_n538_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G57gat), .B1(new_n541_), .B2(KEYINPUT104), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n632_), .B(new_n633_), .C1(KEYINPUT104), .C2(G57gat), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n373_), .A2(new_n631_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(new_n539_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n636_), .A2(new_n541_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n634_), .B1(G57gat), .B2(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT105), .Z(G1332gat));
  INV_X1    g438(.A(G64gat), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n632_), .B2(new_n608_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT48), .Z(new_n642_));
  INV_X1    g441(.A(new_n636_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n643_), .A2(new_n640_), .A3(new_n608_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n642_), .A2(new_n644_), .ZN(G1333gat));
  AOI21_X1  g444(.A(new_n315_), .B1(new_n632_), .B2(new_n355_), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT49), .Z(new_n647_));
  NAND3_X1  g446(.A1(new_n643_), .A2(new_n315_), .A3(new_n355_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT106), .Z(G1334gat));
  NAND2_X1  g449(.A1(new_n632_), .A2(new_n624_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G78gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n574_), .A2(G78gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(new_n636_), .B2(new_n655_), .ZN(G1335gat));
  AND2_X1   g455(.A1(new_n635_), .A2(new_n600_), .ZN(new_n657_));
  AOI21_X1  g456(.A(G85gat), .B1(new_n657_), .B2(new_n593_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT108), .Z(new_n659_));
  NAND2_X1  g458(.A1(new_n630_), .A2(new_n538_), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT109), .B1(new_n590_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT109), .ZN(new_n662_));
  INV_X1    g461(.A(new_n660_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n596_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n661_), .A2(new_n664_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n541_), .A2(new_n415_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n659_), .B1(new_n665_), .B2(new_n666_), .ZN(G1336gat));
  NAND3_X1  g466(.A1(new_n661_), .A2(new_n664_), .A3(new_n608_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n668_), .A2(G92gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n657_), .A2(new_n416_), .A3(new_n260_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT110), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT110), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n669_), .A2(new_n673_), .A3(new_n670_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n674_), .ZN(G1337gat));
  INV_X1    g474(.A(G99gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n660_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(new_n355_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n657_), .A2(new_n411_), .A3(new_n355_), .ZN(new_n679_));
  OAI22_X1  g478(.A1(new_n678_), .A2(new_n679_), .B1(KEYINPUT111), .B2(KEYINPUT51), .ZN(new_n680_));
  NAND2_X1  g479(.A1(KEYINPUT111), .A2(KEYINPUT51), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT112), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n680_), .B(new_n682_), .ZN(G1338gat));
  NAND3_X1  g482(.A1(new_n657_), .A2(new_n412_), .A3(new_n624_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n596_), .A2(new_n624_), .A3(new_n663_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT52), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(new_n686_), .A3(G106gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n685_), .B2(G106gat), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n684_), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT53), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT53), .ZN(new_n691_));
  OAI211_X1 g490(.A(new_n691_), .B(new_n684_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(G1339gat));
  NAND3_X1  g492(.A1(new_n474_), .A2(new_n478_), .A3(new_n486_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n408_), .A2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT55), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n474_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n458_), .A2(new_n465_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n410_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n699_), .B(new_n473_), .C1(new_n477_), .C2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n468_), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n466_), .A2(new_n469_), .A3(KEYINPUT55), .A4(new_n473_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n698_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n486_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n704_), .A2(KEYINPUT56), .A3(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT56), .B1(new_n704_), .B2(new_n705_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n696_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT114), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(KEYINPUT114), .B(new_n696_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n488_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT116), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n391_), .A2(new_n399_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n385_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n399_), .B1(new_n715_), .B2(new_n394_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(new_n397_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT115), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n714_), .A2(new_n717_), .A3(new_n718_), .A4(new_n377_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n403_), .A2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n378_), .B1(new_n716_), .B2(new_n397_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n718_), .B1(new_n721_), .B2(new_n714_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n713_), .B1(new_n720_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n721_), .A2(new_n714_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT115), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n725_), .A2(KEYINPUT116), .A3(new_n403_), .A4(new_n719_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n723_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n712_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n710_), .A2(new_n711_), .A3(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n548_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT57), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT117), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT117), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n733_), .B(KEYINPUT57), .C1(new_n729_), .C2(new_n548_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n547_), .A2(new_n731_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n729_), .A2(KEYINPUT119), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT119), .B1(new_n729_), .B2(new_n736_), .ZN(new_n738_));
  AND2_X1   g537(.A1(new_n727_), .A2(new_n694_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n739_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT58), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT58), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n742_), .B(new_n739_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n585_), .B1(new_n741_), .B2(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n744_), .A2(KEYINPUT118), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT118), .ZN(new_n746_));
  AOI211_X1 g545(.A(new_n746_), .B(new_n585_), .C1(new_n741_), .C2(new_n743_), .ZN(new_n747_));
  OAI22_X1  g546(.A1(new_n737_), .A2(new_n738_), .B1(new_n745_), .B2(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(KEYINPUT120), .B1(new_n735_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n704_), .A2(new_n705_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT56), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n704_), .A2(KEYINPUT56), .A3(new_n705_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n695_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n728_), .B1(new_n754_), .B2(KEYINPUT114), .ZN(new_n755_));
  INV_X1    g554(.A(new_n711_), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n736_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT119), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n729_), .A2(KEYINPUT119), .A3(new_n736_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n752_), .A2(new_n753_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n742_), .B1(new_n761_), .B2(new_n739_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n743_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n525_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n746_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n744_), .A2(KEYINPUT118), .ZN(new_n766_));
  AOI22_X1  g565(.A1(new_n759_), .A2(new_n760_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  AOI22_X1  g566(.A1(new_n708_), .A2(new_n709_), .B1(new_n712_), .B2(new_n727_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n547_), .B1(new_n768_), .B2(new_n711_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n733_), .B1(new_n769_), .B2(KEYINPUT57), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n730_), .A2(KEYINPUT117), .A3(new_n731_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT120), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n767_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n749_), .A2(new_n538_), .A3(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n539_), .A2(new_n409_), .A3(new_n629_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777_));
  OR3_X1    g576(.A1(new_n776_), .A2(new_n777_), .A3(KEYINPUT54), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(KEYINPUT54), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n776_), .A2(KEYINPUT54), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n778_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n775_), .A2(new_n781_), .ZN(new_n782_));
  NOR3_X1   g581(.A1(new_n541_), .A2(new_n357_), .A3(new_n260_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT59), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n759_), .A2(new_n760_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n744_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n537_), .B1(new_n786_), .B2(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n781_), .B1(new_n788_), .B2(KEYINPUT121), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n788_), .A2(KEYINPUT121), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NOR4_X1   g590(.A1(new_n541_), .A2(KEYINPUT59), .A3(new_n357_), .A4(new_n260_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n785_), .A2(new_n408_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(G113gat), .ZN(new_n795_));
  OR3_X1    g594(.A1(new_n784_), .A2(G113gat), .A3(new_n409_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(G1340gat));
  NAND3_X1  g596(.A1(new_n785_), .A2(new_n491_), .A3(new_n793_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(G120gat), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT60), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n800_), .A2(G120gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(G120gat), .B1(new_n491_), .B2(new_n800_), .ZN(new_n802_));
  OR3_X1    g601(.A1(new_n784_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n799_), .A2(new_n803_), .ZN(G1341gat));
  INV_X1    g603(.A(G127gat), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n805_), .B1(new_n784_), .B2(new_n538_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT122), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  OAI211_X1 g607(.A(KEYINPUT122), .B(new_n805_), .C1(new_n784_), .C2(new_n538_), .ZN(new_n809_));
  AOI22_X1  g608(.A1(new_n784_), .A2(KEYINPUT59), .B1(new_n791_), .B2(new_n792_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n538_), .A2(new_n805_), .ZN(new_n811_));
  AOI22_X1  g610(.A1(new_n808_), .A2(new_n809_), .B1(new_n810_), .B2(new_n811_), .ZN(G1342gat));
  NAND3_X1  g611(.A1(new_n785_), .A2(new_n525_), .A3(new_n793_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(G134gat), .ZN(new_n814_));
  OR3_X1    g613(.A1(new_n784_), .A2(G134gat), .A3(new_n548_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(G1343gat));
  NOR3_X1   g615(.A1(new_n608_), .A2(new_n541_), .A3(new_n353_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n782_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n408_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n819_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n491_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g621(.A1(new_n782_), .A2(new_n817_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n823_), .A2(new_n538_), .ZN(new_n824_));
  XOR2_X1   g623(.A(KEYINPUT61), .B(G155gat), .Z(new_n825_));
  XNOR2_X1  g624(.A(new_n824_), .B(new_n825_), .ZN(G1346gat));
  OR3_X1    g625(.A1(new_n823_), .A2(G162gat), .A3(new_n548_), .ZN(new_n827_));
  OAI21_X1  g626(.A(G162gat), .B1(new_n823_), .B2(new_n585_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(G1347gat));
  NOR2_X1   g628(.A1(new_n593_), .A2(new_n607_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n355_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n409_), .ZN(new_n832_));
  XOR2_X1   g631(.A(new_n832_), .B(KEYINPUT123), .Z(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(new_n574_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n789_), .A2(new_n790_), .ZN(new_n835_));
  OAI21_X1  g634(.A(G169gat), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n836_), .A2(KEYINPUT62), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(KEYINPUT62), .ZN(new_n838_));
  NOR3_X1   g637(.A1(new_n593_), .A2(new_n607_), .A3(new_n357_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n791_), .A2(new_n839_), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n409_), .A2(new_n212_), .ZN(new_n841_));
  OAI22_X1  g640(.A1(new_n837_), .A2(new_n838_), .B1(new_n840_), .B2(new_n841_), .ZN(G1348gat));
  AND2_X1   g641(.A1(new_n791_), .A2(new_n839_), .ZN(new_n843_));
  AOI21_X1  g642(.A(G176gat), .B1(new_n843_), .B2(new_n491_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n781_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n767_), .A2(new_n772_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n537_), .B1(new_n846_), .B2(KEYINPUT120), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n845_), .B1(new_n847_), .B2(new_n774_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n624_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n831_), .A2(new_n215_), .A3(new_n629_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n844_), .B1(new_n849_), .B2(new_n850_), .ZN(G1349gat));
  NOR3_X1   g650(.A1(new_n840_), .A2(new_n218_), .A3(new_n538_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n831_), .A2(new_n538_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n782_), .A2(new_n574_), .A3(new_n853_), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n854_), .A2(KEYINPUT124), .ZN(new_n855_));
  AOI21_X1  g654(.A(G183gat), .B1(new_n854_), .B2(KEYINPUT124), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n852_), .B1(new_n855_), .B2(new_n856_), .ZN(G1350gat));
  NAND3_X1  g656(.A1(new_n843_), .A2(new_n547_), .A3(new_n219_), .ZN(new_n858_));
  OAI21_X1  g657(.A(G190gat), .B1(new_n840_), .B2(new_n585_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1351gat));
  INV_X1    g659(.A(KEYINPUT126), .ZN(new_n861_));
  OR3_X1    g660(.A1(new_n593_), .A2(KEYINPUT125), .A3(new_n353_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT125), .B1(new_n593_), .B2(new_n353_), .ZN(new_n863_));
  AND3_X1   g662(.A1(new_n862_), .A2(new_n608_), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n861_), .B1(new_n848_), .B2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n782_), .A2(KEYINPUT126), .A3(new_n864_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G197gat), .B1(new_n868_), .B2(new_n408_), .ZN(new_n869_));
  INV_X1    g668(.A(G197gat), .ZN(new_n870_));
  AOI211_X1 g669(.A(new_n870_), .B(new_n409_), .C1(new_n866_), .C2(new_n867_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n869_), .A2(new_n871_), .ZN(G1352gat));
  AOI21_X1  g671(.A(KEYINPUT126), .B1(new_n782_), .B2(new_n864_), .ZN(new_n873_));
  AOI211_X1 g672(.A(new_n861_), .B(new_n865_), .C1(new_n775_), .C2(new_n781_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n491_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(G204gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n868_), .A2(new_n226_), .A3(new_n491_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1353gat));
  NOR3_X1   g677(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n879_));
  AOI211_X1 g678(.A(new_n879_), .B(new_n538_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n881_));
  OAI21_X1  g680(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n868_), .A2(new_n882_), .A3(new_n880_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1354gat));
  INV_X1    g685(.A(G218gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n868_), .A2(new_n887_), .A3(new_n547_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n585_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n887_), .B2(new_n889_), .ZN(G1355gat));
endmodule


