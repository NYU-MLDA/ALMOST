//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_c1355" written by ABC on Sun Mar 26 01:26:03 2023

module locked_c1355 ( 
    KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5,
    KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11,
    KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17,
    KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23,
    KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29,
    KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35,
    KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41,
    KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47,
    KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53,
    KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59,
    KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat,
    G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat,
    G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat,
    G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat,
    G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat,
    G229gat, G230gat, G231gat, G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT0, KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4,
    KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10,
    KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16,
    KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22,
    KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28,
    KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34,
    KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40,
    KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46,
    KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52,
    KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58,
    KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat,
    G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat,
    G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat,
    G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat,
    G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat,
    G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n138_, new_n139_, new_n140_, new_n141_, new_n142_, new_n143_,
    new_n144_, new_n145_, new_n146_, new_n147_, new_n148_, new_n149_,
    new_n150_, new_n151_, new_n152_, new_n153_, new_n154_, new_n155_,
    new_n156_, new_n157_, new_n158_, new_n159_, new_n160_, new_n161_,
    new_n162_, new_n163_, new_n164_, new_n165_, new_n166_, new_n167_,
    new_n168_, new_n169_, new_n170_, new_n171_, new_n172_, new_n173_,
    new_n174_, new_n175_, new_n176_, new_n177_, new_n178_, new_n179_,
    new_n180_, new_n181_, new_n182_, new_n183_, new_n184_, new_n185_,
    new_n186_, new_n187_, new_n188_, new_n189_, new_n190_, new_n191_,
    new_n192_, new_n193_, new_n194_, new_n195_, new_n196_, new_n197_,
    new_n198_, new_n199_, new_n200_, new_n201_, new_n202_, new_n203_,
    new_n204_, new_n205_, new_n206_, new_n207_, new_n208_, new_n209_,
    new_n210_, new_n211_, new_n212_, new_n213_, new_n214_, new_n215_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n229_, new_n230_, new_n231_, new_n232_, new_n233_,
    new_n234_, new_n235_, new_n236_, new_n237_, new_n238_, new_n239_,
    new_n240_, new_n241_, new_n242_, new_n243_, new_n244_, new_n245_,
    new_n246_, new_n247_, new_n248_, new_n249_, new_n250_, new_n251_,
    new_n252_, new_n253_, new_n254_, new_n255_, new_n256_, new_n257_,
    new_n258_, new_n259_, new_n260_, new_n261_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n271_, new_n272_, new_n273_, new_n274_, new_n275_,
    new_n276_, new_n277_, new_n278_, new_n279_, new_n280_, new_n281_,
    new_n282_, new_n283_, new_n284_, new_n285_, new_n286_, new_n287_,
    new_n288_, new_n289_, new_n290_, new_n291_, new_n292_, new_n293_,
    new_n294_, new_n295_, new_n296_, new_n297_, new_n298_, new_n299_,
    new_n300_, new_n301_, new_n302_, new_n303_, new_n304_, new_n305_,
    new_n306_, new_n307_, new_n308_, new_n309_, new_n310_, new_n311_,
    new_n312_, new_n313_, new_n314_, new_n315_, new_n316_, new_n317_,
    new_n318_, new_n319_, new_n320_, new_n321_, new_n322_, new_n323_,
    new_n324_, new_n325_, new_n326_, new_n327_, new_n328_, new_n329_,
    new_n330_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n492_,
    new_n493_, new_n494_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n523_, new_n524_, new_n525_, new_n526_, new_n527_,
    new_n528_, new_n530_, new_n531_, new_n533_, new_n534_, new_n535_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n603_, new_n604_, new_n605_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n613_, new_n615_,
    new_n616_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n644_,
    new_n645_, new_n646_, new_n648_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n138_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n139_));
  XNOR2_X1  g002(.A(new_n138_), .B(new_n139_), .ZN(new_n140_));
  XNOR2_X1  g003(.A(G15gat), .B(G43gat), .ZN(new_n141_));
  XNOR2_X1  g004(.A(new_n140_), .B(new_n141_), .ZN(new_n142_));
  XNOR2_X1  g005(.A(G71gat), .B(G99gat), .ZN(new_n143_));
  XNOR2_X1  g006(.A(new_n142_), .B(new_n143_), .ZN(new_n144_));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n145_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n146_));
  XNOR2_X1  g009(.A(new_n145_), .B(new_n146_), .ZN(new_n147_));
  INV_X1    g010(.A(G169gat), .ZN(new_n148_));
  INV_X1    g011(.A(G176gat), .ZN(new_n149_));
  NAND2_X1  g012(.A1(new_n148_), .A2(new_n149_), .ZN(new_n150_));
  NOR2_X1   g013(.A1(new_n150_), .A2(KEYINPUT24), .ZN(new_n151_));
  NOR2_X1   g014(.A1(new_n147_), .A2(new_n151_), .ZN(new_n152_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n153_));
  NAND3_X1  g016(.A1(new_n150_), .A2(KEYINPUT24), .A3(new_n153_), .ZN(new_n154_));
  XNOR2_X1  g017(.A(KEYINPUT25), .B(G183gat), .ZN(new_n155_));
  XNOR2_X1  g018(.A(KEYINPUT26), .B(G190gat), .ZN(new_n156_));
  NAND2_X1  g019(.A1(new_n155_), .A2(new_n156_), .ZN(new_n157_));
  NAND3_X1  g020(.A1(new_n152_), .A2(new_n154_), .A3(new_n157_), .ZN(new_n158_));
  XNOR2_X1  g021(.A(KEYINPUT22), .B(G169gat), .ZN(new_n159_));
  NAND2_X1  g022(.A1(new_n159_), .A2(new_n149_), .ZN(new_n160_));
  NOR2_X1   g023(.A1(G183gat), .A2(G190gat), .ZN(new_n161_));
  OAI211_X1 g024(.A(new_n160_), .B(new_n153_), .C1(new_n147_), .C2(new_n161_), .ZN(new_n162_));
  NAND2_X1  g025(.A1(new_n158_), .A2(new_n162_), .ZN(new_n163_));
  XOR2_X1   g026(.A(new_n163_), .B(KEYINPUT30), .Z(new_n164_));
  OR2_X1    g027(.A1(new_n144_), .A2(new_n164_), .ZN(new_n165_));
  NAND2_X1  g028(.A1(G227gat), .A2(G233gat), .ZN(new_n166_));
  XOR2_X1   g029(.A(new_n166_), .B(KEYINPUT31), .Z(new_n167_));
  NAND2_X1  g030(.A1(new_n144_), .A2(new_n164_), .ZN(new_n168_));
  AND3_X1   g031(.A1(new_n165_), .A2(new_n167_), .A3(new_n168_), .ZN(new_n169_));
  AOI21_X1  g032(.A(new_n167_), .B1(new_n165_), .B2(new_n168_), .ZN(new_n170_));
  NOR2_X1   g033(.A1(new_n169_), .A2(new_n170_), .ZN(new_n171_));
  NAND2_X1  g034(.A1(G226gat), .A2(G233gat), .ZN(new_n172_));
  XOR2_X1   g035(.A(new_n172_), .B(KEYINPUT19), .Z(new_n173_));
  INV_X1    g036(.A(new_n173_), .ZN(new_n174_));
  XOR2_X1   g037(.A(G197gat), .B(G204gat), .Z(new_n175_));
  XNOR2_X1  g038(.A(G211gat), .B(G218gat), .ZN(new_n176_));
  OAI21_X1  g039(.A(new_n175_), .B1(KEYINPUT21), .B2(new_n176_), .ZN(new_n177_));
  NAND2_X1  g040(.A1(new_n176_), .A2(KEYINPUT21), .ZN(new_n178_));
  XOR2_X1   g041(.A(new_n177_), .B(new_n178_), .Z(new_n179_));
  NAND2_X1  g042(.A1(new_n179_), .A2(new_n163_), .ZN(new_n180_));
  INV_X1    g043(.A(new_n180_), .ZN(new_n181_));
  OAI21_X1  g044(.A(KEYINPUT20), .B1(new_n179_), .B2(new_n163_), .ZN(new_n182_));
  OAI21_X1  g045(.A(new_n174_), .B1(new_n181_), .B2(new_n182_), .ZN(new_n183_));
  INV_X1    g046(.A(KEYINPUT20), .ZN(new_n184_));
  INV_X1    g047(.A(new_n163_), .ZN(new_n185_));
  XNOR2_X1  g048(.A(new_n177_), .B(new_n178_), .ZN(new_n186_));
  AOI21_X1  g049(.A(new_n184_), .B1(new_n185_), .B2(new_n186_), .ZN(new_n187_));
  NAND3_X1  g050(.A1(new_n187_), .A2(new_n173_), .A3(new_n180_), .ZN(new_n188_));
  XOR2_X1   g051(.A(G8gat), .B(G36gat), .Z(new_n189_));
  XNOR2_X1  g052(.A(new_n189_), .B(KEYINPUT18), .ZN(new_n190_));
  XNOR2_X1  g053(.A(G64gat), .B(G92gat), .ZN(new_n191_));
  XNOR2_X1  g054(.A(new_n190_), .B(new_n191_), .ZN(new_n192_));
  NAND2_X1  g055(.A1(new_n192_), .A2(KEYINPUT32), .ZN(new_n193_));
  AND3_X1   g056(.A1(new_n183_), .A2(new_n188_), .A3(new_n193_), .ZN(new_n194_));
  AOI21_X1  g057(.A(new_n193_), .B1(new_n183_), .B2(new_n188_), .ZN(new_n195_));
  NOR2_X1   g058(.A1(new_n194_), .A2(new_n195_), .ZN(new_n196_));
  NOR2_X1   g059(.A1(G141gat), .A2(G148gat), .ZN(new_n197_));
  XNOR2_X1  g060(.A(new_n197_), .B(KEYINPUT3), .ZN(new_n198_));
  NAND2_X1  g061(.A1(G141gat), .A2(G148gat), .ZN(new_n199_));
  XNOR2_X1  g062(.A(new_n199_), .B(KEYINPUT2), .ZN(new_n200_));
  NAND2_X1  g063(.A1(new_n198_), .A2(new_n200_), .ZN(new_n201_));
  AND2_X1   g064(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  NOR2_X1   g065(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  NOR2_X1   g066(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g067(.A(KEYINPUT1), .ZN(new_n205_));
  AOI21_X1  g068(.A(new_n203_), .B1(new_n202_), .B2(new_n205_), .ZN(new_n206_));
  OAI21_X1  g069(.A(new_n206_), .B1(new_n205_), .B2(new_n202_), .ZN(new_n207_));
  INV_X1    g070(.A(new_n197_), .ZN(new_n208_));
  AND2_X1   g071(.A1(new_n208_), .A2(new_n199_), .ZN(new_n209_));
  AOI22_X1  g072(.A1(new_n201_), .A2(new_n204_), .B1(new_n207_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g073(.A(new_n210_), .ZN(new_n211_));
  INV_X1    g074(.A(new_n140_), .ZN(new_n212_));
  NAND3_X1  g075(.A1(new_n211_), .A2(KEYINPUT4), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n214_));
  OAI21_X1  g077(.A(new_n214_), .B1(new_n210_), .B2(new_n140_), .ZN(new_n215_));
  NAND2_X1  g078(.A1(new_n210_), .A2(new_n140_), .ZN(new_n216_));
  NAND3_X1  g079(.A1(new_n213_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  NAND2_X1  g080(.A1(G225gat), .A2(G233gat), .ZN(new_n218_));
  INV_X1    g081(.A(new_n218_), .ZN(new_n219_));
  NAND2_X1  g082(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g083(.A1(new_n211_), .A2(new_n212_), .ZN(new_n221_));
  NAND3_X1  g084(.A1(new_n221_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n222_));
  NAND2_X1  g085(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g086(.A(G1gat), .B(G29gat), .ZN(new_n224_));
  XNOR2_X1  g087(.A(new_n224_), .B(KEYINPUT0), .ZN(new_n225_));
  XNOR2_X1  g088(.A(G57gat), .B(G85gat), .ZN(new_n226_));
  XNOR2_X1  g089(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  NAND2_X1  g090(.A1(new_n223_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g091(.A(new_n227_), .ZN(new_n229_));
  NAND3_X1  g092(.A1(new_n220_), .A2(new_n222_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g093(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g094(.A1(new_n196_), .A2(new_n231_), .ZN(new_n232_));
  OR2_X1    g095(.A1(new_n211_), .A2(KEYINPUT29), .ZN(new_n233_));
  XOR2_X1   g096(.A(G78gat), .B(G106gat), .Z(new_n234_));
  XNOR2_X1  g097(.A(new_n234_), .B(KEYINPUT28), .ZN(new_n235_));
  XNOR2_X1  g098(.A(new_n233_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g099(.A(new_n236_), .ZN(new_n237_));
  INV_X1    g100(.A(G228gat), .ZN(new_n238_));
  INV_X1    g101(.A(G233gat), .ZN(new_n239_));
  NOR2_X1   g102(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  AND2_X1   g103(.A1(new_n211_), .A2(KEYINPUT29), .ZN(new_n241_));
  OAI21_X1  g104(.A(new_n240_), .B1(new_n241_), .B2(new_n186_), .ZN(new_n242_));
  AOI21_X1  g105(.A(new_n186_), .B1(new_n211_), .B2(KEYINPUT29), .ZN(new_n243_));
  INV_X1    g106(.A(new_n240_), .ZN(new_n244_));
  NAND2_X1  g107(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g108(.A(G22gat), .B(G50gat), .ZN(new_n246_));
  INV_X1    g109(.A(new_n246_), .ZN(new_n247_));
  NAND3_X1  g110(.A1(new_n242_), .A2(new_n245_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g111(.A(new_n248_), .ZN(new_n249_));
  AOI21_X1  g112(.A(new_n247_), .B1(new_n242_), .B2(new_n245_), .ZN(new_n250_));
  OAI21_X1  g113(.A(new_n237_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g114(.A1(new_n242_), .A2(new_n245_), .ZN(new_n252_));
  NAND2_X1  g115(.A1(new_n252_), .A2(new_n246_), .ZN(new_n253_));
  NAND3_X1  g116(.A1(new_n253_), .A2(new_n236_), .A3(new_n248_), .ZN(new_n254_));
  NAND2_X1  g117(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g118(.A1(new_n232_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g119(.A(new_n192_), .ZN(new_n257_));
  INV_X1    g120(.A(new_n188_), .ZN(new_n258_));
  AOI21_X1  g121(.A(new_n173_), .B1(new_n187_), .B2(new_n180_), .ZN(new_n259_));
  OAI21_X1  g122(.A(new_n257_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g123(.A1(new_n183_), .A2(new_n188_), .A3(new_n192_), .ZN(new_n261_));
  NAND2_X1  g124(.A1(new_n217_), .A2(new_n218_), .ZN(new_n262_));
  NAND3_X1  g125(.A1(new_n221_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n263_));
  NAND3_X1  g126(.A1(new_n262_), .A2(new_n227_), .A3(new_n263_), .ZN(new_n264_));
  NAND3_X1  g127(.A1(new_n260_), .A2(new_n261_), .A3(new_n264_), .ZN(new_n265_));
  INV_X1    g128(.A(KEYINPUT33), .ZN(new_n266_));
  NAND2_X1  g129(.A1(new_n230_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g130(.A(new_n267_), .ZN(new_n268_));
  NOR2_X1   g131(.A1(new_n230_), .A2(new_n266_), .ZN(new_n269_));
  NOR3_X1   g132(.A1(new_n265_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  OAI21_X1  g133(.A(new_n171_), .B1(new_n256_), .B2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g134(.A(new_n144_), .B(new_n164_), .ZN(new_n272_));
  INV_X1    g135(.A(new_n167_), .ZN(new_n273_));
  XNOR2_X1  g136(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  NAND2_X1  g137(.A1(new_n274_), .A2(new_n255_), .ZN(new_n275_));
  INV_X1    g138(.A(new_n261_), .ZN(new_n276_));
  AOI21_X1  g139(.A(new_n192_), .B1(new_n183_), .B2(new_n188_), .ZN(new_n277_));
  NOR2_X1   g140(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g141(.A1(new_n278_), .A2(KEYINPUT27), .ZN(new_n279_));
  INV_X1    g142(.A(new_n231_), .ZN(new_n280_));
  INV_X1    g143(.A(KEYINPUT27), .ZN(new_n281_));
  OAI21_X1  g144(.A(new_n281_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n282_));
  NAND3_X1  g145(.A1(new_n279_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g146(.A1(new_n171_), .A2(new_n255_), .ZN(new_n284_));
  AOI22_X1  g147(.A1(new_n271_), .A2(new_n275_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g148(.A1(G229gat), .A2(G233gat), .ZN(new_n286_));
  XNOR2_X1  g149(.A(G15gat), .B(G22gat), .ZN(new_n287_));
  INV_X1    g150(.A(G1gat), .ZN(new_n288_));
  INV_X1    g151(.A(G8gat), .ZN(new_n289_));
  OAI21_X1  g152(.A(KEYINPUT14), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g153(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g154(.A(G1gat), .B(G8gat), .Z(new_n292_));
  XNOR2_X1  g155(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g156(.A(G43gat), .B(G50gat), .ZN(new_n294_));
  XNOR2_X1  g157(.A(G29gat), .B(G36gat), .ZN(new_n295_));
  XNOR2_X1  g158(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  NAND2_X1  g159(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  XOR2_X1   g160(.A(new_n296_), .B(KEYINPUT15), .Z(new_n298_));
  OAI211_X1 g161(.A(new_n286_), .B(new_n297_), .C1(new_n298_), .C2(new_n293_), .ZN(new_n299_));
  XNOR2_X1  g162(.A(G113gat), .B(G141gat), .ZN(new_n300_));
  XNOR2_X1  g163(.A(G169gat), .B(G197gat), .ZN(new_n301_));
  XOR2_X1   g164(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  XNOR2_X1  g165(.A(new_n293_), .B(new_n296_), .ZN(new_n303_));
  NAND3_X1  g166(.A1(new_n303_), .A2(G229gat), .A3(G233gat), .ZN(new_n304_));
  NAND3_X1  g167(.A1(new_n299_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g168(.A(new_n305_), .ZN(new_n306_));
  AOI21_X1  g169(.A(new_n302_), .B1(new_n299_), .B2(new_n304_), .ZN(new_n307_));
  NOR2_X1   g170(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g171(.A(new_n308_), .ZN(new_n309_));
  NAND2_X1  g172(.A1(new_n285_), .A2(new_n309_), .ZN(new_n310_));
  XOR2_X1   g173(.A(G71gat), .B(G78gat), .Z(new_n311_));
  NAND2_X1  g174(.A1(new_n311_), .A2(KEYINPUT11), .ZN(new_n312_));
  XNOR2_X1  g175(.A(G71gat), .B(G78gat), .ZN(new_n313_));
  INV_X1    g176(.A(KEYINPUT11), .ZN(new_n314_));
  NAND2_X1  g177(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g178(.A(G57gat), .B(G64gat), .ZN(new_n316_));
  NAND3_X1  g179(.A1(new_n312_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  OR3_X1    g180(.A1(new_n313_), .A2(new_n316_), .A3(new_n314_), .ZN(new_n318_));
  NAND2_X1  g181(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  XOR2_X1   g182(.A(new_n319_), .B(new_n293_), .Z(new_n320_));
  NAND2_X1  g183(.A1(G231gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g184(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g185(.A(G127gat), .B(G155gat), .ZN(new_n323_));
  XNOR2_X1  g186(.A(new_n323_), .B(KEYINPUT16), .ZN(new_n324_));
  XOR2_X1   g187(.A(G183gat), .B(G211gat), .Z(new_n325_));
  XNOR2_X1  g188(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  INV_X1    g189(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g190(.A1(new_n322_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g191(.A(KEYINPUT17), .ZN(new_n329_));
  NAND2_X1  g192(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g193(.A1(new_n322_), .A2(KEYINPUT17), .A3(new_n327_), .ZN(new_n331_));
  OR2_X1    g194(.A1(new_n322_), .A2(new_n327_), .ZN(new_n332_));
  NAND3_X1  g195(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  INV_X1    g196(.A(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g197(.A(G134gat), .B(G162gat), .ZN(new_n335_));
  XNOR2_X1  g198(.A(G190gat), .B(G218gat), .ZN(new_n336_));
  XOR2_X1   g199(.A(new_n335_), .B(new_n336_), .Z(new_n337_));
  XNOR2_X1  g200(.A(new_n337_), .B(KEYINPUT36), .ZN(new_n338_));
  NAND2_X1  g201(.A1(G232gat), .A2(G233gat), .ZN(new_n339_));
  XOR2_X1   g202(.A(new_n339_), .B(KEYINPUT34), .Z(new_n340_));
  INV_X1    g203(.A(KEYINPUT35), .ZN(new_n341_));
  NOR2_X1   g204(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g205(.A(G85gat), .B(G92gat), .ZN(new_n343_));
  OAI21_X1  g206(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n344_));
  INV_X1    g207(.A(new_n344_), .ZN(new_n345_));
  NOR3_X1   g208(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n346_));
  NOR2_X1   g209(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g210(.A1(G99gat), .A2(G106gat), .ZN(new_n348_));
  NAND2_X1  g211(.A1(new_n348_), .A2(KEYINPUT6), .ZN(new_n349_));
  INV_X1    g212(.A(KEYINPUT6), .ZN(new_n350_));
  NAND3_X1  g213(.A1(new_n350_), .A2(G99gat), .A3(G106gat), .ZN(new_n351_));
  NAND2_X1  g214(.A1(new_n349_), .A2(new_n351_), .ZN(new_n352_));
  AOI211_X1 g215(.A(KEYINPUT8), .B(new_n343_), .C1(new_n347_), .C2(new_n352_), .ZN(new_n353_));
  INV_X1    g216(.A(KEYINPUT8), .ZN(new_n354_));
  NOR2_X1   g217(.A1(G99gat), .A2(G106gat), .ZN(new_n355_));
  INV_X1    g218(.A(KEYINPUT7), .ZN(new_n356_));
  NAND2_X1  g219(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g220(.A(new_n350_), .B1(G99gat), .B2(G106gat), .ZN(new_n358_));
  NOR2_X1   g221(.A1(new_n348_), .A2(KEYINPUT6), .ZN(new_n359_));
  OAI211_X1 g222(.A(new_n344_), .B(new_n357_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  INV_X1    g223(.A(new_n343_), .ZN(new_n361_));
  AOI21_X1  g224(.A(new_n354_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  OR2_X1    g225(.A1(new_n353_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g226(.A(KEYINPUT9), .ZN(new_n364_));
  INV_X1    g227(.A(G85gat), .ZN(new_n365_));
  INV_X1    g228(.A(G92gat), .ZN(new_n366_));
  OAI21_X1  g229(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g230(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n368_));
  OAI211_X1 g231(.A(new_n367_), .B(new_n368_), .C1(G85gat), .C2(G92gat), .ZN(new_n369_));
  XNOR2_X1  g232(.A(KEYINPUT10), .B(G99gat), .ZN(new_n370_));
  OAI211_X1 g233(.A(new_n369_), .B(new_n352_), .C1(G106gat), .C2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g234(.A(new_n298_), .B1(new_n363_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g235(.A1(new_n340_), .A2(new_n341_), .ZN(new_n373_));
  OAI21_X1  g236(.A(new_n371_), .B1(new_n353_), .B2(new_n362_), .ZN(new_n374_));
  INV_X1    g237(.A(new_n296_), .ZN(new_n375_));
  OAI21_X1  g238(.A(new_n373_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g239(.A(new_n342_), .B1(new_n372_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g240(.A(new_n377_), .ZN(new_n378_));
  NOR3_X1   g241(.A1(new_n372_), .A2(new_n376_), .A3(new_n342_), .ZN(new_n379_));
  OAI21_X1  g242(.A(new_n338_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g243(.A(new_n379_), .ZN(new_n381_));
  INV_X1    g244(.A(new_n337_), .ZN(new_n382_));
  NOR2_X1   g245(.A1(new_n382_), .A2(KEYINPUT36), .ZN(new_n383_));
  NAND3_X1  g246(.A1(new_n381_), .A2(new_n377_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g247(.A(KEYINPUT37), .ZN(new_n385_));
  NAND3_X1  g248(.A1(new_n380_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g249(.A(new_n386_), .ZN(new_n387_));
  AOI21_X1  g250(.A(new_n385_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n388_));
  NOR2_X1   g251(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NOR3_X1   g252(.A1(new_n310_), .A2(new_n334_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g253(.A1(G230gat), .A2(G233gat), .ZN(new_n391_));
  INV_X1    g254(.A(new_n319_), .ZN(new_n392_));
  NAND2_X1  g255(.A1(new_n374_), .A2(new_n392_), .ZN(new_n393_));
  OAI211_X1 g256(.A(new_n319_), .B(new_n371_), .C1(new_n362_), .C2(new_n353_), .ZN(new_n394_));
  AOI21_X1  g257(.A(new_n391_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g258(.A1(new_n393_), .A2(KEYINPUT12), .A3(new_n394_), .ZN(new_n396_));
  INV_X1    g259(.A(KEYINPUT12), .ZN(new_n397_));
  NAND3_X1  g260(.A1(new_n374_), .A2(new_n392_), .A3(new_n397_), .ZN(new_n398_));
  NAND2_X1  g261(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g262(.A(new_n395_), .B1(new_n399_), .B2(new_n391_), .ZN(new_n400_));
  XNOR2_X1  g263(.A(G176gat), .B(G204gat), .ZN(new_n401_));
  XNOR2_X1  g264(.A(new_n401_), .B(KEYINPUT5), .ZN(new_n402_));
  XNOR2_X1  g265(.A(G120gat), .B(G148gat), .ZN(new_n403_));
  XOR2_X1   g266(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  INV_X1    g267(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g268(.A1(new_n400_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g269(.A(new_n406_), .ZN(new_n407_));
  INV_X1    g270(.A(KEYINPUT13), .ZN(new_n408_));
  NOR2_X1   g271(.A1(new_n400_), .A2(new_n405_), .ZN(new_n409_));
  OR3_X1    g272(.A1(new_n407_), .A2(new_n408_), .A3(new_n409_), .ZN(new_n410_));
  OAI21_X1  g273(.A(new_n408_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n411_));
  NAND2_X1  g274(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g275(.A1(new_n412_), .A2(new_n280_), .ZN(new_n413_));
  NAND3_X1  g276(.A1(new_n390_), .A2(new_n288_), .A3(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g277(.A(new_n414_), .B(KEYINPUT38), .ZN(new_n415_));
  AND3_X1   g278(.A1(new_n381_), .A2(new_n377_), .A3(new_n383_), .ZN(new_n416_));
  INV_X1    g279(.A(new_n338_), .ZN(new_n417_));
  AOI21_X1  g280(.A(new_n417_), .B1(new_n381_), .B2(new_n377_), .ZN(new_n418_));
  NOR2_X1   g281(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g282(.A1(new_n410_), .A2(new_n333_), .A3(new_n411_), .ZN(new_n420_));
  NOR3_X1   g283(.A1(new_n310_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g284(.A(new_n421_), .ZN(new_n422_));
  OAI21_X1  g285(.A(G1gat), .B1(new_n422_), .B2(new_n280_), .ZN(new_n423_));
  NAND2_X1  g286(.A1(new_n415_), .A2(new_n423_), .ZN(G1324gat));
  NAND2_X1  g287(.A1(new_n279_), .A2(new_n282_), .ZN(new_n425_));
  INV_X1    g288(.A(new_n412_), .ZN(new_n426_));
  NAND4_X1  g289(.A1(new_n390_), .A2(new_n289_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  AND2_X1   g290(.A1(new_n285_), .A2(new_n309_), .ZN(new_n428_));
  NOR2_X1   g291(.A1(new_n420_), .A2(new_n419_), .ZN(new_n429_));
  NAND3_X1  g292(.A1(new_n428_), .A2(new_n425_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g293(.A(KEYINPUT39), .ZN(new_n431_));
  AND3_X1   g294(.A1(new_n430_), .A2(new_n431_), .A3(G8gat), .ZN(new_n432_));
  AOI21_X1  g295(.A(new_n431_), .B1(new_n430_), .B2(G8gat), .ZN(new_n433_));
  OAI21_X1  g296(.A(new_n427_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g297(.A(KEYINPUT40), .ZN(new_n435_));
  XNOR2_X1  g298(.A(new_n434_), .B(new_n435_), .ZN(G1325gat));
  NOR3_X1   g299(.A1(new_n412_), .A2(G15gat), .A3(new_n171_), .ZN(new_n437_));
  NAND2_X1  g300(.A1(new_n390_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g301(.A(G15gat), .B1(new_n422_), .B2(new_n171_), .ZN(new_n439_));
  INV_X1    g302(.A(KEYINPUT41), .ZN(new_n440_));
  AND2_X1   g303(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NOR2_X1   g304(.A1(new_n439_), .A2(new_n440_), .ZN(new_n442_));
  OAI21_X1  g305(.A(new_n438_), .B1(new_n441_), .B2(new_n442_), .ZN(G1326gat));
  NOR3_X1   g306(.A1(new_n412_), .A2(G22gat), .A3(new_n255_), .ZN(new_n444_));
  NAND2_X1  g307(.A1(new_n390_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g308(.A(G22gat), .B1(new_n422_), .B2(new_n255_), .ZN(new_n446_));
  AND2_X1   g309(.A1(new_n446_), .A2(KEYINPUT42), .ZN(new_n447_));
  NOR2_X1   g310(.A1(new_n446_), .A2(KEYINPUT42), .ZN(new_n448_));
  OAI21_X1  g311(.A(new_n445_), .B1(new_n447_), .B2(new_n448_), .ZN(G1327gat));
  NAND2_X1  g312(.A1(new_n283_), .A2(new_n284_), .ZN(new_n450_));
  AOI22_X1  g313(.A1(new_n196_), .A2(new_n231_), .B1(new_n251_), .B2(new_n254_), .ZN(new_n451_));
  INV_X1    g314(.A(new_n269_), .ZN(new_n452_));
  NAND4_X1  g315(.A1(new_n278_), .A2(new_n452_), .A3(new_n267_), .A4(new_n264_), .ZN(new_n453_));
  AOI21_X1  g316(.A(new_n274_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g317(.A(new_n255_), .ZN(new_n455_));
  NOR2_X1   g318(.A1(new_n455_), .A2(new_n171_), .ZN(new_n456_));
  OAI211_X1 g319(.A(new_n450_), .B(new_n389_), .C1(new_n454_), .C2(new_n456_), .ZN(new_n457_));
  INV_X1    g320(.A(KEYINPUT43), .ZN(new_n458_));
  NAND2_X1  g321(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g322(.A1(new_n271_), .A2(new_n275_), .ZN(new_n460_));
  NAND4_X1  g323(.A1(new_n460_), .A2(KEYINPUT43), .A3(new_n450_), .A4(new_n389_), .ZN(new_n461_));
  NOR2_X1   g324(.A1(new_n412_), .A2(new_n308_), .ZN(new_n462_));
  NAND4_X1  g325(.A1(new_n459_), .A2(new_n461_), .A3(new_n334_), .A4(new_n462_), .ZN(new_n463_));
  INV_X1    g326(.A(KEYINPUT44), .ZN(new_n464_));
  NAND2_X1  g327(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  AOI21_X1  g328(.A(new_n333_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n466_));
  NAND4_X1  g329(.A1(new_n466_), .A2(KEYINPUT44), .A3(new_n461_), .A4(new_n462_), .ZN(new_n467_));
  AND3_X1   g330(.A1(new_n465_), .A2(new_n231_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g331(.A(G29gat), .ZN(new_n469_));
  NAND4_X1  g332(.A1(new_n285_), .A2(new_n309_), .A3(new_n419_), .A4(new_n334_), .ZN(new_n470_));
  NAND2_X1  g333(.A1(new_n413_), .A2(new_n469_), .ZN(new_n471_));
  OAI22_X1  g334(.A1(new_n468_), .A2(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(G1328gat));
  NAND3_X1  g335(.A1(new_n465_), .A2(new_n425_), .A3(new_n467_), .ZN(new_n473_));
  NAND2_X1  g336(.A1(new_n473_), .A2(G36gat), .ZN(new_n474_));
  INV_X1    g337(.A(new_n425_), .ZN(new_n475_));
  OR3_X1    g338(.A1(new_n412_), .A2(new_n475_), .A3(G36gat), .ZN(new_n476_));
  OR2_X1    g339(.A1(new_n470_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g340(.A(new_n477_), .B(KEYINPUT45), .ZN(new_n478_));
  NAND2_X1  g341(.A1(new_n474_), .A2(new_n478_), .ZN(new_n479_));
  INV_X1    g342(.A(KEYINPUT46), .ZN(new_n480_));
  NAND2_X1  g343(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g344(.A1(new_n474_), .A2(new_n478_), .A3(KEYINPUT46), .ZN(new_n482_));
  NAND2_X1  g345(.A1(new_n481_), .A2(new_n482_), .ZN(G1329gat));
  NAND3_X1  g346(.A1(new_n465_), .A2(new_n274_), .A3(new_n467_), .ZN(new_n484_));
  NAND2_X1  g347(.A1(new_n484_), .A2(G43gat), .ZN(new_n485_));
  OR4_X1    g348(.A1(G43gat), .A2(new_n470_), .A3(new_n171_), .A4(new_n412_), .ZN(new_n486_));
  NAND2_X1  g349(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g350(.A(KEYINPUT47), .ZN(new_n488_));
  NAND2_X1  g351(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g352(.A1(new_n485_), .A2(new_n486_), .A3(KEYINPUT47), .ZN(new_n490_));
  NAND2_X1  g353(.A1(new_n489_), .A2(new_n490_), .ZN(G1330gat));
  AND3_X1   g354(.A1(new_n465_), .A2(new_n455_), .A3(new_n467_), .ZN(new_n492_));
  INV_X1    g355(.A(G50gat), .ZN(new_n493_));
  NAND3_X1  g356(.A1(new_n426_), .A2(new_n493_), .A3(new_n455_), .ZN(new_n494_));
  OAI22_X1  g357(.A1(new_n492_), .A2(new_n493_), .B1(new_n470_), .B2(new_n494_), .ZN(G1331gat));
  NAND2_X1  g358(.A1(new_n285_), .A2(new_n333_), .ZN(new_n496_));
  OAI21_X1  g359(.A(new_n308_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n497_));
  NOR2_X1   g360(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g361(.A(G57gat), .ZN(new_n499_));
  NOR2_X1   g362(.A1(new_n426_), .A2(new_n280_), .ZN(new_n500_));
  NAND3_X1  g363(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  NOR2_X1   g364(.A1(new_n426_), .A2(new_n309_), .ZN(new_n502_));
  INV_X1    g365(.A(new_n419_), .ZN(new_n503_));
  NAND2_X1  g366(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NOR3_X1   g367(.A1(new_n496_), .A2(new_n504_), .A3(new_n280_), .ZN(new_n505_));
  OAI21_X1  g368(.A(new_n501_), .B1(new_n505_), .B2(new_n499_), .ZN(G1332gat));
  INV_X1    g369(.A(G64gat), .ZN(new_n507_));
  NOR2_X1   g370(.A1(new_n496_), .A2(new_n504_), .ZN(new_n508_));
  AOI21_X1  g371(.A(new_n507_), .B1(new_n508_), .B2(new_n425_), .ZN(new_n509_));
  XOR2_X1   g372(.A(new_n509_), .B(KEYINPUT48), .Z(new_n510_));
  NAND4_X1  g373(.A1(new_n498_), .A2(new_n507_), .A3(new_n425_), .A4(new_n412_), .ZN(new_n511_));
  NAND2_X1  g374(.A1(new_n510_), .A2(new_n511_), .ZN(G1333gat));
  INV_X1    g375(.A(G71gat), .ZN(new_n513_));
  AOI21_X1  g376(.A(new_n513_), .B1(new_n508_), .B2(new_n274_), .ZN(new_n514_));
  XOR2_X1   g377(.A(new_n514_), .B(KEYINPUT49), .Z(new_n515_));
  NAND4_X1  g378(.A1(new_n498_), .A2(new_n513_), .A3(new_n274_), .A4(new_n412_), .ZN(new_n516_));
  NAND2_X1  g379(.A1(new_n515_), .A2(new_n516_), .ZN(G1334gat));
  INV_X1    g380(.A(G78gat), .ZN(new_n518_));
  AOI21_X1  g381(.A(new_n518_), .B1(new_n508_), .B2(new_n455_), .ZN(new_n519_));
  XOR2_X1   g382(.A(new_n519_), .B(KEYINPUT50), .Z(new_n520_));
  NAND4_X1  g383(.A1(new_n498_), .A2(new_n518_), .A3(new_n455_), .A4(new_n412_), .ZN(new_n521_));
  NAND2_X1  g384(.A1(new_n520_), .A2(new_n521_), .ZN(G1335gat));
  NOR3_X1   g385(.A1(new_n503_), .A2(new_n309_), .A3(new_n333_), .ZN(new_n523_));
  NAND2_X1  g386(.A1(new_n285_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g387(.A(new_n524_), .ZN(new_n525_));
  NAND3_X1  g388(.A1(new_n525_), .A2(new_n365_), .A3(new_n500_), .ZN(new_n526_));
  AND2_X1   g389(.A1(new_n466_), .A2(new_n461_), .ZN(new_n527_));
  AND3_X1   g390(.A1(new_n527_), .A2(new_n231_), .A3(new_n502_), .ZN(new_n528_));
  OAI21_X1  g391(.A(new_n526_), .B1(new_n528_), .B2(new_n365_), .ZN(G1336gat));
  NAND4_X1  g392(.A1(new_n525_), .A2(new_n366_), .A3(new_n425_), .A4(new_n412_), .ZN(new_n530_));
  AND3_X1   g393(.A1(new_n527_), .A2(new_n425_), .A3(new_n502_), .ZN(new_n531_));
  OAI21_X1  g394(.A(new_n530_), .B1(new_n531_), .B2(new_n366_), .ZN(G1337gat));
  NAND4_X1  g395(.A1(new_n466_), .A2(new_n274_), .A3(new_n461_), .A4(new_n502_), .ZN(new_n533_));
  NOR3_X1   g396(.A1(new_n426_), .A2(new_n171_), .A3(new_n370_), .ZN(new_n534_));
  AOI22_X1  g397(.A1(new_n533_), .A2(G99gat), .B1(new_n525_), .B2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g398(.A(new_n535_), .B(KEYINPUT51), .Z(G1338gat));
  OR4_X1    g399(.A1(G106gat), .A2(new_n524_), .A3(new_n255_), .A4(new_n426_), .ZN(new_n537_));
  NAND4_X1  g400(.A1(new_n466_), .A2(new_n455_), .A3(new_n461_), .A4(new_n502_), .ZN(new_n538_));
  INV_X1    g401(.A(KEYINPUT52), .ZN(new_n539_));
  AND3_X1   g402(.A1(new_n538_), .A2(new_n539_), .A3(G106gat), .ZN(new_n540_));
  AOI21_X1  g403(.A(new_n539_), .B1(new_n538_), .B2(G106gat), .ZN(new_n541_));
  OAI21_X1  g404(.A(new_n537_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g405(.A1(new_n542_), .A2(KEYINPUT53), .ZN(new_n543_));
  INV_X1    g406(.A(KEYINPUT53), .ZN(new_n544_));
  OAI211_X1 g407(.A(new_n544_), .B(new_n537_), .C1(new_n540_), .C2(new_n541_), .ZN(new_n545_));
  NAND2_X1  g408(.A1(new_n543_), .A2(new_n545_), .ZN(G1339gat));
  OAI21_X1  g409(.A(KEYINPUT37), .B1(new_n416_), .B2(new_n418_), .ZN(new_n547_));
  AOI21_X1  g410(.A(new_n309_), .B1(new_n547_), .B2(new_n386_), .ZN(new_n548_));
  INV_X1    g411(.A(KEYINPUT54), .ZN(new_n549_));
  NAND4_X1  g412(.A1(new_n426_), .A2(new_n548_), .A3(new_n549_), .A4(new_n333_), .ZN(new_n550_));
  OAI21_X1  g413(.A(KEYINPUT54), .B1(new_n497_), .B2(new_n420_), .ZN(new_n551_));
  NAND2_X1  g414(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g415(.A(new_n552_), .ZN(new_n553_));
  NOR2_X1   g416(.A1(new_n407_), .A2(new_n308_), .ZN(new_n554_));
  INV_X1    g417(.A(new_n391_), .ZN(new_n555_));
  NAND3_X1  g418(.A1(new_n396_), .A2(new_n555_), .A3(new_n398_), .ZN(new_n556_));
  INV_X1    g419(.A(KEYINPUT55), .ZN(new_n557_));
  AOI21_X1  g420(.A(new_n557_), .B1(new_n399_), .B2(new_n391_), .ZN(new_n558_));
  AOI211_X1 g421(.A(KEYINPUT55), .B(new_n555_), .C1(new_n396_), .C2(new_n398_), .ZN(new_n559_));
  OAI21_X1  g422(.A(new_n556_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  AND3_X1   g423(.A1(new_n560_), .A2(KEYINPUT56), .A3(new_n404_), .ZN(new_n561_));
  AOI21_X1  g424(.A(KEYINPUT56), .B1(new_n560_), .B2(new_n404_), .ZN(new_n562_));
  OAI21_X1  g425(.A(new_n554_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g426(.A(new_n302_), .B1(new_n303_), .B2(new_n286_), .ZN(new_n564_));
  OAI21_X1  g427(.A(new_n297_), .B1(new_n298_), .B2(new_n293_), .ZN(new_n565_));
  OAI21_X1  g428(.A(new_n564_), .B1(new_n565_), .B2(new_n286_), .ZN(new_n566_));
  OAI211_X1 g429(.A(new_n305_), .B(new_n566_), .C1(new_n407_), .C2(new_n409_), .ZN(new_n567_));
  NAND2_X1  g430(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g431(.A1(new_n568_), .A2(new_n503_), .ZN(new_n569_));
  INV_X1    g432(.A(KEYINPUT57), .ZN(new_n570_));
  NAND2_X1  g433(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  AND3_X1   g434(.A1(new_n406_), .A2(new_n305_), .A3(new_n566_), .ZN(new_n572_));
  OAI21_X1  g435(.A(new_n572_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n573_));
  INV_X1    g436(.A(KEYINPUT58), .ZN(new_n574_));
  NAND2_X1  g437(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  OAI211_X1 g438(.A(KEYINPUT58), .B(new_n572_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n576_));
  NAND3_X1  g439(.A1(new_n575_), .A2(new_n389_), .A3(new_n576_), .ZN(new_n577_));
  NAND3_X1  g440(.A1(new_n568_), .A2(KEYINPUT57), .A3(new_n503_), .ZN(new_n578_));
  NAND3_X1  g441(.A1(new_n571_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  AOI21_X1  g442(.A(new_n553_), .B1(new_n579_), .B2(new_n334_), .ZN(new_n580_));
  NOR2_X1   g443(.A1(new_n425_), .A2(new_n280_), .ZN(new_n581_));
  INV_X1    g444(.A(new_n581_), .ZN(new_n582_));
  NOR3_X1   g445(.A1(new_n580_), .A2(new_n275_), .A3(new_n582_), .ZN(new_n583_));
  INV_X1    g446(.A(G113gat), .ZN(new_n584_));
  NAND3_X1  g447(.A1(new_n583_), .A2(new_n584_), .A3(new_n309_), .ZN(new_n585_));
  AOI21_X1  g448(.A(KEYINPUT57), .B1(new_n568_), .B2(new_n503_), .ZN(new_n586_));
  AOI211_X1 g449(.A(new_n570_), .B(new_n419_), .C1(new_n563_), .C2(new_n567_), .ZN(new_n587_));
  NOR2_X1   g450(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  AOI21_X1  g451(.A(new_n333_), .B1(new_n588_), .B2(new_n577_), .ZN(new_n589_));
  OAI211_X1 g452(.A(new_n456_), .B(new_n581_), .C1(new_n589_), .C2(new_n553_), .ZN(new_n590_));
  INV_X1    g453(.A(KEYINPUT59), .ZN(new_n591_));
  NAND2_X1  g454(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g455(.A1(new_n579_), .A2(new_n334_), .ZN(new_n593_));
  NAND2_X1  g456(.A1(new_n593_), .A2(new_n552_), .ZN(new_n594_));
  NAND4_X1  g457(.A1(new_n594_), .A2(KEYINPUT59), .A3(new_n456_), .A4(new_n581_), .ZN(new_n595_));
  AOI21_X1  g458(.A(new_n308_), .B1(new_n592_), .B2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g459(.A(new_n585_), .B1(new_n596_), .B2(new_n584_), .ZN(G1340gat));
  INV_X1    g460(.A(G120gat), .ZN(new_n598_));
  OAI21_X1  g461(.A(new_n598_), .B1(new_n426_), .B2(KEYINPUT60), .ZN(new_n599_));
  OAI211_X1 g462(.A(new_n583_), .B(new_n599_), .C1(KEYINPUT60), .C2(new_n598_), .ZN(new_n600_));
  AOI21_X1  g463(.A(new_n426_), .B1(new_n592_), .B2(new_n595_), .ZN(new_n601_));
  OAI21_X1  g464(.A(new_n600_), .B1(new_n601_), .B2(new_n598_), .ZN(G1341gat));
  AOI21_X1  g465(.A(G127gat), .B1(new_n583_), .B2(new_n333_), .ZN(new_n603_));
  NAND2_X1  g466(.A1(new_n592_), .A2(new_n595_), .ZN(new_n604_));
  AND2_X1   g467(.A1(new_n333_), .A2(G127gat), .ZN(new_n605_));
  AOI21_X1  g468(.A(new_n603_), .B1(new_n604_), .B2(new_n605_), .ZN(G1342gat));
  AOI21_X1  g469(.A(G134gat), .B1(new_n583_), .B2(new_n419_), .ZN(new_n607_));
  AND2_X1   g470(.A1(new_n389_), .A2(G134gat), .ZN(new_n608_));
  AOI21_X1  g471(.A(new_n607_), .B1(new_n604_), .B2(new_n608_), .ZN(G1343gat));
  NOR2_X1   g472(.A1(new_n274_), .A2(new_n255_), .ZN(new_n610_));
  NAND4_X1  g473(.A1(new_n594_), .A2(new_n309_), .A3(new_n581_), .A4(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g474(.A(new_n611_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g475(.A1(new_n594_), .A2(new_n412_), .A3(new_n581_), .A4(new_n610_), .ZN(new_n613_));
  XNOR2_X1  g476(.A(new_n613_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g477(.A1(new_n594_), .A2(new_n333_), .A3(new_n581_), .A4(new_n610_), .ZN(new_n615_));
  XNOR2_X1  g478(.A(KEYINPUT61), .B(G155gat), .ZN(new_n616_));
  XNOR2_X1  g479(.A(new_n615_), .B(new_n616_), .ZN(G1346gat));
  NAND2_X1  g480(.A1(new_n594_), .A2(new_n610_), .ZN(new_n618_));
  INV_X1    g481(.A(new_n618_), .ZN(new_n619_));
  NAND3_X1  g482(.A1(new_n619_), .A2(new_n419_), .A3(new_n581_), .ZN(new_n620_));
  INV_X1    g483(.A(G162gat), .ZN(new_n621_));
  NOR2_X1   g484(.A1(new_n618_), .A2(new_n582_), .ZN(new_n622_));
  INV_X1    g485(.A(new_n389_), .ZN(new_n623_));
  NOR2_X1   g486(.A1(new_n623_), .A2(new_n621_), .ZN(new_n624_));
  AOI22_X1  g487(.A1(new_n620_), .A2(new_n621_), .B1(new_n622_), .B2(new_n624_), .ZN(G1347gat));
  NOR2_X1   g488(.A1(new_n580_), .A2(new_n275_), .ZN(new_n626_));
  NOR2_X1   g489(.A1(new_n475_), .A2(new_n231_), .ZN(new_n627_));
  NAND3_X1  g490(.A1(new_n626_), .A2(new_n309_), .A3(new_n627_), .ZN(new_n628_));
  NAND3_X1  g491(.A1(new_n628_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n629_));
  INV_X1    g492(.A(KEYINPUT62), .ZN(new_n630_));
  INV_X1    g493(.A(new_n627_), .ZN(new_n631_));
  NOR4_X1   g494(.A1(new_n580_), .A2(new_n308_), .A3(new_n275_), .A4(new_n631_), .ZN(new_n632_));
  OAI21_X1  g495(.A(new_n630_), .B1(new_n632_), .B2(new_n148_), .ZN(new_n633_));
  NAND2_X1  g496(.A1(new_n632_), .A2(new_n159_), .ZN(new_n634_));
  NAND3_X1  g497(.A1(new_n629_), .A2(new_n633_), .A3(new_n634_), .ZN(G1348gat));
  NAND3_X1  g498(.A1(new_n626_), .A2(new_n412_), .A3(new_n627_), .ZN(new_n636_));
  XNOR2_X1  g499(.A(new_n636_), .B(G176gat), .ZN(G1349gat));
  NAND3_X1  g500(.A1(new_n626_), .A2(new_n333_), .A3(new_n627_), .ZN(new_n638_));
  INV_X1    g501(.A(G183gat), .ZN(new_n639_));
  NAND2_X1  g502(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g503(.A(new_n155_), .ZN(new_n641_));
  NAND4_X1  g504(.A1(new_n626_), .A2(new_n641_), .A3(new_n333_), .A4(new_n627_), .ZN(new_n642_));
  AND2_X1   g505(.A1(new_n640_), .A2(new_n642_), .ZN(G1350gat));
  NAND2_X1  g506(.A1(new_n626_), .A2(new_n627_), .ZN(new_n644_));
  OAI21_X1  g507(.A(G190gat), .B1(new_n644_), .B2(new_n623_), .ZN(new_n645_));
  NAND2_X1  g508(.A1(new_n419_), .A2(new_n156_), .ZN(new_n646_));
  OAI21_X1  g509(.A(new_n645_), .B1(new_n644_), .B2(new_n646_), .ZN(G1351gat));
  NAND4_X1  g510(.A1(new_n594_), .A2(new_n309_), .A3(new_n610_), .A4(new_n627_), .ZN(new_n648_));
  XNOR2_X1  g511(.A(new_n648_), .B(G197gat), .ZN(G1352gat));
  NAND4_X1  g512(.A1(new_n594_), .A2(new_n412_), .A3(new_n610_), .A4(new_n627_), .ZN(new_n650_));
  XNOR2_X1  g513(.A(new_n650_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g514(.A(KEYINPUT63), .B(G211gat), .ZN(new_n652_));
  NAND4_X1  g515(.A1(new_n619_), .A2(new_n333_), .A3(new_n627_), .A4(new_n652_), .ZN(new_n653_));
  NOR3_X1   g516(.A1(new_n618_), .A2(new_n334_), .A3(new_n631_), .ZN(new_n654_));
  NOR2_X1   g517(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n655_));
  OAI21_X1  g518(.A(new_n653_), .B1(new_n654_), .B2(new_n655_), .ZN(G1354gat));
  NAND3_X1  g519(.A1(new_n619_), .A2(new_n419_), .A3(new_n627_), .ZN(new_n657_));
  INV_X1    g520(.A(G218gat), .ZN(new_n658_));
  NOR2_X1   g521(.A1(new_n618_), .A2(new_n631_), .ZN(new_n659_));
  NOR2_X1   g522(.A1(new_n623_), .A2(new_n658_), .ZN(new_n660_));
  AOI22_X1  g523(.A1(new_n657_), .A2(new_n658_), .B1(new_n659_), .B2(new_n660_), .ZN(G1355gat));
endmodule


