//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n592_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT78), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT78), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G169gat), .A3(G176gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(new_n210_), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G183gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT25), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT25), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(G183gat), .ZN(new_n217_));
  INV_X1    g016(.A(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT26), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT26), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n220_), .A2(G190gat), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n215_), .A2(new_n217_), .A3(new_n219_), .A4(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  OR3_X1    g025(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n213_), .A2(new_n222_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n231_), .B(new_n223_), .C1(G183gat), .C2(G190gat), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n210_), .A2(new_n212_), .ZN(new_n233_));
  INV_X1    g032(.A(G169gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT22), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT22), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(G169gat), .ZN(new_n237_));
  INV_X1    g036(.A(G176gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n235_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n232_), .A2(new_n233_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n228_), .A2(new_n240_), .ZN(new_n241_));
  OR2_X1    g040(.A1(G197gat), .A2(G204gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G197gat), .A2(G204gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT21), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n242_), .A2(KEYINPUT21), .A3(new_n243_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G211gat), .B(G218gat), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n247_), .A2(new_n248_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n241_), .A2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT20), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n254_));
  NAND2_X1  g053(.A1(G226gat), .A2(G233gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n254_), .B(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n253_), .A2(new_n256_), .ZN(new_n257_));
  AOI211_X1 g056(.A(new_n225_), .B(new_n224_), .C1(new_n209_), .C2(new_n208_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n258_), .A2(new_n227_), .A3(new_n222_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT87), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n235_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n210_), .A2(new_n212_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT86), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT86), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n233_), .A2(new_n264_), .A3(new_n239_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n260_), .B1(new_n266_), .B2(new_n232_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n232_), .ZN(new_n268_));
  AOI211_X1 g067(.A(KEYINPUT87), .B(new_n268_), .C1(new_n263_), .C2(new_n265_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n259_), .B1(new_n267_), .B2(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n257_), .B1(new_n270_), .B2(new_n251_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n251_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n228_), .A2(new_n249_), .A3(new_n240_), .A4(new_n250_), .ZN(new_n273_));
  AND3_X1   g072(.A1(new_n273_), .A2(KEYINPUT85), .A3(KEYINPUT20), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT85), .B1(new_n273_), .B2(KEYINPUT20), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT88), .B1(new_n277_), .B2(new_n256_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT88), .ZN(new_n279_));
  INV_X1    g078(.A(new_n256_), .ZN(new_n280_));
  AOI211_X1 g079(.A(new_n279_), .B(new_n280_), .C1(new_n272_), .C2(new_n276_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n206_), .B(new_n271_), .C1(new_n278_), .C2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT90), .ZN(new_n283_));
  INV_X1    g082(.A(new_n251_), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n261_), .A2(KEYINPUT86), .A3(new_n262_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n264_), .B1(new_n233_), .B2(new_n239_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n232_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT87), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n268_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n260_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n284_), .B1(new_n291_), .B2(new_n259_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n275_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n273_), .A2(KEYINPUT85), .A3(KEYINPUT20), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n256_), .B1(new_n292_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n279_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n277_), .A2(KEYINPUT88), .A3(new_n256_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n206_), .B1(new_n299_), .B2(new_n271_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n283_), .A2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n271_), .B1(new_n278_), .B2(new_n281_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n206_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n304_), .A2(KEYINPUT90), .A3(new_n282_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT27), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n301_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n272_), .A2(new_n280_), .A3(new_n276_), .ZN(new_n308_));
  AND3_X1   g107(.A1(new_n284_), .A2(new_n287_), .A3(new_n259_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n256_), .B1(new_n309_), .B2(new_n253_), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n282_), .B(KEYINPUT27), .C1(new_n206_), .C2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313_));
  INV_X1    g112(.A(G141gat), .ZN(new_n314_));
  INV_X1    g113(.A(G148gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT1), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT80), .ZN(new_n319_));
  INV_X1    g118(.A(G155gat), .ZN(new_n320_));
  INV_X1    g119(.A(G162gat), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT80), .B1(G155gat), .B2(G162gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n313_), .B(new_n316_), .C1(new_n318_), .C2(new_n324_), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n322_), .A2(new_n323_), .A3(new_n317_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT81), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT2), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n313_), .A2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n329_), .A2(new_n331_), .A3(new_n332_), .A4(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n326_), .A2(new_n327_), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n327_), .B1(new_n326_), .B2(new_n334_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n325_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT29), .ZN(new_n339_));
  OAI211_X1 g138(.A(KEYINPUT83), .B(new_n251_), .C1(new_n338_), .C2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G228gat), .A2(G233gat), .ZN(new_n341_));
  XOR2_X1   g140(.A(new_n341_), .B(G78gat), .Z(new_n342_));
  INV_X1    g141(.A(G106gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n340_), .B(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(G22gat), .B(G50gat), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n338_), .A2(new_n339_), .ZN(new_n349_));
  XOR2_X1   g148(.A(KEYINPUT82), .B(KEYINPUT28), .Z(new_n350_));
  OR2_X1    g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n349_), .A2(new_n350_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n348_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n351_), .A2(new_n348_), .A3(new_n352_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n346_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n355_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n345_), .B1(new_n357_), .B2(new_n353_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n356_), .A2(new_n358_), .ZN(new_n359_));
  XOR2_X1   g158(.A(KEYINPUT79), .B(G15gat), .Z(new_n360_));
  NAND2_X1  g159(.A1(G227gat), .A2(G233gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n241_), .B(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G127gat), .B(G134gat), .Z(new_n364_));
  XOR2_X1   g163(.A(G113gat), .B(G120gat), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n363_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G71gat), .B(G99gat), .ZN(new_n369_));
  INV_X1    g168(.A(G43gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT30), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT31), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n368_), .B(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT92), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n337_), .A2(new_n367_), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n366_), .B(new_n325_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n376_), .A2(KEYINPUT4), .A3(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(KEYINPUT91), .B(KEYINPUT4), .Z(new_n379_));
  NAND3_X1  g178(.A1(new_n337_), .A2(new_n367_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n375_), .B1(new_n378_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n376_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n376_), .A2(KEYINPUT4), .A3(new_n377_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n386_), .A2(KEYINPUT92), .A3(new_n382_), .A4(new_n380_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G85gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT0), .B(G57gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n393_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n384_), .A2(new_n392_), .A3(new_n385_), .A4(new_n387_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n359_), .A2(new_n374_), .A3(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n307_), .A2(new_n312_), .A3(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT97), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n396_), .ZN(new_n401_));
  AND4_X1   g200(.A1(new_n359_), .A2(new_n307_), .A3(new_n401_), .A4(new_n312_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n395_), .A2(KEYINPUT93), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT33), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n395_), .A2(KEYINPUT93), .A3(KEYINPUT33), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT94), .ZN(new_n407_));
  INV_X1    g206(.A(new_n376_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n377_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n407_), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n376_), .A2(KEYINPUT94), .A3(new_n377_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n411_), .A3(new_n382_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n380_), .A2(new_n381_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n392_), .B1(new_n413_), .B2(new_n386_), .ZN(new_n414_));
  AOI22_X1  g213(.A1(new_n405_), .A2(new_n406_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n283_), .A2(new_n300_), .ZN(new_n416_));
  AOI211_X1 g215(.A(KEYINPUT90), .B(new_n206_), .C1(new_n299_), .C2(new_n271_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT95), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT95), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n420_), .B(new_n415_), .C1(new_n416_), .C2(new_n417_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n206_), .A2(KEYINPUT32), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n423_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n299_), .A2(new_n271_), .A3(new_n422_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT96), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n424_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n426_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n419_), .A2(new_n421_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n359_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n402_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n374_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n400_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G29gat), .B(G36gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G43gat), .B(G50gat), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  XOR2_X1   g236(.A(new_n437_), .B(KEYINPUT15), .Z(new_n438_));
  XNOR2_X1  g237(.A(G15gat), .B(G22gat), .ZN(new_n439_));
  INV_X1    g238(.A(G1gat), .ZN(new_n440_));
  INV_X1    g239(.A(G8gat), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT14), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n439_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(G1gat), .B(G8gat), .ZN(new_n444_));
  XOR2_X1   g243(.A(new_n443_), .B(new_n444_), .Z(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n438_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n437_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G229gat), .A2(G233gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n447_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n445_), .B(new_n437_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n451_), .B1(new_n452_), .B2(new_n450_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G113gat), .B(G141gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G169gat), .B(G197gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n454_), .B(new_n455_), .Z(new_n456_));
  XNOR2_X1  g255(.A(new_n453_), .B(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n457_), .A2(KEYINPUT77), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(KEYINPUT77), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n434_), .A2(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G85gat), .B(G92gat), .Z(new_n462_));
  NAND2_X1  g261(.A1(G99gat), .A2(G106gat), .ZN(new_n463_));
  XOR2_X1   g262(.A(new_n463_), .B(KEYINPUT6), .Z(new_n464_));
  AND2_X1   g263(.A1(new_n464_), .A2(KEYINPUT68), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n464_), .A2(KEYINPUT68), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT69), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(G99gat), .A2(G106gat), .ZN(new_n468_));
  XOR2_X1   g267(.A(new_n468_), .B(KEYINPUT7), .Z(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n467_), .A2(new_n470_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n465_), .A2(new_n466_), .A3(KEYINPUT69), .ZN(new_n472_));
  OAI211_X1 g271(.A(KEYINPUT8), .B(new_n462_), .C1(new_n471_), .C2(new_n472_), .ZN(new_n473_));
  NOR2_X1   g272(.A1(new_n462_), .A2(KEYINPUT8), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT65), .ZN(new_n475_));
  XOR2_X1   g274(.A(KEYINPUT10), .B(G99gat), .Z(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n477_), .B2(G106gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(KEYINPUT65), .A3(new_n343_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n462_), .A2(KEYINPUT9), .ZN(new_n480_));
  XOR2_X1   g279(.A(KEYINPUT66), .B(G92gat), .Z(new_n481_));
  INV_X1    g280(.A(KEYINPUT9), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(G85gat), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n478_), .A2(new_n479_), .A3(new_n480_), .A4(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n484_), .B1(KEYINPUT8), .B2(new_n469_), .ZN(new_n485_));
  XOR2_X1   g284(.A(new_n464_), .B(KEYINPUT67), .Z(new_n486_));
  AOI21_X1  g285(.A(new_n474_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n473_), .A2(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G57gat), .B(G64gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT70), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT11), .ZN(new_n491_));
  OR2_X1    g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G71gat), .B(G78gat), .Z(new_n493_));
  OR2_X1    g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n491_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n492_), .A2(new_n495_), .A3(new_n493_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n488_), .A2(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n488_), .A2(new_n497_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n499_), .A2(KEYINPUT71), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT12), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n498_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n502_), .B1(new_n501_), .B2(new_n500_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G230gat), .A2(G233gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT64), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n498_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(new_n499_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n506_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G120gat), .B(G148gat), .Z(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT5), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G176gat), .B(G204gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n509_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n509_), .A2(new_n513_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT13), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n514_), .A2(KEYINPUT13), .A3(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT75), .ZN(new_n522_));
  XOR2_X1   g321(.A(G190gat), .B(G218gat), .Z(new_n523_));
  XNOR2_X1  g322(.A(G134gat), .B(G162gat), .ZN(new_n524_));
  OR2_X1    g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n524_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT36), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n488_), .A2(new_n438_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT73), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G232gat), .A2(G233gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n532_), .B(KEYINPUT34), .Z(new_n533_));
  INV_X1    g332(.A(KEYINPUT35), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n531_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  OAI211_X1 g334(.A(new_n530_), .B(new_n535_), .C1(new_n437_), .C2(new_n488_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n533_), .A2(new_n534_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n537_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n529_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(KEYINPUT74), .ZN(new_n542_));
  AOI21_X1  g341(.A(KEYINPUT36), .B1(new_n525_), .B2(new_n526_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n543_), .B(KEYINPUT72), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n538_), .A2(new_n539_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT74), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n545_), .B1(new_n540_), .B2(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n522_), .B1(new_n548_), .B2(KEYINPUT37), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n522_), .B(KEYINPUT37), .C1(new_n542_), .C2(new_n547_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n541_), .A2(new_n545_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n550_), .B1(KEYINPUT37), .B2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n549_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G231gat), .A2(G233gat), .ZN(new_n556_));
  XOR2_X1   g355(.A(new_n445_), .B(new_n556_), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n497_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G127gat), .B(G155gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT16), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G183gat), .B(G211gat), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n560_), .B(new_n561_), .Z(new_n562_));
  AOI21_X1  g361(.A(new_n555_), .B1(new_n558_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n558_), .A2(KEYINPUT76), .ZN(new_n564_));
  INV_X1    g363(.A(new_n562_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n564_), .B2(new_n565_), .ZN(new_n566_));
  AOI211_X1 g365(.A(new_n555_), .B(new_n562_), .C1(new_n558_), .C2(KEYINPUT76), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n554_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n461_), .A2(new_n521_), .A3(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(new_n570_), .B(KEYINPUT98), .Z(new_n571_));
  NAND3_X1  g370(.A1(new_n571_), .A2(new_n440_), .A3(new_n396_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT38), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n434_), .A2(new_n552_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n568_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n575_), .A2(new_n521_), .A3(new_n460_), .A4(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(G1gat), .B1(new_n577_), .B2(new_n401_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n572_), .A2(new_n573_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n574_), .A2(new_n578_), .A3(new_n579_), .ZN(G1324gat));
  AND2_X1   g379(.A1(new_n307_), .A2(new_n312_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n571_), .A2(new_n441_), .A3(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(G8gat), .B1(new_n577_), .B2(new_n581_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT39), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g386(.A(G15gat), .B1(new_n577_), .B2(new_n374_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT99), .B(KEYINPUT41), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n589_), .ZN(new_n591_));
  OR3_X1    g390(.A1(new_n570_), .A2(G15gat), .A3(new_n374_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .ZN(G1326gat));
  OAI21_X1  g392(.A(G22gat), .B1(new_n577_), .B2(new_n431_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT100), .B(KEYINPUT42), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n431_), .A2(G22gat), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n596_), .B1(new_n570_), .B2(new_n597_), .ZN(G1327gat));
  NAND2_X1  g397(.A1(new_n551_), .A2(new_n568_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT105), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n520_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n461_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(G29gat), .B1(new_n603_), .B2(new_n396_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT104), .ZN(new_n605_));
  INV_X1    g404(.A(new_n460_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n520_), .A2(new_n606_), .A3(new_n576_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT102), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n421_), .A2(new_n429_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n301_), .A2(new_n305_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n420_), .B1(new_n611_), .B2(new_n415_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n431_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n581_), .A2(new_n359_), .A3(new_n401_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n433_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n398_), .B(KEYINPUT97), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n609_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(KEYINPUT102), .B(new_n400_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(new_n554_), .A3(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(KEYINPUT101), .B(KEYINPUT43), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT103), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(KEYINPUT103), .A3(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n554_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n626_), .A2(KEYINPUT43), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(new_n434_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n608_), .B1(new_n625_), .B2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n605_), .B1(new_n629_), .B2(KEYINPUT44), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n619_), .A2(KEYINPUT103), .A3(new_n620_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT103), .B1(new_n619_), .B2(new_n620_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n607_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT44), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(KEYINPUT104), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n630_), .A2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n633_), .A2(KEYINPUT44), .A3(new_n607_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n396_), .A2(G29gat), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n604_), .B1(new_n639_), .B2(new_n640_), .ZN(G1328gat));
  INV_X1    g440(.A(G36gat), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n603_), .A2(new_n642_), .A3(new_n582_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT45), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n638_), .A2(new_n582_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n645_), .B1(new_n630_), .B2(new_n636_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT106), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n646_), .A2(new_n647_), .A3(new_n642_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n581_), .B1(new_n629_), .B2(KEYINPUT44), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT104), .B1(new_n634_), .B2(new_n635_), .ZN(new_n650_));
  AOI211_X1 g449(.A(new_n605_), .B(KEYINPUT44), .C1(new_n633_), .C2(new_n607_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n649_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT106), .B1(new_n652_), .B2(G36gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n644_), .B1(new_n648_), .B2(new_n653_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  OAI211_X1 g456(.A(new_n644_), .B(new_n655_), .C1(new_n648_), .C2(new_n653_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1329gat));
  NAND4_X1  g458(.A1(new_n637_), .A2(G43gat), .A3(new_n433_), .A4(new_n638_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n370_), .B1(new_n602_), .B2(new_n374_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g462(.A1(new_n639_), .A2(new_n359_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G50gat), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n431_), .A2(G50gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT108), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n665_), .B1(new_n602_), .B2(new_n667_), .ZN(G1331gat));
  NAND4_X1  g467(.A1(new_n575_), .A2(new_n606_), .A3(new_n520_), .A4(new_n576_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT110), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G57gat), .B1(new_n671_), .B2(new_n401_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n434_), .A2(new_n606_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(new_n520_), .A3(new_n569_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT109), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n401_), .A2(G57gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n672_), .B1(new_n676_), .B2(new_n677_), .ZN(G1332gat));
  INV_X1    g477(.A(G64gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n679_), .B1(new_n670_), .B2(new_n582_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT48), .Z(new_n681_));
  NAND3_X1  g480(.A1(new_n675_), .A2(new_n679_), .A3(new_n582_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(G1333gat));
  OAI21_X1  g482(.A(G71gat), .B1(new_n671_), .B2(new_n374_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n374_), .A2(G71gat), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT112), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n686_), .B1(new_n676_), .B2(new_n688_), .ZN(G1334gat));
  OAI21_X1  g488(.A(G78gat), .B1(new_n671_), .B2(new_n431_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT50), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n431_), .A2(G78gat), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n691_), .B1(new_n676_), .B2(new_n692_), .ZN(G1335gat));
  NOR2_X1   g492(.A1(new_n521_), .A2(new_n600_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n673_), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n695_), .A2(G85gat), .A3(new_n401_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n520_), .A2(new_n606_), .A3(new_n568_), .ZN(new_n697_));
  AOI22_X1  g496(.A1(new_n623_), .A2(new_n624_), .B1(new_n434_), .B2(new_n627_), .ZN(new_n698_));
  OR2_X1    g497(.A1(new_n698_), .A2(KEYINPUT113), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(KEYINPUT113), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n697_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(new_n396_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n696_), .B1(new_n702_), .B2(G85gat), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT114), .Z(G1336gat));
  INV_X1    g503(.A(new_n695_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G92gat), .B1(new_n705_), .B2(new_n582_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n582_), .A2(new_n481_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n706_), .B1(new_n701_), .B2(new_n707_), .ZN(G1337gat));
  NOR3_X1   g507(.A1(new_n695_), .A2(new_n374_), .A3(new_n477_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n701_), .A2(new_n433_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(G99gat), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT51), .Z(G1338gat));
  OR2_X1    g511(.A1(new_n697_), .A2(new_n431_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G106gat), .B1(new_n698_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT52), .ZN(new_n715_));
  OR2_X1    g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n715_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n695_), .A2(G106gat), .A3(new_n431_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT115), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n716_), .A2(new_n717_), .A3(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g520(.A(KEYINPUT55), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n506_), .A2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n503_), .A2(KEYINPUT55), .A3(new_n505_), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n723_), .B(new_n724_), .C1(new_n505_), .C2(new_n503_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n513_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT56), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n725_), .A2(KEYINPUT56), .A3(new_n513_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n514_), .A2(new_n460_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n456_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n453_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n452_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n456_), .B1(new_n734_), .B2(new_n450_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n735_), .A2(KEYINPUT116), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n450_), .B1(new_n445_), .B2(new_n448_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n447_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n735_), .A2(KEYINPUT116), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n733_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  AOI22_X1  g539(.A1(new_n730_), .A2(new_n731_), .B1(new_n516_), .B2(new_n740_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n741_), .A2(new_n551_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT57), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(KEYINPUT117), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n514_), .A2(new_n740_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT58), .B1(new_n730_), .B2(new_n746_), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n747_), .A2(new_n626_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n730_), .A2(KEYINPUT58), .A3(new_n746_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT117), .B(new_n743_), .C1(new_n741_), .C2(new_n551_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n745_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n521_), .A2(new_n569_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT54), .B1(new_n753_), .B2(new_n460_), .ZN(new_n754_));
  OR3_X1    g553(.A1(new_n753_), .A2(KEYINPUT54), .A3(new_n460_), .ZN(new_n755_));
  AOI22_X1  g554(.A1(new_n752_), .A2(new_n568_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n582_), .A2(new_n401_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n757_), .A2(new_n433_), .A3(new_n431_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(G113gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(new_n460_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n756_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n758_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(KEYINPUT59), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT59), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n765_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n606_), .B1(new_n764_), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n761_), .B1(new_n767_), .B2(new_n760_), .ZN(G1340gat));
  INV_X1    g567(.A(G120gat), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n769_), .B1(new_n521_), .B2(KEYINPUT60), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n759_), .B(new_n770_), .C1(KEYINPUT60), .C2(new_n769_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n521_), .B1(new_n764_), .B2(new_n766_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(new_n769_), .ZN(G1341gat));
  AOI21_X1  g572(.A(new_n568_), .B1(new_n764_), .B2(new_n766_), .ZN(new_n774_));
  INV_X1    g573(.A(G127gat), .ZN(new_n775_));
  INV_X1    g574(.A(new_n759_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n576_), .A2(new_n775_), .ZN(new_n777_));
  OAI22_X1  g576(.A1(new_n774_), .A2(new_n775_), .B1(new_n776_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(KEYINPUT118), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780_));
  OAI221_X1 g579(.A(new_n780_), .B1(new_n776_), .B2(new_n777_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n779_), .A2(new_n781_), .ZN(G1342gat));
  INV_X1    g581(.A(G134gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n776_), .B2(new_n552_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n784_), .A2(KEYINPUT119), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(KEYINPUT119), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n764_), .A2(new_n766_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n626_), .A2(new_n783_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n785_), .A2(new_n786_), .B1(new_n787_), .B2(new_n788_), .ZN(G1343gat));
  NOR2_X1   g588(.A1(new_n431_), .A2(new_n433_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n757_), .A2(new_n790_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT120), .Z(new_n792_));
  NAND2_X1  g591(.A1(new_n762_), .A2(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n793_), .A2(new_n606_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(new_n794_), .B(new_n314_), .ZN(G1344gat));
  NOR2_X1   g594(.A1(new_n793_), .A2(new_n521_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(new_n315_), .ZN(G1345gat));
  NOR2_X1   g596(.A1(new_n793_), .A2(new_n568_), .ZN(new_n798_));
  XOR2_X1   g597(.A(KEYINPUT61), .B(G155gat), .Z(new_n799_));
  XNOR2_X1  g598(.A(new_n798_), .B(new_n799_), .ZN(G1346gat));
  OAI21_X1  g599(.A(G162gat), .B1(new_n793_), .B2(new_n626_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n551_), .A2(new_n321_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n793_), .B2(new_n802_), .ZN(G1347gat));
  AND2_X1   g602(.A1(new_n582_), .A2(new_n397_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n762_), .A2(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(G169gat), .B1(new_n805_), .B2(new_n606_), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n806_), .A2(KEYINPUT62), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(KEYINPUT62), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n460_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT121), .ZN(new_n810_));
  OAI22_X1  g609(.A1(new_n807_), .A2(new_n808_), .B1(new_n805_), .B2(new_n810_), .ZN(G1348gat));
  NOR2_X1   g610(.A1(new_n805_), .A2(new_n521_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(new_n238_), .ZN(G1349gat));
  NAND2_X1  g612(.A1(new_n215_), .A2(new_n217_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n762_), .A2(new_n814_), .A3(new_n576_), .A4(new_n804_), .ZN(new_n815_));
  OR2_X1    g614(.A1(new_n815_), .A2(KEYINPUT122), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n214_), .B1(new_n805_), .B2(new_n568_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n818_), .B1(KEYINPUT122), .B2(new_n815_), .ZN(G1350gat));
  OAI21_X1  g618(.A(G190gat), .B1(new_n805_), .B2(new_n626_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n551_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n820_), .B1(new_n805_), .B2(new_n821_), .ZN(G1351gat));
  INV_X1    g621(.A(KEYINPUT123), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n582_), .A2(new_n401_), .A3(new_n790_), .ZN(new_n824_));
  OR3_X1    g623(.A1(new_n756_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n823_), .B1(new_n756_), .B2(new_n824_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n460_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n521_), .B1(new_n830_), .B2(G204gat), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n827_), .A2(new_n831_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n830_), .A2(G204gat), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n832_), .B(new_n833_), .Z(G1353gat));
  AOI21_X1  g633(.A(new_n568_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n835_));
  XOR2_X1   g634(.A(new_n835_), .B(KEYINPUT125), .Z(new_n836_));
  NOR2_X1   g635(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n836_), .B1(KEYINPUT126), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n827_), .A2(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n837_), .A2(KEYINPUT126), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1354gat));
  INV_X1    g640(.A(G218gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n827_), .A2(new_n842_), .A3(new_n551_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n626_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n844_), .B2(new_n842_), .ZN(G1355gat));
endmodule


