//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n820_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n867_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n881_, new_n882_;
  AOI21_X1  g000(.A(G176gat), .B1(KEYINPUT83), .B2(KEYINPUT22), .ZN(new_n202_));
  INV_X1    g001(.A(G169gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G183gat), .A2(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT23), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n207_), .B1(new_n208_), .B2(new_n206_), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n209_), .B1(G183gat), .B2(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT84), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n204_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n212_), .B1(new_n211_), .B2(new_n210_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G169gat), .A2(G176gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n214_), .B(KEYINPUT80), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216_));
  INV_X1    g015(.A(G176gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n203_), .A2(new_n217_), .ZN(new_n218_));
  NOR3_X1   g017(.A1(new_n215_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT25), .B(G183gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT82), .B1(new_n205_), .B2(KEYINPUT23), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n208_), .A2(new_n205_), .ZN(new_n224_));
  MUX2_X1   g023(.A(KEYINPUT82), .B(new_n223_), .S(new_n224_), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n215_), .A2(new_n216_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n222_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n213_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT30), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT85), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G71gat), .B(G99gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(G43gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G227gat), .A2(G233gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(G15gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n234_), .B(new_n236_), .ZN(new_n237_));
  OR2_X1    g036(.A1(new_n232_), .A2(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n230_), .A2(new_n231_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n232_), .A2(new_n237_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G113gat), .B(G120gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n242_), .B(new_n243_), .Z(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT31), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n241_), .A2(KEYINPUT86), .A3(new_n246_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n241_), .A2(KEYINPUT86), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n245_), .B1(new_n241_), .B2(KEYINPUT86), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G197gat), .B(G204gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT21), .ZN(new_n252_));
  OR2_X1    g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G211gat), .B(G218gat), .Z(new_n254_));
  AND2_X1   g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n251_), .A2(new_n252_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n254_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n228_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n225_), .B1(G183gat), .B2(G190gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT22), .B(G169gat), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n218_), .B1(new_n261_), .B2(new_n217_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n226_), .A2(new_n209_), .A3(KEYINPUT94), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n226_), .A2(new_n209_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT94), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n222_), .A2(new_n264_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n263_), .A2(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n259_), .B(KEYINPUT20), .C1(new_n258_), .C2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G226gat), .A2(G233gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT19), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT20), .B1(new_n228_), .B2(new_n258_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT95), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n269_), .A2(new_n276_), .A3(new_n258_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n276_), .B1(new_n269_), .B2(new_n258_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n275_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n273_), .B1(new_n280_), .B2(new_n272_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(G8gat), .B(G36gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT18), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G64gat), .B(G92gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n283_), .B(new_n284_), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n285_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n272_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n269_), .A2(new_n258_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT95), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n277_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n288_), .B1(new_n291_), .B2(new_n275_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n287_), .B1(new_n292_), .B2(new_n273_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n286_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT27), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n295_), .B1(new_n281_), .B2(new_n285_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n288_), .B(new_n275_), .C1(new_n278_), .C2(new_n279_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n270_), .A2(new_n272_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n287_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n296_), .A2(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G78gat), .B(G106gat), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT89), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G141gat), .A2(G148gat), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT2), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT3), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n308_), .A2(new_n309_), .B1(new_n310_), .B2(KEYINPUT88), .ZN(new_n311_));
  NOR2_X1   g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n312_), .B1(KEYINPUT88), .B2(new_n310_), .ZN(new_n313_));
  OR3_X1    g112(.A1(new_n312_), .A2(KEYINPUT88), .A3(new_n310_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n307_), .A2(new_n311_), .A3(new_n313_), .A4(new_n314_), .ZN(new_n315_));
  AND2_X1   g114(.A1(G155gat), .A2(G162gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G155gat), .A2(G162gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT90), .B1(new_n315_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n318_), .A2(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n312_), .A2(KEYINPUT87), .ZN(new_n322_));
  AOI21_X1  g121(.A(new_n312_), .B1(KEYINPUT87), .B2(new_n308_), .ZN(new_n323_));
  AOI211_X1 g122(.A(new_n322_), .B(new_n323_), .C1(KEYINPUT1), .C2(new_n316_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n319_), .B1(new_n321_), .B2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n315_), .A2(KEYINPUT90), .A3(new_n318_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT29), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT92), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n258_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n328_), .A2(KEYINPUT92), .ZN(new_n331_));
  OAI211_X1 g130(.A(G228gat), .B(G233gat), .C1(new_n330_), .C2(new_n331_), .ZN(new_n332_));
  OR2_X1    g131(.A1(new_n328_), .A2(KEYINPUT91), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n328_), .A2(KEYINPUT91), .ZN(new_n334_));
  INV_X1    g133(.A(new_n258_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n335_), .B1(G228gat), .B2(G233gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n333_), .A2(new_n334_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n305_), .B1(new_n332_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n332_), .A2(new_n337_), .A3(new_n305_), .ZN(new_n340_));
  OR3_X1    g139(.A1(new_n327_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n341_));
  OAI21_X1  g140(.A(KEYINPUT28), .B1(new_n327_), .B2(KEYINPUT29), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G22gat), .B(G50gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n343_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n345_), .A2(KEYINPUT93), .A3(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT93), .B1(new_n345_), .B2(new_n346_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n339_), .B(new_n340_), .C1(new_n347_), .C2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n340_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n348_), .B1(new_n351_), .B2(new_n338_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n244_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n325_), .A2(new_n354_), .A3(new_n326_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(G225gat), .A2(G233gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n355_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n360_), .B(KEYINPUT96), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n363_), .B(new_n364_), .C1(new_n358_), .C2(new_n362_), .ZN(new_n365_));
  XOR2_X1   g164(.A(G1gat), .B(G29gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G57gat), .B(G85gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n368_), .B(new_n369_), .Z(new_n370_));
  NAND3_X1  g169(.A1(new_n361_), .A2(new_n365_), .A3(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(KEYINPUT98), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT98), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n361_), .A2(new_n365_), .A3(new_n373_), .A4(new_n370_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n361_), .A2(new_n365_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n370_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n372_), .A2(new_n374_), .A3(new_n377_), .ZN(new_n378_));
  NOR4_X1   g177(.A1(new_n250_), .A2(new_n303_), .A3(new_n353_), .A4(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT99), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n285_), .A2(KEYINPUT32), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n381_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n382_), .B1(new_n281_), .B2(new_n381_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n378_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT33), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n360_), .B(new_n363_), .C1(new_n358_), .C2(new_n362_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n370_), .B1(new_n359_), .B2(new_n364_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n371_), .A2(new_n385_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n361_), .A2(new_n365_), .A3(KEYINPUT33), .A4(new_n370_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n388_), .A2(new_n286_), .A3(new_n293_), .A4(new_n389_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n384_), .A2(new_n350_), .A3(new_n390_), .A4(new_n352_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n250_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n294_), .A2(new_n295_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n378_), .ZN(new_n394_));
  AOI22_X1  g193(.A1(new_n393_), .A2(new_n394_), .B1(new_n350_), .B2(new_n352_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n380_), .B1(new_n392_), .B2(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n353_), .B1(new_n303_), .B2(new_n378_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n397_), .A2(KEYINPUT99), .A3(new_n391_), .A4(new_n250_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n379_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT69), .ZN(new_n400_));
  AND2_X1   g199(.A1(G85gat), .A2(G92gat), .ZN(new_n401_));
  NOR2_X1   g200(.A1(G85gat), .A2(G92gat), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n401_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(G99gat), .A2(G106gat), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT68), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT7), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT7), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(KEYINPUT68), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n405_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  AOI211_X1 g209(.A(G99gat), .B(G106gat), .C1(new_n406_), .C2(KEYINPUT7), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(G99gat), .A2(G106gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(KEYINPUT6), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT6), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(G99gat), .A3(G106gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n404_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT8), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n400_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n407_), .A2(new_n405_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT68), .B(KEYINPUT7), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n417_), .B(new_n421_), .C1(new_n405_), .C2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n403_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n414_), .A2(new_n416_), .A3(KEYINPUT66), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT66), .B1(new_n414_), .B2(new_n416_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n412_), .A3(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n430_), .A2(new_n419_), .A3(new_n403_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n420_), .A2(new_n425_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT67), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n426_), .A2(new_n428_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n435_), .B1(new_n402_), .B2(KEYINPUT65), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT65), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n437_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n438_));
  INV_X1    g237(.A(G92gat), .ZN(new_n439_));
  OR2_X1    g238(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n440_));
  NAND2_X1  g239(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  OAI211_X1 g241(.A(new_n436_), .B(new_n438_), .C1(new_n442_), .C2(KEYINPUT9), .ZN(new_n443_));
  AND2_X1   g242(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n444_));
  NOR2_X1   g243(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n444_), .A2(new_n445_), .A3(G106gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  AND4_X1   g246(.A1(new_n433_), .A2(new_n434_), .A3(new_n443_), .A4(new_n447_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n426_), .A2(new_n428_), .A3(new_n446_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n433_), .B1(new_n449_), .B2(new_n443_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G29gat), .B(G36gat), .Z(new_n452_));
  XOR2_X1   g251(.A(G43gat), .B(G50gat), .Z(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n432_), .A2(new_n451_), .A3(new_n454_), .ZN(new_n455_));
  OR2_X1    g254(.A1(new_n455_), .A2(KEYINPUT73), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(KEYINPUT73), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n432_), .A2(new_n451_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n454_), .B(KEYINPUT15), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT35), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G232gat), .A2(G233gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT34), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  AOI22_X1  g262(.A1(new_n458_), .A2(new_n459_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n456_), .A2(new_n457_), .A3(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n463_), .A2(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n466_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n456_), .A2(new_n468_), .A3(new_n457_), .A4(new_n464_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G190gat), .B(G218gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G134gat), .B(G162gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n471_), .B(new_n472_), .ZN(new_n473_));
  NOR3_X1   g272(.A1(new_n470_), .A2(KEYINPUT36), .A3(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n473_), .B(KEYINPUT36), .Z(new_n475_));
  AND2_X1   g274(.A1(new_n470_), .A2(new_n475_), .ZN(new_n476_));
  OAI22_X1  g275(.A1(new_n474_), .A2(new_n476_), .B1(KEYINPUT74), .B2(KEYINPUT37), .ZN(new_n477_));
  NAND2_X1  g276(.A1(KEYINPUT74), .A2(KEYINPUT37), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n478_), .B(KEYINPUT75), .Z(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G127gat), .B(G155gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT16), .ZN(new_n483_));
  XOR2_X1   g282(.A(G183gat), .B(G211gat), .Z(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT78), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n486_), .B(KEYINPUT17), .Z(new_n487_));
  XNOR2_X1  g286(.A(G15gat), .B(G22gat), .ZN(new_n488_));
  INV_X1    g287(.A(G1gat), .ZN(new_n489_));
  INV_X1    g288(.A(G8gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT14), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G1gat), .B(G8gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G231gat), .A2(G233gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G57gat), .B(G64gat), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n497_), .A2(KEYINPUT11), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(KEYINPUT11), .ZN(new_n499_));
  XOR2_X1   g298(.A(G71gat), .B(G78gat), .Z(new_n500_));
  NAND3_X1  g299(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n499_), .A2(new_n500_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n496_), .B(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT77), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n504_), .A2(KEYINPUT77), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n487_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(KEYINPUT76), .B(KEYINPUT17), .ZN(new_n508_));
  OR3_X1    g307(.A1(new_n504_), .A2(new_n485_), .A3(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n507_), .A2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  OAI221_X1 g310(.A(new_n479_), .B1(KEYINPUT74), .B2(KEYINPUT37), .C1(new_n474_), .C2(new_n476_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n481_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT79), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G230gat), .A2(G233gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n503_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n458_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n432_), .A2(new_n451_), .A3(new_n503_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n516_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n520_), .A2(KEYINPUT70), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n518_), .A2(new_n519_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n516_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(KEYINPUT70), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n521_), .A2(new_n524_), .ZN(new_n525_));
  AND3_X1   g324(.A1(new_n432_), .A2(new_n503_), .A3(new_n451_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n503_), .B1(new_n432_), .B2(new_n451_), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT12), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT12), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n518_), .A2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n516_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n525_), .A2(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G120gat), .B(G148gat), .Z(new_n534_));
  XNOR2_X1  g333(.A(G176gat), .B(G204gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n538_), .A2(KEYINPUT71), .ZN(new_n539_));
  INV_X1    g338(.A(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n533_), .A2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n539_), .B1(new_n525_), .B2(new_n532_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT13), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(KEYINPUT13), .A3(new_n542_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n459_), .A2(new_n494_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n454_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n549_), .A2(new_n494_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G229gat), .A2(G233gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n549_), .B(new_n494_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n554_), .A2(G229gat), .A3(G233gat), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G113gat), .B(G141gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G169gat), .B(G197gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  OR2_X1    g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n556_), .A2(new_n559_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n547_), .A2(new_n562_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n399_), .A2(new_n515_), .A3(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(new_n489_), .A3(new_n378_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n565_), .B(KEYINPUT38), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n474_), .A2(new_n476_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n567_), .A2(KEYINPUT101), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(KEYINPUT101), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OR3_X1    g369(.A1(new_n563_), .A2(KEYINPUT100), .A3(new_n510_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT100), .B1(new_n563_), .B2(new_n510_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n396_), .A2(new_n398_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n379_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(new_n378_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(G1gat), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n579_), .A2(KEYINPUT102), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(KEYINPUT102), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n566_), .B1(new_n580_), .B2(new_n581_), .ZN(G1324gat));
  NAND3_X1  g381(.A1(new_n564_), .A2(new_n490_), .A3(new_n303_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT39), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n577_), .A2(new_n303_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n584_), .B1(new_n585_), .B2(G8gat), .ZN(new_n586_));
  AOI211_X1 g385(.A(KEYINPUT39), .B(new_n490_), .C1(new_n577_), .C2(new_n303_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n583_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT40), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(G1325gat));
  INV_X1    g389(.A(G15gat), .ZN(new_n591_));
  INV_X1    g390(.A(new_n250_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n564_), .A2(new_n591_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n577_), .A2(new_n592_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n594_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n595_));
  AOI21_X1  g394(.A(KEYINPUT41), .B1(new_n594_), .B2(G15gat), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n593_), .B1(new_n595_), .B2(new_n596_), .ZN(G1326gat));
  INV_X1    g396(.A(G22gat), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n564_), .A2(new_n598_), .A3(new_n353_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n577_), .A2(new_n353_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(G22gat), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n601_), .A2(KEYINPUT42), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(KEYINPUT42), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n599_), .B1(new_n602_), .B2(new_n603_), .ZN(G1327gat));
  NOR2_X1   g403(.A1(new_n567_), .A2(new_n511_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT103), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n399_), .A2(new_n563_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(G29gat), .B1(new_n607_), .B2(new_n378_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n563_), .A2(new_n511_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT43), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n481_), .A2(new_n512_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n610_), .B1(new_n576_), .B2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n611_), .ZN(new_n613_));
  NOR3_X1   g412(.A1(new_n399_), .A2(KEYINPUT43), .A3(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n609_), .B1(new_n612_), .B2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT44), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(KEYINPUT44), .B(new_n609_), .C1(new_n612_), .C2(new_n614_), .ZN(new_n618_));
  AND2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n378_), .A2(G29gat), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n608_), .B1(new_n619_), .B2(new_n620_), .ZN(G1328gat));
  INV_X1    g420(.A(KEYINPUT46), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(KEYINPUT104), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n617_), .A2(new_n303_), .A3(new_n618_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G36gat), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n622_), .A2(KEYINPUT104), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT45), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n393_), .A2(G36gat), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n607_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n628_), .B1(new_n607_), .B2(new_n629_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n627_), .B1(new_n630_), .B2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n624_), .B1(new_n626_), .B2(new_n633_), .ZN(new_n634_));
  AOI211_X1 g433(.A(new_n623_), .B(new_n632_), .C1(new_n625_), .C2(G36gat), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(G1329gat));
  NAND4_X1  g435(.A1(new_n617_), .A2(G43gat), .A3(new_n592_), .A4(new_n618_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n607_), .A2(new_n592_), .ZN(new_n638_));
  OR2_X1    g437(.A1(new_n638_), .A2(G43gat), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g440(.A(G50gat), .B1(new_n607_), .B2(new_n353_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n353_), .A2(G50gat), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n642_), .B1(new_n619_), .B2(new_n643_), .ZN(G1331gat));
  INV_X1    g443(.A(KEYINPUT105), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n515_), .B2(new_n547_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n399_), .A2(new_n562_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n545_), .A2(new_n546_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n514_), .A2(KEYINPUT105), .A3(new_n648_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n646_), .A2(new_n647_), .A3(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(G57gat), .B1(new_n651_), .B2(new_n378_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n547_), .A2(new_n562_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  NOR4_X1   g453(.A1(new_n399_), .A2(new_n510_), .A3(new_n570_), .A4(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n394_), .A2(KEYINPUT106), .ZN(new_n656_));
  MUX2_X1   g455(.A(KEYINPUT106), .B(new_n656_), .S(G57gat), .Z(new_n657_));
  AOI21_X1  g456(.A(new_n652_), .B1(new_n655_), .B2(new_n657_), .ZN(G1332gat));
  INV_X1    g457(.A(G64gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n659_), .B1(new_n655_), .B2(new_n303_), .ZN(new_n660_));
  XOR2_X1   g459(.A(new_n660_), .B(KEYINPUT48), .Z(new_n661_));
  NAND2_X1  g460(.A1(new_n303_), .A2(new_n659_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT107), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n661_), .B1(new_n650_), .B2(new_n663_), .ZN(G1333gat));
  INV_X1    g463(.A(G71gat), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n665_), .B1(new_n655_), .B2(new_n592_), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT49), .Z(new_n667_));
  NAND2_X1  g466(.A1(new_n592_), .A2(new_n665_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n667_), .B1(new_n650_), .B2(new_n668_), .ZN(G1334gat));
  INV_X1    g468(.A(G78gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n655_), .B2(new_n353_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT50), .Z(new_n672_));
  NAND3_X1  g471(.A1(new_n651_), .A2(new_n670_), .A3(new_n353_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(G1335gat));
  NOR2_X1   g473(.A1(new_n612_), .A2(new_n614_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n654_), .A2(new_n511_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n440_), .A2(new_n441_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n378_), .A3(new_n679_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n399_), .A2(new_n606_), .A3(new_n654_), .ZN(new_n681_));
  AOI21_X1  g480(.A(G85gat), .B1(new_n681_), .B2(new_n378_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n683_), .A2(KEYINPUT108), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(KEYINPUT108), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n680_), .A2(new_n684_), .A3(new_n685_), .ZN(G1336gat));
  NAND3_X1  g485(.A1(new_n678_), .A2(G92gat), .A3(new_n303_), .ZN(new_n687_));
  AOI21_X1  g486(.A(G92gat), .B1(new_n681_), .B2(new_n303_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n687_), .B1(KEYINPUT109), .B2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(KEYINPUT109), .B2(new_n688_), .ZN(G1337gat));
  NOR2_X1   g489(.A1(new_n444_), .A2(new_n445_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n681_), .A2(new_n592_), .A3(new_n691_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT110), .Z(new_n693_));
  INV_X1    g492(.A(G99gat), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n675_), .A2(new_n250_), .A3(new_n677_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT51), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT51), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n693_), .B(new_n698_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1338gat));
  INV_X1    g499(.A(G106gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n681_), .A2(new_n701_), .A3(new_n353_), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n353_), .B(new_n676_), .C1(new_n612_), .C2(new_n614_), .ZN(new_n703_));
  XNOR2_X1  g502(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n703_), .A2(G106gat), .A3(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n703_), .B2(G106gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n702_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g507(.A(KEYINPUT55), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n531_), .A2(new_n709_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n528_), .A2(KEYINPUT55), .A3(new_n530_), .A4(new_n516_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n529_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n527_), .A2(KEYINPUT12), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n523_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n710_), .A2(new_n711_), .A3(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT112), .ZN(new_n716_));
  INV_X1    g515(.A(new_n538_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT112), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n710_), .A2(new_n718_), .A3(new_n711_), .A4(new_n714_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n716_), .A2(KEYINPUT56), .A3(new_n717_), .A4(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT113), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n719_), .A2(new_n717_), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n723_), .A2(KEYINPUT113), .A3(KEYINPUT56), .A4(new_n716_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT56), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n719_), .A2(new_n717_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n516_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n709_), .B2(new_n531_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n718_), .B1(new_n728_), .B2(new_n711_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n726_), .B2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n722_), .A2(new_n724_), .A3(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n559_), .B1(new_n554_), .B2(new_n552_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n551_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n552_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n561_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n533_), .B2(new_n538_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n731_), .A2(KEYINPUT58), .A3(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n611_), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT58), .B1(new_n731_), .B2(new_n736_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n533_), .A2(new_n538_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n562_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n730_), .B2(new_n720_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n735_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n567_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT57), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  OAI211_X1 g546(.A(KEYINPUT57), .B(new_n567_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n510_), .B1(new_n740_), .B2(new_n749_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n562_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n545_), .A2(new_n751_), .A3(new_n546_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n513_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT54), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n513_), .A2(new_n752_), .A3(KEYINPUT54), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n750_), .A2(new_n758_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n250_), .A2(new_n353_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n303_), .A2(new_n394_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n759_), .A2(new_n763_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n764_), .A2(KEYINPUT114), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(KEYINPUT114), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n765_), .A2(new_n562_), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(G113gat), .ZN(new_n768_));
  OAI211_X1 g567(.A(new_n747_), .B(new_n748_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n769_), .A2(KEYINPUT116), .A3(new_n510_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT116), .B1(new_n769_), .B2(new_n510_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n758_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  XOR2_X1   g571(.A(KEYINPUT115), .B(KEYINPUT59), .Z(new_n773_));
  NOR2_X1   g572(.A1(new_n762_), .A2(new_n773_), .ZN(new_n774_));
  AOI22_X1  g573(.A1(new_n772_), .A2(new_n774_), .B1(new_n764_), .B2(KEYINPUT59), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n562_), .A2(G113gat), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT117), .Z(new_n777_));
  AOI22_X1  g576(.A1(new_n767_), .A2(new_n768_), .B1(new_n775_), .B2(new_n777_), .ZN(G1340gat));
  AOI21_X1  g577(.A(new_n757_), .B1(new_n510_), .B2(new_n769_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT59), .B1(new_n779_), .B2(new_n762_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n750_), .A2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n769_), .A2(KEYINPUT116), .A3(new_n510_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n757_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n774_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n648_), .B(new_n780_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT118), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT60), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n547_), .B2(G120gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n765_), .A2(new_n766_), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n772_), .A2(new_n774_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n648_), .A4(new_n780_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n787_), .A2(new_n790_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(G120gat), .ZN(new_n795_));
  OR2_X1    g594(.A1(new_n790_), .A2(KEYINPUT60), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(G1341gat));
  NAND3_X1  g596(.A1(new_n765_), .A2(new_n511_), .A3(new_n766_), .ZN(new_n798_));
  INV_X1    g597(.A(G127gat), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n511_), .A2(G127gat), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT119), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n798_), .A2(new_n799_), .B1(new_n775_), .B2(new_n801_), .ZN(G1342gat));
  NAND2_X1  g601(.A1(new_n775_), .A2(new_n611_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(G134gat), .ZN(new_n804_));
  INV_X1    g603(.A(new_n570_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(G134gat), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n765_), .A2(new_n766_), .A3(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(KEYINPUT120), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT120), .ZN(new_n809_));
  INV_X1    g608(.A(new_n807_), .ZN(new_n810_));
  INV_X1    g609(.A(G134gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n775_), .B2(new_n611_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n809_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n808_), .A2(new_n813_), .ZN(G1343gat));
  INV_X1    g613(.A(new_n353_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n779_), .A2(new_n815_), .A3(new_n592_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n761_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(new_n751_), .ZN(new_n818_));
  XOR2_X1   g617(.A(new_n818_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g618(.A1(new_n817_), .A2(new_n547_), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(G148gat), .Z(G1345gat));
  XNOR2_X1  g620(.A(KEYINPUT61), .B(G155gat), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT121), .B1(new_n817_), .B2(new_n510_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n817_), .A2(KEYINPUT121), .A3(new_n510_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n823_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n826_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(new_n824_), .A3(new_n822_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(G1346gat));
  INV_X1    g629(.A(G162gat), .ZN(new_n831_));
  NOR3_X1   g630(.A1(new_n817_), .A2(new_n831_), .A3(new_n613_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n817_), .A2(new_n805_), .ZN(new_n833_));
  OR3_X1    g632(.A1(new_n833_), .A2(KEYINPUT122), .A3(G162gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(KEYINPUT122), .B1(new_n833_), .B2(G162gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n832_), .B1(new_n834_), .B2(new_n835_), .ZN(G1347gat));
  NOR2_X1   g635(.A1(new_n393_), .A2(new_n378_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n760_), .A2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n784_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(new_n261_), .A3(new_n562_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT62), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n250_), .A2(new_n378_), .A3(new_n393_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  OR3_X1    g642(.A1(new_n843_), .A2(KEYINPUT123), .A3(new_n751_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT123), .B1(new_n843_), .B2(new_n751_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n353_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n772_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n841_), .B1(new_n847_), .B2(G169gat), .ZN(new_n848_));
  AOI211_X1 g647(.A(KEYINPUT62), .B(new_n203_), .C1(new_n772_), .C2(new_n846_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n840_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT124), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT124), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n852_), .B(new_n840_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(G1348gat));
  NOR2_X1   g653(.A1(new_n779_), .A2(new_n353_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n843_), .A2(new_n217_), .A3(new_n547_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NOR3_X1   g656(.A1(new_n784_), .A2(new_n547_), .A3(new_n838_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(G176gat), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT125), .ZN(G1349gat));
  NOR2_X1   g659(.A1(new_n843_), .A2(new_n510_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G183gat), .B1(new_n855_), .B2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n510_), .A2(new_n220_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n839_), .B2(new_n863_), .ZN(G1350gat));
  NAND3_X1  g663(.A1(new_n839_), .A2(new_n221_), .A3(new_n570_), .ZN(new_n865_));
  INV_X1    g664(.A(G190gat), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n784_), .A2(new_n613_), .A3(new_n838_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n865_), .B1(new_n866_), .B2(new_n867_), .ZN(G1351gat));
  NAND2_X1  g667(.A1(new_n816_), .A2(new_n837_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n562_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g671(.A1(new_n869_), .A2(new_n547_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT126), .B(G204gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1353gat));
  AOI21_X1  g674(.A(new_n510_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n876_));
  XOR2_X1   g675(.A(new_n876_), .B(KEYINPUT127), .Z(new_n877_));
  NAND2_X1  g676(.A1(new_n870_), .A2(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n879_));
  XOR2_X1   g678(.A(new_n878_), .B(new_n879_), .Z(G1354gat));
  OR3_X1    g679(.A1(new_n869_), .A2(G218gat), .A3(new_n805_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G218gat), .B1(new_n869_), .B2(new_n613_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1355gat));
endmodule


