//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n736_, new_n737_, new_n738_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n920_, new_n921_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  INV_X1    g002(.A(G36gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(G29gat), .ZN(new_n205_));
  INV_X1    g004(.A(G29gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(G36gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT74), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n203_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n206_), .A2(G36gat), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n204_), .A2(G29gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT74), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(new_n202_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT15), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n211_), .A2(new_n216_), .A3(KEYINPUT15), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G99gat), .A2(G106gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT6), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT6), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(G99gat), .A3(G106gat), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT7), .ZN(new_n228_));
  INV_X1    g027(.A(G99gat), .ZN(new_n229_));
  INV_X1    g028(.A(G106gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n222_), .B1(new_n227_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n224_), .A2(new_n226_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n235_), .A2(KEYINPUT67), .A3(new_n232_), .A4(new_n231_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT68), .B(KEYINPUT8), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  INV_X1    g037(.A(G85gat), .ZN(new_n239_));
  INV_X1    g038(.A(G92gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n237_), .A2(new_n238_), .A3(new_n241_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n234_), .A2(new_n236_), .A3(new_n242_), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n241_), .A2(new_n238_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n244_), .B1(new_n227_), .B2(new_n233_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT8), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n241_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT9), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n238_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n238_), .A2(KEYINPUT66), .A3(new_n250_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n249_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT10), .B(G99gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(KEYINPUT65), .B(G106gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n235_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n255_), .A2(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n221_), .B1(new_n247_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT75), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G232gat), .A2(G233gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(KEYINPUT34), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n263_), .B2(KEYINPUT35), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n259_), .B1(new_n243_), .B2(new_n246_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n217_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n260_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n263_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT35), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n260_), .B(new_n267_), .C1(new_n270_), .C2(new_n269_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G190gat), .B(G218gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G134gat), .B(G162gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XOR2_X1   g076(.A(new_n277_), .B(KEYINPUT36), .Z(new_n278_));
  NAND2_X1  g077(.A1(new_n274_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n277_), .A2(KEYINPUT36), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n272_), .A2(new_n273_), .A3(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n274_), .A2(KEYINPUT76), .A3(new_n278_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n281_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT37), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(KEYINPUT77), .ZN(new_n287_));
  INV_X1    g086(.A(new_n279_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n283_), .ZN(new_n289_));
  OR3_X1    g088(.A1(new_n288_), .A2(KEYINPUT37), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT77), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n284_), .A2(new_n283_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT76), .B1(new_n274_), .B2(new_n278_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n291_), .B(KEYINPUT37), .C1(new_n292_), .C2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n287_), .A2(new_n290_), .A3(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G57gat), .B(G64gat), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n296_), .A2(KEYINPUT11), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(KEYINPUT11), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G71gat), .B(G78gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n297_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(new_n298_), .B2(new_n300_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G15gat), .B(G22gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G1gat), .A2(G8gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT14), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G1gat), .ZN(new_n307_));
  INV_X1    g106(.A(G8gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(new_n304_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n306_), .A2(new_n310_), .ZN(new_n311_));
  NAND4_X1  g110(.A1(new_n303_), .A2(new_n304_), .A3(new_n309_), .A4(new_n305_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n302_), .B(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G231gat), .A2(G233gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(G127gat), .B(G155gat), .Z(new_n317_));
  XNOR2_X1  g116(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G183gat), .B(G211gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT17), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n316_), .A2(new_n322_), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n321_), .A2(KEYINPUT17), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n316_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n295_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT79), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G113gat), .B(G141gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(G169gat), .B(G197gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n330_), .B(new_n331_), .Z(new_n332_));
  INV_X1    g131(.A(KEYINPUT81), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n211_), .A2(new_n216_), .A3(new_n311_), .A4(new_n312_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n334_), .B2(KEYINPUT80), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(KEYINPUT80), .A3(new_n333_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n336_), .A2(new_n313_), .A3(new_n217_), .A4(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n217_), .A2(new_n313_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n337_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(new_n335_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n338_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G229gat), .A2(G233gat), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n221_), .A2(new_n313_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n346_), .A2(new_n343_), .A3(new_n334_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n332_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n343_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n347_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n332_), .ZN(new_n351_));
  NOR3_X1   g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G57gat), .B(G85gat), .Z(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT97), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(new_n307_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(new_n206_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n357_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G141gat), .A2(G148gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT85), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT2), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n367_), .B1(new_n365_), .B2(new_n362_), .ZN(new_n368_));
  NOR3_X1   g167(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(G155gat), .A2(G162gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G155gat), .A2(G162gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT87), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n372_), .A2(KEYINPUT87), .A3(new_n373_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n371_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT88), .ZN(new_n379_));
  NOR2_X1   g178(.A1(G155gat), .A2(G162gat), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n373_), .B1(new_n380_), .B2(KEYINPUT1), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT86), .ZN(new_n382_));
  OR2_X1    g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n373_), .A2(KEYINPUT1), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n364_), .B1(G141gat), .B2(G148gat), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n378_), .B(new_n379_), .C1(new_n386_), .C2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n387_), .B1(new_n383_), .B2(new_n385_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n376_), .A2(new_n377_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n390_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT88), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G127gat), .B(G134gat), .Z(new_n393_));
  XOR2_X1   g192(.A(G113gat), .B(G120gat), .Z(new_n394_));
  XOR2_X1   g193(.A(new_n393_), .B(new_n394_), .Z(new_n395_));
  NAND3_X1  g194(.A1(new_n388_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n389_), .A2(new_n391_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n395_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n396_), .A2(KEYINPUT4), .A3(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT4), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n388_), .A2(new_n392_), .A3(new_n403_), .A4(new_n395_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n400_), .A2(KEYINPUT95), .A3(new_n402_), .A4(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n396_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n404_), .A2(new_n402_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(KEYINPUT95), .B1(new_n409_), .B2(new_n400_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n361_), .B1(new_n407_), .B2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT98), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT95), .ZN(new_n413_));
  INV_X1    g212(.A(new_n400_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n413_), .B1(new_n414_), .B2(new_n408_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n415_), .A2(new_n360_), .A3(new_n406_), .A4(new_n405_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n411_), .A2(new_n412_), .A3(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(KEYINPUT89), .B(G204gat), .Z(new_n418_));
  NAND3_X1  g217(.A1(new_n418_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n419_));
  INV_X1    g218(.A(G197gat), .ZN(new_n420_));
  AOI21_X1  g219(.A(KEYINPUT90), .B1(new_n420_), .B2(G204gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT89), .B(G204gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n421_), .B1(new_n422_), .B2(new_n420_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n419_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G211gat), .B(G218gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n422_), .A2(G197gat), .ZN(new_n429_));
  INV_X1    g228(.A(G204gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(KEYINPUT21), .B1(new_n420_), .B2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n428_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n419_), .A2(KEYINPUT92), .A3(new_n423_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n428_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n433_), .A2(KEYINPUT21), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT92), .B1(new_n419_), .B2(new_n423_), .ZN(new_n436_));
  OAI22_X1  g235(.A1(new_n427_), .A2(new_n432_), .B1(new_n435_), .B2(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(G169gat), .A2(G176gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT82), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(G169gat), .A2(G176gat), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n440_), .A2(KEYINPUT24), .A3(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT25), .B(G183gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT26), .B(G190gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G183gat), .A2(G190gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n446_), .B(KEYINPUT23), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT24), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n438_), .A2(new_n448_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n442_), .A2(new_n445_), .A3(new_n447_), .A4(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(G183gat), .ZN(new_n451_));
  INV_X1    g250(.A(G190gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n447_), .A2(new_n453_), .ZN(new_n454_));
  XOR2_X1   g253(.A(new_n441_), .B(KEYINPUT83), .Z(new_n455_));
  XOR2_X1   g254(.A(KEYINPUT22), .B(G169gat), .Z(new_n456_));
  OAI211_X1 g255(.A(new_n454_), .B(new_n455_), .C1(G176gat), .C2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n450_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n437_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n436_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n460_), .A2(KEYINPUT21), .A3(new_n434_), .A4(new_n433_), .ZN(new_n461_));
  INV_X1    g260(.A(G176gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT84), .ZN(new_n463_));
  INV_X1    g262(.A(G169gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT22), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  OR2_X1    g264(.A1(new_n464_), .A2(KEYINPUT22), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n462_), .B(new_n465_), .C1(new_n466_), .C2(new_n463_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n454_), .A2(new_n455_), .A3(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n446_), .B(KEYINPUT23), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n445_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n470_), .B1(new_n448_), .B2(new_n439_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n440_), .A2(KEYINPUT24), .A3(new_n455_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n468_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n426_), .B(new_n428_), .C1(new_n429_), .C2(new_n431_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n461_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n459_), .A2(KEYINPUT20), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G226gat), .A2(G233gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT19), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n471_), .A2(new_n472_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n468_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n437_), .A2(new_n482_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n461_), .A2(new_n474_), .A3(new_n450_), .A4(new_n457_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n478_), .ZN(new_n485_));
  NAND4_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(KEYINPUT20), .A4(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n479_), .A2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G8gat), .B(G36gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT18), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G64gat), .B(G92gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  AND2_X1   g290(.A1(new_n491_), .A2(KEYINPUT32), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n487_), .A2(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT20), .B1(new_n437_), .B2(new_n458_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n473_), .B1(new_n474_), .B2(new_n461_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n478_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n459_), .A2(new_n475_), .A3(KEYINPUT20), .A4(new_n485_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n493_), .B1(new_n498_), .B2(new_n492_), .ZN(new_n499_));
  OAI211_X1 g298(.A(KEYINPUT98), .B(new_n361_), .C1(new_n407_), .C2(new_n410_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n417_), .A2(new_n499_), .A3(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n407_), .A2(new_n410_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(KEYINPUT33), .A3(new_n360_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n491_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n487_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n479_), .A2(new_n491_), .A3(new_n486_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n400_), .A2(new_n401_), .A3(new_n404_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n396_), .A2(new_n399_), .A3(new_n402_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n361_), .A3(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n505_), .A2(new_n506_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT33), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n416_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n503_), .A2(new_n510_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n501_), .A2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n388_), .A2(new_n392_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT29), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n517_), .A2(KEYINPUT28), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT28), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n515_), .A2(new_n519_), .A3(new_n516_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G22gat), .B(G50gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n518_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n521_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n519_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n524_));
  AOI211_X1 g323(.A(KEYINPUT28), .B(KEYINPUT29), .C1(new_n388_), .C2(new_n392_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n522_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G228gat), .A2(G233gat), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n437_), .B(new_n528_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n437_), .B1(new_n516_), .B2(new_n397_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n528_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n529_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G78gat), .B(G106gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT93), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n535_), .A2(KEYINPUT93), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n529_), .A2(new_n532_), .A3(new_n536_), .A4(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n527_), .A2(new_n538_), .A3(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n535_), .A2(KEYINPUT94), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n533_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n529_), .B(new_n532_), .C1(KEYINPUT94), .C2(new_n535_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n543_), .A2(new_n522_), .A3(new_n526_), .A4(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G71gat), .B(G99gat), .ZN(new_n547_));
  INV_X1    g346(.A(G43gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n482_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n549_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n473_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n395_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G227gat), .A2(G233gat), .ZN(new_n555_));
  INV_X1    g354(.A(G15gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n555_), .B(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT30), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT31), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n550_), .A2(new_n398_), .A3(new_n552_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n554_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n559_), .B1(new_n554_), .B2(new_n560_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n546_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n514_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n417_), .A2(new_n500_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT27), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT99), .ZN(new_n568_));
  AOI22_X1  g367(.A1(new_n506_), .A2(new_n568_), .B1(new_n498_), .B2(new_n504_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n479_), .A2(KEYINPUT99), .A3(new_n491_), .A4(new_n486_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n567_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  AND3_X1   g370(.A1(new_n505_), .A2(new_n567_), .A3(new_n506_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n563_), .B1(new_n541_), .B2(new_n545_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n541_), .A2(new_n545_), .A3(new_n563_), .ZN(new_n574_));
  OAI221_X1 g373(.A(new_n566_), .B1(new_n571_), .B2(new_n572_), .C1(new_n573_), .C2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n354_), .B1(new_n565_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT69), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n577_), .B1(new_n265_), .B2(new_n302_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(KEYINPUT12), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G230gat), .A2(G233gat), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT64), .Z(new_n581_));
  NAND2_X1  g380(.A1(new_n265_), .A2(new_n302_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT12), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n577_), .B(new_n583_), .C1(new_n265_), .C2(new_n302_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n579_), .A2(new_n581_), .A3(new_n582_), .A4(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n581_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n582_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n265_), .A2(new_n302_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n586_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n585_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G176gat), .B(G204gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT71), .ZN(new_n592_));
  XNOR2_X1  g391(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n592_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G120gat), .B(G148gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n590_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n596_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n585_), .A2(new_n589_), .A3(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n597_), .B1(KEYINPUT72), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(KEYINPUT72), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n598_), .B1(new_n585_), .B2(new_n589_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n604_));
  NOR2_X1   g403(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NOR3_X1   g405(.A1(new_n600_), .A2(new_n603_), .A3(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n600_), .A2(new_n603_), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n608_), .B1(new_n609_), .B2(new_n604_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n329_), .A2(new_n576_), .A3(new_n610_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n611_), .A2(G1gat), .A3(new_n566_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(KEYINPUT38), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT101), .ZN(new_n614_));
  OR3_X1    g413(.A1(new_n288_), .A2(KEYINPUT100), .A3(new_n289_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT100), .B1(new_n288_), .B2(new_n289_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n617_), .B1(new_n565_), .B2(new_n575_), .ZN(new_n618_));
  AND4_X1   g417(.A1(new_n353_), .A2(new_n618_), .A3(new_n610_), .A4(new_n327_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n566_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n307_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n621_), .B1(new_n612_), .B2(KEYINPUT38), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n614_), .A2(new_n622_), .ZN(G1324gat));
  NOR2_X1   g422(.A1(new_n571_), .A2(new_n572_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n619_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(G8gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT39), .ZN(new_n627_));
  INV_X1    g426(.A(new_n611_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n308_), .A3(new_n624_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n627_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n630_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1325gat));
  AOI21_X1  g433(.A(new_n556_), .B1(new_n619_), .B2(new_n563_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT41), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n628_), .A2(new_n556_), .A3(new_n563_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1326gat));
  NAND2_X1  g437(.A1(new_n619_), .A2(new_n546_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(G22gat), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT42), .ZN(new_n641_));
  INV_X1    g440(.A(new_n546_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n642_), .A2(G22gat), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n641_), .B1(new_n611_), .B2(new_n643_), .ZN(G1327gat));
  NOR2_X1   g443(.A1(new_n609_), .A2(new_n604_), .ZN(new_n645_));
  OAI211_X1 g444(.A(new_n353_), .B(new_n326_), .C1(new_n645_), .C2(new_n607_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT103), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n647_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n294_), .A2(new_n290_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n291_), .B1(new_n285_), .B2(KEYINPUT37), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI22_X1  g452(.A1(new_n574_), .A2(new_n573_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(new_n620_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n563_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n642_), .A2(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n501_), .B2(new_n513_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n653_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n653_), .B2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n659_), .A2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT43), .B1(new_n295_), .B2(KEYINPUT104), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n565_), .A2(new_n575_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n664_), .B1(new_n665_), .B2(new_n653_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n650_), .B1(new_n663_), .B2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT44), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n659_), .A2(new_n662_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n665_), .A2(new_n664_), .A3(new_n653_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(KEYINPUT44), .A3(new_n650_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n669_), .A2(new_n673_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n566_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n645_), .A2(new_n607_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n617_), .A2(new_n326_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n576_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n620_), .A2(new_n206_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n675_), .B1(new_n679_), .B2(new_n680_), .ZN(G1328gat));
  INV_X1    g480(.A(new_n624_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(G36gat), .ZN(new_n683_));
  INV_X1    g482(.A(new_n683_), .ZN(new_n684_));
  OR3_X1    g483(.A1(new_n679_), .A2(KEYINPUT106), .A3(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT106), .B1(new_n679_), .B2(new_n684_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(KEYINPUT45), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT45), .B1(new_n685_), .B2(new_n686_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AOI221_X4 g488(.A(new_n668_), .B1(new_n648_), .B2(new_n649_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n690_));
  AOI21_X1  g489(.A(KEYINPUT44), .B1(new_n672_), .B2(new_n650_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT105), .B1(new_n692_), .B2(new_n624_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n669_), .A2(KEYINPUT105), .A3(new_n624_), .A4(new_n673_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(G36gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n689_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n689_), .B(KEYINPUT46), .C1(new_n693_), .C2(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1329gat));
  NOR3_X1   g499(.A1(new_n679_), .A2(G43gat), .A3(new_n656_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n674_), .A2(new_n656_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(new_n548_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT47), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(KEYINPUT47), .B(new_n702_), .C1(new_n703_), .C2(new_n548_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1330gat));
  OAI21_X1  g507(.A(G50gat), .B1(new_n674_), .B2(new_n642_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n642_), .A2(G50gat), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT107), .Z(new_n711_));
  OAI21_X1  g510(.A(new_n709_), .B1(new_n679_), .B2(new_n711_), .ZN(G1331gat));
  NOR2_X1   g511(.A1(new_n353_), .A2(new_n326_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n676_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n618_), .A2(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G57gat), .B1(new_n715_), .B2(new_n566_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n665_), .A2(KEYINPUT108), .A3(new_n354_), .ZN(new_n717_));
  AOI21_X1  g516(.A(KEYINPUT108), .B1(new_n665_), .B2(new_n354_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n329_), .A2(new_n676_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n566_), .A2(G57gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n716_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT109), .Z(G1332gat));
  INV_X1    g523(.A(G64gat), .ZN(new_n725_));
  INV_X1    g524(.A(new_n715_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n725_), .B1(new_n726_), .B2(new_n624_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728_));
  OR2_X1    g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n728_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n729_), .A2(KEYINPUT48), .A3(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n624_), .A2(new_n725_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n731_), .B1(new_n721_), .B2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT48), .B1(new_n729_), .B2(new_n730_), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n733_), .A2(new_n734_), .ZN(G1333gat));
  OAI21_X1  g534(.A(G71gat), .B1(new_n715_), .B2(new_n656_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT49), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n656_), .A2(G71gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n721_), .B2(new_n738_), .ZN(G1334gat));
  OAI21_X1  g538(.A(G78gat), .B1(new_n715_), .B2(new_n642_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT50), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n642_), .A2(G78gat), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n741_), .B1(new_n721_), .B2(new_n742_), .ZN(G1335gat));
  NAND3_X1  g542(.A1(new_n676_), .A2(new_n354_), .A3(new_n326_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT111), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n672_), .A2(new_n745_), .A3(KEYINPUT112), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(KEYINPUT112), .B1(new_n672_), .B2(new_n745_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(G85gat), .B1(new_n749_), .B2(new_n566_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n610_), .A2(new_n677_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n719_), .A2(new_n239_), .A3(new_n620_), .A4(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT113), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT113), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n750_), .A2(new_n755_), .A3(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1336gat));
  OAI21_X1  g556(.A(G92gat), .B1(new_n749_), .B2(new_n682_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n719_), .A2(new_n751_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n624_), .A2(new_n240_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n759_), .B2(new_n760_), .ZN(G1337gat));
  NAND2_X1  g560(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n762_));
  OR2_X1    g561(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n672_), .A2(new_n745_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT112), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n746_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n229_), .B1(new_n767_), .B2(new_n563_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n656_), .A2(new_n256_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n751_), .B(new_n769_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT114), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  OAI211_X1 g571(.A(new_n762_), .B(new_n763_), .C1(new_n768_), .C2(new_n772_), .ZN(new_n773_));
  OAI21_X1  g572(.A(G99gat), .B1(new_n749_), .B2(new_n656_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n774_), .A2(KEYINPUT115), .A3(KEYINPUT51), .A4(new_n771_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1338gat));
  OR3_X1    g575(.A1(new_n759_), .A2(new_n642_), .A3(new_n257_), .ZN(new_n777_));
  OAI21_X1  g576(.A(G106gat), .B1(new_n764_), .B2(new_n642_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n778_), .A2(KEYINPUT52), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(KEYINPUT52), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n777_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT53), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT53), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n777_), .B(new_n783_), .C1(new_n779_), .C2(new_n780_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1339gat));
  NOR2_X1   g584(.A1(new_n624_), .A2(new_n566_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n574_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n585_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n579_), .A2(new_n582_), .A3(new_n584_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n586_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n578_), .A2(KEYINPUT12), .B1(new_n265_), .B2(new_n302_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n793_), .A2(KEYINPUT55), .A3(new_n581_), .A4(new_n584_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n790_), .A2(new_n792_), .A3(new_n794_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n795_), .A2(KEYINPUT56), .A3(new_n596_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT119), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT56), .B1(new_n795_), .B2(new_n596_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n795_), .A2(new_n596_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n349_), .A2(new_n350_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n342_), .A2(new_n343_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n334_), .A2(new_n344_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n332_), .B1(new_n346_), .B2(new_n806_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n804_), .A2(new_n332_), .B1(new_n805_), .B2(new_n807_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n808_), .A2(new_n599_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n803_), .A2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n788_), .B1(new_n799_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n800_), .A2(new_n802_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(KEYINPUT119), .A3(new_n796_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n813_), .A2(KEYINPUT58), .A3(new_n803_), .A4(new_n809_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n811_), .A2(new_n653_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT57), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n597_), .A2(KEYINPUT72), .A3(new_n599_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n601_), .A2(new_n602_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n808_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT117), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n795_), .A2(new_n820_), .A3(new_n596_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT118), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n802_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n599_), .B1(new_n348_), .B2(new_n352_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT117), .B1(new_n822_), .B2(KEYINPUT56), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n825_), .B1(new_n800_), .B2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n819_), .B1(new_n824_), .B2(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n816_), .B1(new_n829_), .B2(new_n617_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n817_), .A2(new_n818_), .A3(new_n808_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n800_), .A2(new_n827_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n832_), .A2(new_n353_), .A3(new_n599_), .ZN(new_n833_));
  AOI21_X1  g632(.A(KEYINPUT56), .B1(new_n821_), .B2(new_n822_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n831_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n617_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(KEYINPUT57), .A3(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n815_), .A2(new_n830_), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT120), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n815_), .A2(new_n830_), .A3(new_n837_), .A4(KEYINPUT120), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n326_), .A3(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n713_), .A2(KEYINPUT116), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n353_), .B2(new_n326_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n610_), .A2(new_n843_), .A3(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT54), .B1(new_n846_), .B2(new_n653_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n843_), .A2(new_n845_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n610_), .A2(new_n849_), .A3(new_n850_), .A4(new_n295_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n847_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n787_), .B1(new_n842_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(G113gat), .B1(new_n853_), .B2(new_n353_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n853_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT59), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n787_), .A2(KEYINPUT59), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n847_), .A2(new_n851_), .ZN(new_n858_));
  AND2_X1   g657(.A1(new_n838_), .A2(new_n326_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n857_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n856_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n354_), .A2(KEYINPUT121), .ZN(new_n863_));
  MUX2_X1   g662(.A(KEYINPUT121), .B(new_n863_), .S(G113gat), .Z(new_n864_));
  AOI21_X1  g663(.A(new_n854_), .B1(new_n862_), .B2(new_n864_), .ZN(G1340gat));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n676_), .B(new_n860_), .C1(new_n853_), .C2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(G120gat), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n610_), .A2(KEYINPUT60), .ZN(new_n869_));
  MUX2_X1   g668(.A(new_n869_), .B(KEYINPUT60), .S(G120gat), .Z(new_n870_));
  NAND2_X1  g669(.A1(new_n853_), .A2(new_n870_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n868_), .A2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n868_), .A2(KEYINPUT122), .A3(new_n871_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1341gat));
  OAI21_X1  g675(.A(G127gat), .B1(new_n861_), .B2(new_n326_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n326_), .A2(G127gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n855_), .B2(new_n878_), .ZN(G1342gat));
  OAI21_X1  g678(.A(G134gat), .B1(new_n861_), .B2(new_n295_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n836_), .A2(G134gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n855_), .B2(new_n881_), .ZN(G1343gat));
  NAND2_X1  g681(.A1(new_n842_), .A2(new_n852_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n573_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n885_), .A2(new_n353_), .A3(new_n786_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g686(.A1(new_n885_), .A2(new_n676_), .A3(new_n786_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g688(.A1(new_n885_), .A2(new_n327_), .A3(new_n786_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT61), .B(G155gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  NOR3_X1   g691(.A1(new_n884_), .A2(new_n566_), .A3(new_n624_), .ZN(new_n893_));
  INV_X1    g692(.A(G162gat), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n893_), .A2(new_n894_), .A3(new_n617_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n893_), .A2(new_n653_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n894_), .ZN(G1347gat));
  NOR2_X1   g696(.A1(new_n858_), .A2(new_n859_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n682_), .A2(new_n620_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n574_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n354_), .A2(new_n456_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT124), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n464_), .B1(new_n901_), .B2(new_n353_), .ZN(new_n905_));
  XOR2_X1   g704(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n906_));
  AND2_X1   g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n905_), .A2(new_n906_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n904_), .B1(new_n907_), .B2(new_n908_), .ZN(G1348gat));
  AOI21_X1  g708(.A(G176gat), .B1(new_n901_), .B2(new_n676_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n546_), .B1(new_n842_), .B2(new_n852_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n899_), .ZN(new_n912_));
  NOR4_X1   g711(.A1(new_n912_), .A2(new_n610_), .A3(new_n462_), .A4(new_n656_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n910_), .B1(new_n911_), .B2(new_n913_), .ZN(G1349gat));
  NAND4_X1  g713(.A1(new_n911_), .A2(new_n563_), .A3(new_n327_), .A4(new_n899_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n326_), .A2(new_n443_), .ZN(new_n916_));
  AOI22_X1  g715(.A1(new_n915_), .A2(new_n451_), .B1(new_n901_), .B2(new_n916_), .ZN(G1350gat));
  NAND3_X1  g716(.A1(new_n901_), .A2(new_n444_), .A3(new_n617_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n452_), .B1(new_n901_), .B2(new_n653_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n919_), .A2(KEYINPUT125), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n919_), .A2(KEYINPUT125), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n918_), .B1(new_n920_), .B2(new_n921_), .ZN(G1351gat));
  NOR2_X1   g721(.A1(new_n884_), .A2(new_n912_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n353_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G197gat), .ZN(G1352gat));
  AOI21_X1  g724(.A(G204gat), .B1(new_n923_), .B2(new_n676_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n923_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n927_), .A2(new_n610_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n422_), .B2(new_n928_), .ZN(G1353gat));
  NAND2_X1  g728(.A1(new_n923_), .A2(new_n327_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n930_), .A2(KEYINPUT126), .A3(new_n931_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n884_), .A2(new_n326_), .A3(new_n912_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n931_), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n933_), .B1(new_n934_), .B2(new_n935_), .ZN(new_n936_));
  XOR2_X1   g735(.A(KEYINPUT63), .B(G211gat), .Z(new_n937_));
  AOI22_X1  g736(.A1(new_n932_), .A2(new_n936_), .B1(new_n934_), .B2(new_n937_), .ZN(G1354gat));
  OAI21_X1  g737(.A(G218gat), .B1(new_n927_), .B2(new_n295_), .ZN(new_n939_));
  INV_X1    g738(.A(G218gat), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n923_), .A2(new_n940_), .A3(new_n617_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n941_), .ZN(G1355gat));
endmodule


