//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:47 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n871_, new_n873_, new_n874_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G78gat), .B(G106gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G211gat), .B(G218gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(KEYINPUT92), .A2(G197gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(KEYINPUT92), .A2(G197gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(G204gat), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G197gat), .A2(G204gat), .ZN(new_n210_));
  INV_X1    g009(.A(new_n210_), .ZN(new_n211_));
  AND4_X1   g010(.A1(KEYINPUT21), .A2(new_n205_), .A3(new_n209_), .A4(new_n211_), .ZN(new_n212_));
  NOR3_X1   g011(.A1(new_n207_), .A2(new_n208_), .A3(G204gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT21), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n214_), .B1(G197gat), .B2(G204gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT93), .B1(new_n213_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT92), .ZN(new_n218_));
  INV_X1    g017(.A(G197gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G204gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(new_n221_), .A3(new_n206_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT93), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n215_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n217_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n209_), .A2(new_n211_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n205_), .B1(new_n226_), .B2(new_n214_), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n212_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT29), .ZN(new_n229_));
  INV_X1    g028(.A(G141gat), .ZN(new_n230_));
  INV_X1    g029(.A(G148gat), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n230_), .B(new_n231_), .C1(KEYINPUT87), .C2(KEYINPUT3), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT87), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n233_), .B(new_n234_), .C1(G141gat), .C2(G148gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G141gat), .A2(G148gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT86), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT86), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(G141gat), .A3(G148gat), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT2), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n238_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n237_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT2), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n236_), .A2(new_n242_), .A3(new_n244_), .ZN(new_n245_));
  AND2_X1   g044(.A1(G155gat), .A2(G162gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(G155gat), .A2(G162gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n230_), .A2(new_n231_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND4_X1  g053(.A1(new_n251_), .A2(new_n238_), .A3(new_n240_), .A4(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n229_), .B1(new_n249_), .B2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n203_), .B1(new_n228_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n220_), .A2(new_n206_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n210_), .B1(new_n258_), .B2(G204gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(KEYINPUT21), .A3(new_n205_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n222_), .A2(new_n223_), .A3(new_n215_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n223_), .B1(new_n222_), .B2(new_n215_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n204_), .B1(new_n259_), .B2(KEYINPUT21), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n260_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n248_), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n232_), .A2(new_n235_), .B1(new_n243_), .B2(KEYINPUT2), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n266_), .B1(new_n267_), .B2(new_n242_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n238_), .A2(new_n240_), .A3(new_n252_), .A4(new_n253_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n269_), .B1(new_n250_), .B2(new_n248_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT29), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n203_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n265_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n257_), .A2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(KEYINPUT90), .B(G228gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(KEYINPUT91), .B(G233gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n278_), .B1(new_n265_), .B2(KEYINPUT94), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n274_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(new_n257_), .A3(new_n273_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n281_), .A2(KEYINPUT89), .A3(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT88), .B(KEYINPUT28), .ZN(new_n284_));
  XOR2_X1   g083(.A(G22gat), .B(G50gat), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n249_), .A2(new_n255_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n285_), .B1(new_n286_), .B2(KEYINPUT29), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(new_n286_), .A2(KEYINPUT29), .A3(new_n285_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n284_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n289_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n284_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n292_), .A3(new_n287_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n290_), .A2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n283_), .A2(KEYINPUT95), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT95), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n279_), .A2(new_n257_), .A3(new_n273_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n265_), .A2(KEYINPUT94), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n257_), .A2(new_n273_), .B1(new_n298_), .B2(new_n277_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n296_), .B1(new_n300_), .B2(KEYINPUT89), .ZN(new_n301_));
  INV_X1    g100(.A(new_n294_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n281_), .A2(new_n296_), .A3(new_n282_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n295_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT99), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT96), .B(KEYINPUT19), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G226gat), .A2(G233gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT83), .ZN(new_n310_));
  INV_X1    g109(.A(G169gat), .ZN(new_n311_));
  INV_X1    g110(.A(G176gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT83), .B1(G169gat), .B2(G176gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT24), .B1(new_n311_), .B2(new_n312_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n313_), .A2(KEYINPUT24), .A3(new_n314_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT82), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT25), .B(G183gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT26), .ZN(new_n322_));
  OAI21_X1  g121(.A(KEYINPUT81), .B1(new_n322_), .B2(G190gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(G190gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT26), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(G190gat), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT81), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n320_), .B1(new_n324_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT81), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n322_), .A2(G190gat), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n325_), .A2(KEYINPUT26), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n330_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n333_), .A2(KEYINPUT82), .A3(new_n321_), .A4(new_n323_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT23), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(G183gat), .A3(G190gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n337_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n338_));
  AOI21_X1  g137(.A(KEYINPUT84), .B1(new_n337_), .B2(KEYINPUT23), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n336_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n319_), .A2(new_n329_), .A3(new_n334_), .A4(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G169gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n337_), .A2(KEYINPUT23), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n344_), .A2(new_n336_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n343_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n341_), .A2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT20), .B1(new_n348_), .B2(new_n265_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n340_), .B1(G183gat), .B2(G190gat), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n331_), .A2(new_n332_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n345_), .B1(new_n351_), .B2(new_n321_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n350_), .A2(new_n343_), .B1(new_n352_), .B2(new_n319_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n228_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n309_), .B1(new_n349_), .B2(new_n354_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G8gat), .B(G36gat), .Z(new_n356_));
  XNOR2_X1  g155(.A(G64gat), .B(G92gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT20), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n228_), .B2(new_n353_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n348_), .A2(new_n265_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n309_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n355_), .A2(new_n360_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT27), .ZN(new_n367_));
  INV_X1    g166(.A(new_n349_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n354_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n364_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n362_), .A2(new_n363_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n371_), .A2(new_n309_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n360_), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n306_), .B1(new_n367_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT27), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n355_), .A2(new_n360_), .A3(new_n365_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n360_), .B1(new_n355_), .B2(new_n365_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n360_), .ZN(new_n379_));
  NOR3_X1   g178(.A1(new_n349_), .A2(new_n309_), .A3(new_n354_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n364_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n379_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n382_), .A2(KEYINPUT99), .A3(KEYINPUT27), .A4(new_n366_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n305_), .A2(new_n374_), .A3(new_n378_), .A4(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G127gat), .B(G134gat), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  XOR2_X1   g186(.A(G113gat), .B(G120gat), .Z(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(G113gat), .B(G120gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n386_), .A2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n389_), .A2(KEYINPUT85), .A3(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n389_), .A2(new_n391_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT85), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n286_), .A2(new_n392_), .A3(new_n395_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n249_), .A2(new_n255_), .A3(new_n393_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n385_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n392_), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT85), .B1(new_n389_), .B2(new_n391_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(KEYINPUT4), .B1(new_n401_), .B2(new_n286_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n398_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n396_), .A2(new_n397_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n403_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G1gat), .B(G29gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT98), .B(KEYINPUT0), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G57gat), .B(G85gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  NOR3_X1   g211(.A1(new_n404_), .A2(new_n407_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G227gat), .A2(G233gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n416_), .B(G15gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT30), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n341_), .A2(new_n418_), .A3(new_n347_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n341_), .B2(new_n347_), .ZN(new_n420_));
  OR3_X1    g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n401_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G71gat), .B(G99gat), .ZN(new_n422_));
  INV_X1    g221(.A(G43gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT31), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n401_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n421_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n425_), .B1(new_n421_), .B2(new_n426_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n414_), .B(new_n415_), .C1(new_n427_), .C2(new_n428_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n202_), .B1(new_n384_), .B2(new_n429_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n374_), .A2(new_n378_), .A3(new_n383_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n429_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n431_), .A2(KEYINPUT100), .A3(new_n305_), .A4(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n430_), .A2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n427_), .A2(new_n428_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n374_), .A2(new_n378_), .A3(new_n383_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n283_), .A2(KEYINPUT95), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n437_), .A2(new_n303_), .A3(new_n302_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n412_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n405_), .A2(KEYINPUT4), .ZN(new_n440_));
  INV_X1    g239(.A(new_n403_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n396_), .A2(new_n385_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n439_), .B1(new_n443_), .B2(new_n406_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n413_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n438_), .A2(new_n445_), .A3(new_n295_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n436_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n441_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n439_), .B1(new_n405_), .B2(new_n403_), .ZN(new_n449_));
  OAI21_X1  g248(.A(KEYINPUT33), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(new_n415_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n376_), .A2(new_n377_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n444_), .A2(KEYINPUT33), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n360_), .A2(KEYINPUT32), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n355_), .A2(new_n365_), .A3(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n380_), .A2(new_n381_), .ZN(new_n457_));
  OAI221_X1 g256(.A(new_n456_), .B1(new_n457_), .B2(new_n455_), .C1(new_n413_), .C2(new_n444_), .ZN(new_n458_));
  AOI22_X1  g257(.A1(new_n454_), .A2(new_n458_), .B1(new_n438_), .B2(new_n295_), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n435_), .B1(new_n447_), .B2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n434_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G113gat), .B(G141gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT79), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G169gat), .B(G197gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(G29gat), .B(G36gat), .Z(new_n467_));
  XOR2_X1   g266(.A(G43gat), .B(G50gat), .Z(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G29gat), .B(G36gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G43gat), .B(G50gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT77), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G15gat), .B(G22gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT75), .B(G1gat), .ZN(new_n476_));
  INV_X1    g275(.A(G8gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT14), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n475_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G8gat), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n475_), .B(new_n481_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n474_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G229gat), .A2(G233gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n473_), .B(KEYINPUT15), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(KEYINPUT78), .B1(new_n490_), .B2(new_n485_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n485_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT78), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(new_n489_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n488_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT77), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n473_), .B(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n492_), .A2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n487_), .B1(new_n498_), .B2(new_n486_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n466_), .B1(new_n495_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n498_), .A2(new_n486_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n487_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n492_), .A2(new_n489_), .A3(new_n493_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n493_), .B1(new_n492_), .B2(new_n489_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n503_), .B(new_n465_), .C1(new_n506_), .C2(new_n488_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT80), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n500_), .A2(new_n507_), .A3(new_n508_), .ZN(new_n509_));
  OAI211_X1 g308(.A(KEYINPUT80), .B(new_n466_), .C1(new_n495_), .C2(new_n499_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(G230gat), .ZN(new_n513_));
  INV_X1    g312(.A(G233gat), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(G71gat), .B(G78gat), .Z(new_n516_));
  XNOR2_X1  g315(.A(G57gat), .B(G64gat), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n516_), .B1(KEYINPUT11), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT69), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n519_), .A3(KEYINPUT11), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n519_), .B1(new_n517_), .B2(KEYINPUT11), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n518_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n517_), .A2(KEYINPUT11), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT69), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n517_), .A2(KEYINPUT11), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n525_), .A2(new_n526_), .A3(new_n516_), .A4(new_n520_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G85gat), .B(G92gat), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n529_), .B1(KEYINPUT9), .B2(G92gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n531_));
  OR2_X1    g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n530_), .A2(new_n531_), .ZN(new_n533_));
  INV_X1    g332(.A(G99gat), .ZN(new_n534_));
  INV_X1    g333(.A(G106gat), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT6), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT6), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n537_), .A2(G99gat), .A3(G106gat), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  XOR2_X1   g338(.A(KEYINPUT10), .B(G99gat), .Z(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT64), .B(G106gat), .Z(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n532_), .A2(new_n533_), .A3(new_n539_), .A4(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT8), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n539_), .A2(KEYINPUT68), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT68), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n536_), .A2(new_n546_), .A3(new_n538_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT66), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT7), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n548_), .B(new_n549_), .C1(G99gat), .C2(G106gat), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n534_), .B(new_n535_), .C1(KEYINPUT66), .C2(KEYINPUT7), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n545_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n529_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n544_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n544_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n552_), .A2(new_n539_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT67), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT67), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n552_), .A2(new_n539_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n556_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n528_), .B(new_n543_), .C1(new_n555_), .C2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT70), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n560_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n559_), .B1(new_n552_), .B2(new_n539_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n539_), .A2(KEYINPUT68), .B1(new_n550_), .B2(new_n551_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n529_), .B1(new_n568_), .B2(new_n547_), .ZN(new_n569_));
  OAI22_X1  g368(.A1(new_n567_), .A2(new_n556_), .B1(new_n569_), .B2(new_n544_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n570_), .A2(KEYINPUT70), .A3(new_n543_), .A4(new_n528_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n564_), .A2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n528_), .B1(new_n570_), .B2(new_n543_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n515_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n562_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n543_), .B1(new_n555_), .B2(new_n561_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n528_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT71), .B(KEYINPUT12), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n577_), .A2(KEYINPUT12), .A3(new_n578_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n576_), .A2(new_n581_), .A3(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n574_), .A2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G120gat), .B(G148gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(G176gat), .B(G204gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n589_), .A2(KEYINPUT72), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n584_), .B(new_n590_), .ZN(new_n591_));
  OR2_X1    g390(.A1(new_n591_), .A2(KEYINPUT13), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(KEYINPUT13), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n485_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(new_n528_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT16), .ZN(new_n600_));
  XOR2_X1   g399(.A(G183gat), .B(G211gat), .Z(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n598_), .A2(KEYINPUT17), .A3(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n598_), .A2(KEYINPUT76), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(KEYINPUT17), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n606_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n604_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n577_), .A2(new_n489_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n570_), .A2(new_n473_), .A3(new_n543_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(G232gat), .A2(G233gat), .ZN(new_n612_));
  XOR2_X1   g411(.A(new_n612_), .B(KEYINPUT34), .Z(new_n613_));
  INV_X1    g412(.A(KEYINPUT35), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n610_), .A2(new_n611_), .A3(KEYINPUT74), .A4(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n613_), .A2(new_n614_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n617_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G190gat), .B(G218gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(new_n623_), .B(KEYINPUT36), .Z(new_n624_));
  NAND2_X1  g423(.A1(new_n620_), .A2(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n623_), .A2(KEYINPUT36), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n618_), .A2(new_n626_), .A3(new_n619_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n625_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n628_), .A2(KEYINPUT37), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT37), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n625_), .A2(new_n630_), .A3(new_n627_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n609_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n461_), .A2(new_n512_), .A3(new_n595_), .A4(new_n632_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT101), .Z(new_n634_));
  INV_X1    g433(.A(new_n445_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n635_), .A2(new_n476_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT102), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT102), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n634_), .A2(new_n639_), .A3(new_n636_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(KEYINPUT38), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n609_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n595_), .A2(new_n512_), .A3(new_n642_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT103), .ZN(new_n644_));
  INV_X1    g443(.A(new_n628_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n645_), .B1(new_n434_), .B2(new_n460_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G1gat), .B1(new_n647_), .B2(new_n445_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n641_), .A2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT38), .B1(new_n638_), .B2(new_n640_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1324gat));
  NAND3_X1  g450(.A1(new_n634_), .A2(new_n477_), .A3(new_n436_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n644_), .A2(new_n436_), .A3(new_n646_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n653_), .A2(new_n654_), .A3(G8gat), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n654_), .B1(new_n653_), .B2(G8gat), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n657_), .B(new_n659_), .ZN(G1325gat));
  OAI21_X1  g459(.A(G15gat), .B1(new_n647_), .B2(new_n435_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT41), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n633_), .A2(G15gat), .A3(new_n435_), .ZN(new_n663_));
  OR2_X1    g462(.A1(new_n662_), .A2(new_n663_), .ZN(G1326gat));
  OAI21_X1  g463(.A(G22gat), .B1(new_n647_), .B2(new_n305_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT42), .ZN(new_n666_));
  OR2_X1    g465(.A1(new_n305_), .A2(G22gat), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT105), .Z(new_n668_));
  OAI21_X1  g467(.A(new_n666_), .B1(new_n633_), .B2(new_n668_), .ZN(G1327gat));
  NOR3_X1   g468(.A1(new_n594_), .A2(new_n511_), .A3(new_n642_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n629_), .A2(new_n631_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n671_), .B1(new_n461_), .B2(new_n673_), .ZN(new_n674_));
  AOI211_X1 g473(.A(KEYINPUT43), .B(new_n672_), .C1(new_n434_), .C2(new_n460_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n670_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT44), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  OAI211_X1 g477(.A(KEYINPUT44), .B(new_n670_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n678_), .A2(new_n680_), .A3(new_n445_), .ZN(new_n681_));
  INV_X1    g480(.A(G29gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n511_), .B1(new_n434_), .B2(new_n460_), .ZN(new_n683_));
  NOR3_X1   g482(.A1(new_n594_), .A2(new_n642_), .A3(new_n628_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n635_), .A2(new_n682_), .ZN(new_n686_));
  OAI22_X1  g485(.A1(new_n681_), .A2(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT106), .ZN(G1328gat));
  NOR3_X1   g487(.A1(new_n685_), .A2(G36gat), .A3(new_n431_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT45), .Z(new_n690_));
  NAND2_X1  g489(.A1(new_n676_), .A2(new_n677_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n691_), .A2(new_n436_), .A3(new_n679_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(new_n693_), .A3(G36gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n692_), .B2(G36gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n690_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT46), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT46), .B(new_n690_), .C1(new_n694_), .C2(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(G1329gat));
  NOR2_X1   g499(.A1(new_n685_), .A2(new_n435_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n701_), .A2(G43gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n678_), .A2(new_n680_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n435_), .A2(new_n423_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n702_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT47), .Z(G1330gat));
  NOR2_X1   g505(.A1(new_n685_), .A2(new_n305_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(G50gat), .ZN(new_n708_));
  INV_X1    g507(.A(new_n305_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(G50gat), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n708_), .B1(new_n703_), .B2(new_n711_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT108), .Z(G1331gat));
  INV_X1    g512(.A(G57gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n512_), .B1(new_n434_), .B2(new_n460_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n594_), .A2(new_n632_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n714_), .B1(new_n717_), .B2(new_n445_), .ZN(new_n718_));
  XOR2_X1   g517(.A(new_n718_), .B(KEYINPUT109), .Z(new_n719_));
  NOR3_X1   g518(.A1(new_n595_), .A2(new_n512_), .A3(new_n609_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n720_), .A2(new_n646_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n721_), .A2(new_n714_), .A3(new_n445_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n719_), .A2(new_n722_), .ZN(G1332gat));
  OAI21_X1  g522(.A(G64gat), .B1(new_n721_), .B2(new_n431_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT48), .ZN(new_n725_));
  OR2_X1    g524(.A1(new_n431_), .A2(G64gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n717_), .B2(new_n726_), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n721_), .B2(new_n435_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT49), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n435_), .A2(G71gat), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n717_), .B2(new_n730_), .ZN(G1334gat));
  OAI21_X1  g530(.A(G78gat), .B1(new_n721_), .B2(new_n305_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT50), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n305_), .A2(G78gat), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n733_), .B1(new_n717_), .B2(new_n734_), .ZN(G1335gat));
  NOR2_X1   g534(.A1(new_n642_), .A2(new_n628_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n715_), .A2(new_n594_), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n635_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT110), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n674_), .A2(new_n675_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n594_), .A2(new_n511_), .A3(new_n609_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n635_), .A2(G85gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1336gat));
  AOI21_X1  g544(.A(G92gat), .B1(new_n738_), .B2(new_n436_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n436_), .A2(G92gat), .ZN(new_n747_));
  XOR2_X1   g546(.A(new_n747_), .B(KEYINPUT111), .Z(new_n748_));
  AOI21_X1  g547(.A(new_n746_), .B1(new_n743_), .B2(new_n748_), .ZN(G1337gat));
  INV_X1    g548(.A(new_n435_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n738_), .A2(new_n750_), .A3(new_n540_), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n741_), .A2(new_n435_), .A3(new_n742_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n752_), .B2(new_n534_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g553(.A(new_n541_), .ZN(new_n755_));
  NOR3_X1   g554(.A1(new_n737_), .A2(new_n305_), .A3(new_n755_), .ZN(new_n756_));
  NOR3_X1   g555(.A1(new_n741_), .A2(new_n305_), .A3(new_n742_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT52), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n759_), .A3(G106gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT52), .B1(new_n757_), .B2(new_n535_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n756_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n762_), .B(new_n764_), .ZN(G1339gat));
  NOR3_X1   g564(.A1(new_n384_), .A2(new_n445_), .A3(new_n435_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT58), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n501_), .A2(new_n487_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n769_), .A2(KEYINPUT115), .A3(new_n466_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT115), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n502_), .B1(new_n498_), .B2(new_n486_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(new_n465_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n486_), .A2(new_n502_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n770_), .B(new_n773_), .C1(new_n506_), .C2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n574_), .A2(new_n583_), .A3(new_n589_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n507_), .A3(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n580_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n582_), .B1(new_n573_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n515_), .B1(new_n779_), .B2(new_n572_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n779_), .B2(new_n575_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n576_), .A2(KEYINPUT55), .A3(new_n581_), .A4(new_n582_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n780_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n589_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n784_), .A2(KEYINPUT56), .A3(new_n785_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n777_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n768_), .B1(new_n790_), .B2(KEYINPUT117), .ZN(new_n791_));
  INV_X1    g590(.A(new_n777_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n784_), .A2(KEYINPUT56), .A3(new_n785_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT56), .B1(new_n784_), .B2(new_n785_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n792_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT117), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(new_n796_), .A3(KEYINPUT58), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n672_), .B1(new_n791_), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n509_), .A2(new_n510_), .A3(new_n776_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n801_));
  AND2_X1   g600(.A1(new_n574_), .A2(new_n583_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n802_), .A2(new_n590_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n590_), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n507_), .B(new_n775_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n645_), .B1(new_n801_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT116), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n807_), .A2(KEYINPUT57), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n808_), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n645_), .B(new_n810_), .C1(new_n801_), .C2(new_n805_), .ZN(new_n811_));
  OAI22_X1  g610(.A1(new_n798_), .A2(new_n799_), .B1(new_n809_), .B2(new_n811_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n795_), .A2(new_n796_), .A3(KEYINPUT58), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT58), .B1(new_n795_), .B2(new_n796_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n673_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n815_), .A2(KEYINPUT118), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n609_), .B1(new_n812_), .B2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT114), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n632_), .A2(new_n593_), .A3(new_n592_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n819_), .B1(new_n820_), .B2(new_n512_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n818_), .A2(KEYINPUT114), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n595_), .A2(new_n511_), .A3(new_n632_), .A4(new_n823_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n821_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n767_), .B1(new_n817_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n512_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT59), .B1(new_n767_), .B2(KEYINPUT119), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n806_), .B(new_n808_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n642_), .B1(new_n830_), .B2(new_n815_), .ZN(new_n831_));
  OAI221_X1 g630(.A(new_n829_), .B1(KEYINPUT119), .B2(new_n767_), .C1(new_n831_), .C2(new_n825_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n832_), .B(new_n833_), .C1(new_n827_), .C2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n815_), .A2(KEYINPUT118), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n798_), .A2(new_n799_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n837_), .A2(new_n838_), .A3(new_n830_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n825_), .B1(new_n839_), .B2(new_n609_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT59), .B1(new_n840_), .B2(new_n767_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n833_), .B1(new_n841_), .B2(new_n832_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n836_), .A2(new_n842_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n512_), .A2(G113gat), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n828_), .B1(new_n843_), .B2(new_n844_), .ZN(G1340gat));
  NAND3_X1  g644(.A1(new_n841_), .A2(new_n594_), .A3(new_n832_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G120gat), .ZN(new_n847_));
  INV_X1    g646(.A(new_n827_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT60), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n594_), .A2(new_n849_), .ZN(new_n850_));
  MUX2_X1   g649(.A(new_n850_), .B(new_n849_), .S(G120gat), .Z(new_n851_));
  OAI21_X1  g650(.A(new_n847_), .B1(new_n848_), .B2(new_n851_), .ZN(G1341gat));
  NOR3_X1   g651(.A1(new_n840_), .A2(new_n609_), .A3(new_n767_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT121), .B1(new_n853_), .B2(G127gat), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n827_), .A2(new_n642_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n856_));
  INV_X1    g655(.A(G127gat), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n855_), .A2(new_n856_), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n854_), .A2(new_n858_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT122), .B(G127gat), .Z(new_n860_));
  NOR2_X1   g659(.A1(new_n609_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n859_), .B1(new_n843_), .B2(new_n861_), .ZN(G1342gat));
  AOI21_X1  g661(.A(G134gat), .B1(new_n827_), .B2(new_n645_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n673_), .A2(G134gat), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n863_), .B1(new_n843_), .B2(new_n864_), .ZN(G1343gat));
  NOR2_X1   g664(.A1(new_n840_), .A2(new_n750_), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n436_), .A2(new_n445_), .A3(new_n305_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n511_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n230_), .ZN(G1344gat));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n595_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(new_n231_), .ZN(G1345gat));
  NOR2_X1   g671(.A1(new_n868_), .A2(new_n609_), .ZN(new_n873_));
  XOR2_X1   g672(.A(KEYINPUT61), .B(G155gat), .Z(new_n874_));
  XNOR2_X1  g673(.A(new_n873_), .B(new_n874_), .ZN(G1346gat));
  OAI21_X1  g674(.A(G162gat), .B1(new_n868_), .B2(new_n672_), .ZN(new_n876_));
  OR2_X1    g675(.A1(new_n628_), .A2(G162gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n868_), .B2(new_n877_), .ZN(G1347gat));
  OR2_X1    g677(.A1(new_n831_), .A2(new_n825_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n431_), .A2(new_n709_), .A3(new_n429_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(new_n512_), .A3(new_n880_), .ZN(new_n881_));
  XOR2_X1   g680(.A(KEYINPUT22), .B(G169gat), .Z(new_n882_));
  NOR2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(KEYINPUT123), .B1(new_n881_), .B2(G169gat), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n883_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n881_), .A2(G169gat), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT62), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n887_), .A2(new_n888_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n886_), .B1(new_n890_), .B2(new_n891_), .ZN(G1348gat));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n879_), .A2(new_n880_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n312_), .B1(new_n894_), .B2(new_n595_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n840_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n305_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n431_), .A2(new_n429_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n594_), .A2(G176gat), .A3(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n893_), .B1(new_n896_), .B2(new_n901_), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n895_), .B(KEYINPUT124), .C1(new_n898_), .C2(new_n900_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1349gat));
  NOR3_X1   g703(.A1(new_n894_), .A2(new_n321_), .A3(new_n609_), .ZN(new_n905_));
  NAND4_X1  g704(.A1(new_n897_), .A2(new_n305_), .A3(new_n642_), .A4(new_n899_), .ZN(new_n906_));
  INV_X1    g705(.A(G183gat), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n905_), .B1(new_n906_), .B2(new_n907_), .ZN(G1350gat));
  OAI21_X1  g707(.A(G190gat), .B1(new_n894_), .B2(new_n672_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n645_), .A2(new_n351_), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT125), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n879_), .A2(new_n880_), .A3(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n909_), .A2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n913_), .A2(new_n914_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n909_), .A2(KEYINPUT126), .A3(new_n912_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1351gat));
  NOR2_X1   g716(.A1(new_n431_), .A2(new_n446_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n866_), .A2(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n511_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(new_n219_), .ZN(G1352gat));
  NOR2_X1   g720(.A1(new_n919_), .A2(new_n595_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n922_), .B(new_n923_), .ZN(G1353gat));
  AOI21_X1  g723(.A(new_n609_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n866_), .A2(new_n918_), .A3(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  XOR2_X1   g726(.A(new_n926_), .B(new_n927_), .Z(G1354gat));
  OAI21_X1  g727(.A(G218gat), .B1(new_n919_), .B2(new_n672_), .ZN(new_n929_));
  OR2_X1    g728(.A1(new_n628_), .A2(G218gat), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n919_), .B2(new_n930_), .ZN(G1355gat));
endmodule


