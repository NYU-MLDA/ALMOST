//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 0 0 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n838_, new_n840_, new_n841_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_, new_n895_;
  INV_X1    g000(.A(KEYINPUT101), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G169gat), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n208_), .A2(KEYINPUT24), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n205_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G169gat), .A2(G176gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(KEYINPUT24), .A3(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NOR2_X1   g013(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT79), .B(G183gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n215_), .B1(new_n216_), .B2(KEYINPUT25), .ZN(new_n217_));
  OAI211_X1 g016(.A(new_n210_), .B(new_n212_), .C1(new_n214_), .C2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n211_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT22), .B(G169gat), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n219_), .B1(new_n220_), .B2(new_n207_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n216_), .A2(G190gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n221_), .B1(new_n222_), .B2(new_n205_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n218_), .A2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(new_n224_), .B(KEYINPUT80), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT30), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n224_), .B(KEYINPUT80), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT30), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NOR3_X1   g030(.A1(new_n227_), .A2(KEYINPUT82), .A3(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT83), .B(G127gat), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n233_), .B(G134gat), .ZN(new_n234_));
  XOR2_X1   g033(.A(G113gat), .B(G120gat), .Z(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n234_), .B(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT82), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n238_), .B1(new_n226_), .B2(new_n230_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G71gat), .B(G99gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G15gat), .B(G43gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G227gat), .A2(G233gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT81), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n242_), .B(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(KEYINPUT31), .B1(new_n239_), .B2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  NOR3_X1   g047(.A1(new_n239_), .A2(KEYINPUT31), .A3(new_n246_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n237_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n249_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n234_), .B(new_n235_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n251_), .A2(new_n247_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n232_), .B1(new_n250_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n250_), .A2(new_n253_), .A3(new_n232_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(G155gat), .ZN(new_n258_));
  INV_X1    g057(.A(G162gat), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n259_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(G141gat), .A2(G148gat), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n263_), .B(KEYINPUT3), .Z(new_n264_));
  NAND2_X1  g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n265_), .B(KEYINPUT2), .Z(new_n266_));
  OAI211_X1 g065(.A(new_n261_), .B(new_n262_), .C1(new_n264_), .C2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n265_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n268_), .A2(new_n263_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT1), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(G155gat), .A3(G162gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT84), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n262_), .B1(new_n260_), .B2(new_n270_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n269_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n267_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  OR3_X1    g075(.A1(new_n276_), .A2(new_n237_), .A3(KEYINPUT4), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n237_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n252_), .A2(new_n275_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n278_), .A2(new_n279_), .A3(KEYINPUT4), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G225gat), .A2(G233gat), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(new_n280_), .A3(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G57gat), .B(G85gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(G1gat), .B(G29gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n285_), .B(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n281_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n278_), .A2(new_n279_), .A3(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n282_), .A2(new_n287_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT93), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n282_), .A2(KEYINPUT93), .A3(new_n287_), .A4(new_n289_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G211gat), .B(G218gat), .Z(new_n295_));
  INV_X1    g094(.A(G197gat), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(G204gat), .ZN(new_n297_));
  INV_X1    g096(.A(G204gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(G197gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n295_), .B1(KEYINPUT21), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n297_), .B(KEYINPUT85), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n299_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n301_), .B1(new_n303_), .B2(KEYINPUT21), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n303_), .A2(KEYINPUT21), .A3(new_n295_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n224_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT88), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT20), .ZN(new_n309_));
  INV_X1    g108(.A(new_n306_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT25), .B(G183gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n213_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n212_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT87), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n210_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n221_), .B1(new_n205_), .B2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n310_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT89), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n309_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  AND2_X1   g120(.A1(new_n316_), .A2(new_n318_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(KEYINPUT89), .A3(new_n310_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G226gat), .A2(G233gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT19), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n308_), .A2(new_n321_), .A3(new_n323_), .A4(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n306_), .A2(new_n224_), .ZN(new_n328_));
  OAI211_X1 g127(.A(KEYINPUT20), .B(new_n328_), .C1(new_n322_), .C2(new_n310_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n325_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT18), .B(G64gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(G92gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(G8gat), .B(G36gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n327_), .A2(new_n330_), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n336_));
  NOR3_X1   g135(.A1(new_n294_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n277_), .A2(new_n280_), .A3(new_n288_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT90), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n278_), .A2(new_n279_), .A3(new_n281_), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n277_), .A2(new_n280_), .A3(KEYINPUT90), .A4(new_n288_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n287_), .ZN(new_n343_));
  NAND4_X1  g142(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .A4(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT33), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n345_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT92), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n344_), .A2(KEYINPUT92), .A3(new_n345_), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n337_), .A2(new_n346_), .A3(new_n349_), .A4(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n340_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(new_n287_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n344_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n308_), .A2(KEYINPUT20), .A3(new_n319_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n355_), .A2(new_n325_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n329_), .A2(new_n325_), .ZN(new_n357_));
  OAI211_X1 g156(.A(KEYINPUT32), .B(new_n334_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n334_), .A2(KEYINPUT32), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n327_), .A2(new_n330_), .A3(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n354_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT94), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT94), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n354_), .A2(new_n358_), .A3(new_n363_), .A4(new_n360_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n351_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  XOR2_X1   g164(.A(KEYINPUT86), .B(KEYINPUT29), .Z(new_n366_));
  OAI21_X1  g165(.A(new_n306_), .B1(new_n276_), .B2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(G228gat), .A3(G233gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G22gat), .B(G50gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT28), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G228gat), .A2(G233gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n306_), .B(new_n372_), .C1(new_n276_), .C2(new_n373_), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n368_), .A2(new_n371_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n371_), .B1(new_n368_), .B2(new_n374_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n276_), .A2(new_n373_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G78gat), .B(G106gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(new_n379_), .Z(new_n380_));
  NAND2_X1  g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n380_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n382_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n381_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n365_), .A2(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n327_), .A2(new_n330_), .A3(new_n334_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n357_), .B1(new_n355_), .B2(new_n325_), .ZN(new_n387_));
  OAI211_X1 g186(.A(KEYINPUT27), .B(new_n386_), .C1(new_n387_), .C2(new_n334_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT95), .B(KEYINPUT27), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n353_), .A2(new_n381_), .A3(new_n344_), .A4(new_n383_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT96), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n392_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT96), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n394_), .A2(new_n395_), .A3(new_n390_), .A4(new_n388_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n393_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n257_), .B1(new_n385_), .B2(new_n397_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n391_), .A2(KEYINPUT97), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n391_), .A2(KEYINPUT97), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n384_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n354_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n256_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n402_), .B1(new_n403_), .B2(new_n254_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n398_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G29gat), .B(G36gat), .ZN(new_n407_));
  INV_X1    g206(.A(G43gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(G50gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT15), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT64), .ZN(new_n413_));
  AND2_X1   g212(.A1(G85gat), .A2(G92gat), .ZN(new_n414_));
  NOR2_X1   g213(.A1(G85gat), .A2(G92gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT9), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G85gat), .A2(G92gat), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT9), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n413_), .B1(new_n416_), .B2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G99gat), .A2(G106gat), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(KEYINPUT10), .B(G99gat), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G106gat), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n426_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n416_), .A2(new_n413_), .A3(new_n419_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n421_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT8), .ZN(new_n433_));
  INV_X1    g232(.A(new_n425_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n437_));
  OAI211_X1 g236(.A(KEYINPUT65), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n439_));
  INV_X1    g238(.A(G99gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n429_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n436_), .A2(new_n437_), .A3(new_n438_), .A4(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n414_), .A2(new_n415_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n433_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n424_), .A2(new_n437_), .A3(new_n425_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n441_), .A2(new_n438_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n433_), .B(new_n443_), .C1(new_n445_), .C2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n432_), .B1(new_n444_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n412_), .A2(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n416_), .A2(new_n413_), .A3(new_n419_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n451_), .A2(new_n420_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n443_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT8), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n430_), .A2(new_n452_), .B1(new_n454_), .B2(new_n447_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n411_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n450_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G232gat), .A2(G233gat), .ZN(new_n458_));
  XOR2_X1   g257(.A(new_n458_), .B(KEYINPUT72), .Z(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT34), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(KEYINPUT35), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(KEYINPUT35), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n460_), .A2(KEYINPUT35), .ZN(new_n463_));
  NAND4_X1  g262(.A1(new_n450_), .A2(new_n462_), .A3(new_n463_), .A4(new_n456_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G190gat), .B(G218gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(G134gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(G162gat), .ZN(new_n468_));
  OAI22_X1  g267(.A1(new_n465_), .A2(KEYINPUT73), .B1(KEYINPUT36), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT73), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n468_), .A2(KEYINPUT36), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n461_), .A2(new_n470_), .A3(new_n464_), .A4(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n465_), .A2(KEYINPUT36), .A3(new_n468_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G15gat), .B(G22gat), .Z(new_n478_));
  NAND2_X1  g277(.A1(G1gat), .A2(G8gat), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n478_), .B1(KEYINPUT14), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT74), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n481_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n479_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(G1gat), .A2(G8gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n484_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n482_), .A2(new_n487_), .A3(new_n483_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G231gat), .A2(G233gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(G57gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(KEYINPUT66), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT66), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G57gat), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n495_), .A2(new_n497_), .A3(G64gat), .ZN(new_n498_));
  AOI21_X1  g297(.A(G64gat), .B1(new_n495_), .B2(new_n497_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT11), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G71gat), .A2(G78gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(G71gat), .A2(G78gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n501_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  OR2_X1    g304(.A1(G71gat), .A2(G78gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT67), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(KEYINPUT11), .A4(new_n502_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(KEYINPUT11), .A3(new_n502_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT67), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n500_), .A2(new_n505_), .B1(new_n508_), .B2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n508_), .ZN(new_n512_));
  INV_X1    g311(.A(G64gat), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n496_), .A2(G57gat), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n494_), .A2(KEYINPUT66), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n513_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n495_), .A2(new_n497_), .A3(G64gat), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n505_), .A3(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n512_), .A2(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n511_), .A2(new_n519_), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n493_), .B(new_n520_), .Z(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT68), .ZN(new_n522_));
  XNOR2_X1  g321(.A(KEYINPUT16), .B(G183gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(G211gat), .ZN(new_n524_));
  XOR2_X1   g323(.A(G127gat), .B(G155gat), .Z(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT17), .ZN(new_n527_));
  XOR2_X1   g326(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n528_));
  NOR2_X1   g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  AOI22_X1  g328(.A1(new_n522_), .A2(new_n527_), .B1(new_n521_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n473_), .A2(new_n474_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT37), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n477_), .A2(new_n530_), .A3(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n406_), .A2(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n500_), .A2(new_n508_), .A3(new_n510_), .A4(new_n505_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n512_), .A2(new_n518_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(KEYINPUT12), .A3(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(KEYINPUT70), .B1(new_n455_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n449_), .A2(new_n520_), .A3(new_n539_), .A4(KEYINPUT12), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT68), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n542_), .B1(new_n511_), .B2(new_n519_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n535_), .A2(KEYINPUT68), .A3(new_n536_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n449_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT12), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(G230gat), .A2(G233gat), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n543_), .A2(new_n544_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n455_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n541_), .A2(new_n547_), .A3(new_n548_), .A4(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(KEYINPUT69), .A3(new_n545_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT69), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n549_), .A2(new_n553_), .A3(new_n455_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n551_), .B1(new_n555_), .B2(new_n548_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT71), .B(G204gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G120gat), .B(G148gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT5), .B(G176gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n556_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT13), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G229gat), .A2(G233gat), .ZN(new_n567_));
  INV_X1    g366(.A(new_n490_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n487_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n411_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n409_), .B(G50gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT15), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n567_), .B(new_n570_), .C1(new_n572_), .C2(new_n491_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n489_), .A2(new_n571_), .A3(new_n490_), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n570_), .A2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n573_), .B1(new_n575_), .B2(new_n567_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G113gat), .B(G141gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n206_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(new_n296_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT76), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT77), .Z(new_n581_));
  XNOR2_X1  g380(.A(new_n576_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT78), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n566_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n534_), .A2(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n585_), .A2(G1gat), .A3(new_n402_), .ZN(new_n586_));
  OR3_X1    g385(.A1(new_n586_), .A2(KEYINPUT100), .A3(KEYINPUT38), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT100), .B1(new_n586_), .B2(KEYINPUT38), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n406_), .A2(new_n531_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n566_), .A2(new_n582_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n530_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT99), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n591_), .A2(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n595_), .B2(new_n402_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n586_), .A2(new_n597_), .A3(KEYINPUT38), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n597_), .B1(new_n586_), .B2(KEYINPUT38), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n596_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n202_), .B1(new_n590_), .B2(new_n600_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n598_), .A2(new_n599_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n602_), .A2(KEYINPUT101), .A3(new_n596_), .A4(new_n589_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(G1324gat));
  OR2_X1    g403(.A1(new_n399_), .A2(new_n400_), .ZN(new_n605_));
  OR3_X1    g404(.A1(new_n585_), .A2(G8gat), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n605_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n591_), .A2(new_n607_), .A3(new_n594_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n609_), .A3(G8gat), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n609_), .B1(new_n608_), .B2(G8gat), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n606_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT102), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT102), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n615_), .B(new_n606_), .C1(new_n611_), .C2(new_n612_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n614_), .A2(KEYINPUT40), .A3(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT40), .B1(new_n614_), .B2(new_n616_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n617_), .A2(new_n618_), .ZN(G1325gat));
  INV_X1    g418(.A(new_n257_), .ZN(new_n620_));
  OAI21_X1  g419(.A(G15gat), .B1(new_n595_), .B2(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n621_), .B(KEYINPUT103), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT41), .ZN(new_n623_));
  INV_X1    g422(.A(new_n585_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(new_n257_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n623_), .B1(G15gat), .B2(new_n625_), .ZN(G1326gat));
  OAI21_X1  g425(.A(G22gat), .B1(new_n595_), .B2(new_n384_), .ZN(new_n627_));
  XOR2_X1   g426(.A(new_n627_), .B(KEYINPUT42), .Z(new_n628_));
  NOR3_X1   g427(.A1(new_n585_), .A2(G22gat), .A3(new_n384_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1327gat));
  NOR2_X1   g429(.A1(new_n406_), .A2(new_n475_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n530_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n632_), .A3(new_n584_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(new_n402_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT43), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n393_), .A2(new_n396_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n636_), .B1(new_n384_), .B2(new_n365_), .ZN(new_n637_));
  OAI22_X1  g436(.A1(new_n637_), .A2(new_n257_), .B1(new_n401_), .B2(new_n404_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n477_), .A2(new_n532_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n635_), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n635_), .B(new_n639_), .C1(new_n398_), .C2(new_n405_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n592_), .B(new_n632_), .C1(new_n640_), .C2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT44), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n639_), .ZN(new_n646_));
  OAI21_X1  g445(.A(KEYINPUT43), .B1(new_n406_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(new_n641_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n648_), .A2(KEYINPUT44), .A3(new_n592_), .A4(new_n632_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n645_), .A2(new_n354_), .A3(new_n649_), .ZN(new_n650_));
  MUX2_X1   g449(.A(new_n634_), .B(new_n650_), .S(G29gat), .Z(G1328gat));
  NAND3_X1  g450(.A1(new_n645_), .A2(new_n607_), .A3(new_n649_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(G36gat), .ZN(new_n653_));
  NAND4_X1  g452(.A1(new_n631_), .A2(new_n607_), .A3(new_n632_), .A4(new_n584_), .ZN(new_n654_));
  OR3_X1    g453(.A1(new_n654_), .A2(KEYINPUT45), .A3(G36gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT45), .B1(new_n654_), .B2(G36gat), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(KEYINPUT105), .A2(KEYINPUT46), .ZN(new_n658_));
  AOI22_X1  g457(.A1(new_n653_), .A2(new_n657_), .B1(KEYINPUT104), .B2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n653_), .A2(KEYINPUT104), .A3(new_n657_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT105), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT46), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(G1329gat));
  NAND4_X1  g462(.A1(new_n645_), .A2(G43gat), .A3(new_n649_), .A4(new_n257_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n408_), .B1(new_n633_), .B2(new_n620_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g466(.A(new_n384_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n645_), .A2(G50gat), .A3(new_n649_), .A4(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n410_), .B1(new_n633_), .B2(new_n384_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1331gat));
  AND2_X1   g470(.A1(new_n564_), .A2(new_n565_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n582_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n534_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G57gat), .B1(new_n676_), .B2(new_n354_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n591_), .A2(new_n566_), .A3(new_n530_), .A4(new_n583_), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n678_), .A2(new_n494_), .A3(new_n402_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1332gat));
  OAI21_X1  g479(.A(G64gat), .B1(new_n678_), .B2(new_n605_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT48), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n605_), .A2(G64gat), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT106), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n682_), .B1(new_n675_), .B2(new_n684_), .ZN(G1333gat));
  OAI21_X1  g484(.A(G71gat), .B1(new_n678_), .B2(new_n620_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT49), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n620_), .A2(G71gat), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT107), .Z(new_n689_));
  OAI21_X1  g488(.A(new_n687_), .B1(new_n675_), .B2(new_n689_), .ZN(G1334gat));
  INV_X1    g489(.A(G78gat), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n672_), .A2(new_n384_), .A3(new_n673_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n534_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G78gat), .B1(new_n678_), .B2(new_n384_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n694_), .A2(KEYINPUT108), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(KEYINPUT108), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n695_), .A2(KEYINPUT50), .A3(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT50), .B1(new_n695_), .B2(new_n696_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n693_), .B1(new_n697_), .B2(new_n698_), .ZN(G1335gat));
  NOR3_X1   g498(.A1(new_n672_), .A2(new_n530_), .A3(new_n673_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n631_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G85gat), .B1(new_n702_), .B2(new_n354_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT109), .B1(new_n640_), .B2(new_n642_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT109), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n647_), .A2(new_n705_), .A3(new_n641_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n707_), .A2(new_n354_), .A3(new_n700_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n703_), .B1(new_n708_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g508(.A(G92gat), .B1(new_n702_), .B2(new_n607_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n707_), .A2(G92gat), .A3(new_n700_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n711_), .B2(new_n607_), .ZN(G1337gat));
  NAND4_X1  g511(.A1(new_n704_), .A2(new_n706_), .A3(new_n257_), .A4(new_n700_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n713_), .A2(KEYINPUT110), .A3(G99gat), .ZN(new_n714_));
  AOI21_X1  g513(.A(KEYINPUT110), .B1(new_n713_), .B2(G99gat), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n714_), .A2(new_n715_), .A3(KEYINPUT111), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT51), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n702_), .A2(new_n257_), .A3(new_n428_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n716_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n715_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT111), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n713_), .A2(KEYINPUT110), .A3(G99gat), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n720_), .A2(new_n721_), .A3(new_n722_), .A4(new_n718_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT51), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n719_), .A2(new_n724_), .ZN(G1338gat));
  NAND3_X1  g524(.A1(new_n702_), .A2(new_n429_), .A3(new_n668_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT52), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n530_), .B1(new_n647_), .B2(new_n641_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n692_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n727_), .B1(new_n729_), .B2(G106gat), .ZN(new_n730_));
  AOI211_X1 g529(.A(KEYINPUT52), .B(new_n429_), .C1(new_n728_), .C2(new_n692_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n726_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(new_n732_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g532(.A(KEYINPUT55), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n551_), .A2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(KEYINPUT113), .ZN(new_n736_));
  AOI22_X1  g535(.A1(new_n538_), .A2(new_n540_), .B1(new_n549_), .B2(new_n455_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n737_), .A2(KEYINPUT55), .A3(new_n548_), .A4(new_n547_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n541_), .A2(new_n547_), .A3(new_n550_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(G230gat), .A3(G233gat), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT113), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n551_), .A2(new_n741_), .A3(new_n734_), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n736_), .A2(new_n738_), .A3(new_n740_), .A4(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT114), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n740_), .A2(new_n738_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n746_), .A2(KEYINPUT114), .A3(new_n736_), .A4(new_n742_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n745_), .A2(new_n561_), .A3(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(KEYINPUT56), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n556_), .A2(new_n561_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT56), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n745_), .A2(new_n751_), .A3(new_n561_), .A4(new_n747_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n749_), .A2(new_n750_), .A3(new_n673_), .A4(new_n752_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n576_), .A2(new_n579_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n755_));
  INV_X1    g554(.A(new_n567_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n755_), .B(new_n579_), .C1(new_n575_), .C2(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n570_), .B2(new_n574_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n579_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT115), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n757_), .A2(new_n760_), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n756_), .B(new_n570_), .C1(new_n572_), .C2(new_n491_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n754_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n763_), .A2(new_n562_), .A3(KEYINPUT116), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(KEYINPUT116), .B1(new_n763_), .B2(new_n562_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n753_), .A2(new_n767_), .ZN(new_n768_));
  AOI21_X1  g567(.A(KEYINPUT57), .B1(new_n768_), .B2(new_n475_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  AOI211_X1 g569(.A(new_n770_), .B(new_n531_), .C1(new_n753_), .C2(new_n767_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n769_), .A2(new_n771_), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n749_), .A2(new_n750_), .A3(new_n752_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(KEYINPUT58), .A4(new_n763_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n749_), .A2(new_n750_), .A3(new_n752_), .A4(new_n763_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT58), .ZN(new_n777_));
  AOI22_X1  g576(.A1(new_n776_), .A2(new_n777_), .B1(new_n477_), .B2(new_n532_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT117), .B1(new_n776_), .B2(new_n777_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n530_), .B1(new_n772_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n672_), .A2(new_n583_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(KEYINPUT112), .A2(KEYINPUT54), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  OR4_X1    g585(.A1(new_n533_), .A2(new_n782_), .A3(new_n783_), .A4(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n784_), .B(new_n785_), .C1(new_n533_), .C2(new_n782_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT118), .B1(new_n781_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n768_), .A2(new_n475_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(new_n770_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n768_), .A2(KEYINPUT57), .A3(new_n475_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n780_), .A2(new_n792_), .A3(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n632_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT118), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n787_), .A2(new_n788_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n795_), .A2(new_n796_), .A3(new_n797_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n620_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n790_), .A2(new_n798_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT59), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT59), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n802_), .B(new_n799_), .C1(new_n781_), .C2(new_n789_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n801_), .A2(G113gat), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n583_), .ZN(new_n805_));
  INV_X1    g604(.A(G113gat), .ZN(new_n806_));
  AND2_X1   g605(.A1(new_n790_), .A2(new_n798_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(new_n673_), .A3(new_n799_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n804_), .A2(new_n805_), .B1(new_n806_), .B2(new_n808_), .ZN(G1340gat));
  INV_X1    g608(.A(G120gat), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n672_), .B2(KEYINPUT60), .ZN(new_n811_));
  OR2_X1    g610(.A1(new_n810_), .A2(KEYINPUT60), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n807_), .A2(new_n799_), .A3(new_n811_), .A4(new_n812_), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n801_), .A2(new_n566_), .A3(new_n803_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n810_), .ZN(G1341gat));
  NAND4_X1  g614(.A1(new_n801_), .A2(G127gat), .A3(new_n530_), .A4(new_n803_), .ZN(new_n816_));
  INV_X1    g615(.A(G127gat), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n800_), .B2(new_n632_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(KEYINPUT119), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n816_), .A2(new_n821_), .A3(new_n818_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n820_), .A2(new_n822_), .ZN(G1342gat));
  NAND3_X1  g622(.A1(new_n807_), .A2(new_n531_), .A3(new_n799_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT120), .ZN(new_n825_));
  INV_X1    g624(.A(G134gat), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n824_), .A2(new_n825_), .A3(new_n826_), .ZN(new_n827_));
  AND4_X1   g626(.A1(G134gat), .A2(new_n801_), .A3(new_n639_), .A4(new_n803_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n825_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n827_), .A2(new_n828_), .A3(new_n829_), .ZN(G1343gat));
  NAND4_X1  g629(.A1(new_n790_), .A2(new_n798_), .A3(new_n605_), .A4(new_n620_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n402_), .A2(new_n384_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n673_), .ZN(new_n835_));
  XNOR2_X1  g634(.A(KEYINPUT121), .B(G141gat), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(G1344gat));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n566_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g638(.A1(new_n834_), .A2(new_n530_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT61), .B(G155gat), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n840_), .B(new_n841_), .ZN(G1346gat));
  NOR3_X1   g641(.A1(new_n831_), .A2(new_n475_), .A3(new_n833_), .ZN(new_n843_));
  OAI21_X1  g642(.A(KEYINPUT122), .B1(new_n843_), .B2(G162gat), .ZN(new_n844_));
  AND3_X1   g643(.A1(new_n790_), .A2(new_n798_), .A3(new_n620_), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n845_), .A2(new_n605_), .A3(new_n531_), .A4(new_n832_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT122), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n259_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n646_), .A2(new_n259_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n844_), .A2(new_n848_), .B1(new_n834_), .B2(new_n849_), .ZN(G1347gat));
  NOR2_X1   g649(.A1(new_n605_), .A2(new_n404_), .ZN(new_n851_));
  OAI211_X1 g650(.A(new_n384_), .B(new_n851_), .C1(new_n781_), .C2(new_n789_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n673_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G169gat), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(KEYINPUT123), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n854_), .A2(new_n857_), .A3(G169gat), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(KEYINPUT62), .A3(new_n858_), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n853_), .A2(new_n220_), .A3(new_n673_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT62), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n855_), .A2(KEYINPUT123), .A3(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n859_), .A2(new_n860_), .A3(new_n862_), .ZN(G1348gat));
  AOI21_X1  g662(.A(G176gat), .B1(new_n853_), .B2(new_n566_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n807_), .A2(new_n384_), .ZN(new_n865_));
  NOR4_X1   g664(.A1(new_n605_), .A2(new_n404_), .A3(new_n207_), .A4(new_n672_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(G1349gat));
  NOR3_X1   g666(.A1(new_n852_), .A2(new_n311_), .A3(new_n632_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n865_), .A2(new_n530_), .A3(new_n851_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n216_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n868_), .B1(new_n869_), .B2(new_n870_), .ZN(G1350gat));
  OAI21_X1  g670(.A(G190gat), .B1(new_n852_), .B2(new_n646_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n531_), .A2(new_n213_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n852_), .B2(new_n873_), .ZN(G1351gat));
  NOR2_X1   g673(.A1(new_n605_), .A2(new_n392_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n790_), .A2(new_n798_), .A3(new_n620_), .A4(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n582_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT124), .B(G197gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1352gat));
  NOR2_X1   g678(.A1(new_n298_), .A2(KEYINPUT125), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n876_), .A2(new_n672_), .A3(new_n880_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n298_), .A2(KEYINPUT125), .ZN(new_n882_));
  XOR2_X1   g681(.A(new_n882_), .B(KEYINPUT126), .Z(new_n883_));
  XOR2_X1   g682(.A(new_n881_), .B(new_n883_), .Z(G1353gat));
  XOR2_X1   g683(.A(KEYINPUT63), .B(G211gat), .Z(new_n885_));
  NAND4_X1  g684(.A1(new_n845_), .A2(new_n530_), .A3(new_n875_), .A4(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT127), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n876_), .B2(new_n632_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT127), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n888_), .B1(new_n886_), .B2(new_n891_), .ZN(G1354gat));
  NOR2_X1   g691(.A1(new_n876_), .A2(new_n475_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n893_), .A2(G218gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n876_), .A2(new_n646_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(G218gat), .B2(new_n895_), .ZN(G1355gat));
endmodule


