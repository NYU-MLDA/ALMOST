//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT0), .B(G57gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  NAND2_X1  g004(.A1(G225gat), .A2(G233gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT79), .ZN(new_n207_));
  INV_X1    g006(.A(G141gat), .ZN(new_n208_));
  INV_X1    g007(.A(G148gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT3), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n211_), .B1(G141gat), .B2(G148gat), .ZN(new_n212_));
  AND2_X1   g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n207_), .B1(new_n213_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n210_), .A2(new_n212_), .ZN(new_n219_));
  AND3_X1   g018(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(new_n214_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n221_), .A3(KEYINPUT79), .ZN(new_n222_));
  OR2_X1    g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n218_), .A2(new_n222_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n224_), .A2(KEYINPUT1), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(G155gat), .A3(G162gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n230_), .A3(new_n223_), .ZN(new_n231_));
  AND2_X1   g030(.A1(G141gat), .A2(G148gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(G141gat), .A2(G148gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n231_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT78), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n231_), .A2(KEYINPUT78), .A3(new_n234_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n227_), .A2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G127gat), .B(G134gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G113gat), .B(G120gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT77), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n241_), .B(new_n242_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n245_), .B1(new_n246_), .B2(new_n244_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n240_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n219_), .A2(new_n221_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n225_), .B1(new_n249_), .B2(new_n207_), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n250_), .A2(new_n222_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n246_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n248_), .A2(new_n252_), .A3(KEYINPUT4), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT87), .B(KEYINPUT4), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n240_), .A2(new_n247_), .A3(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n206_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n206_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n257_), .B1(new_n248_), .B2(new_n252_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n205_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT88), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT33), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT33), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n259_), .A2(new_n260_), .A3(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n265_));
  AND2_X1   g064(.A1(G226gat), .A2(G233gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT84), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT21), .ZN(new_n270_));
  AND2_X1   g069(.A1(G197gat), .A2(G204gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(G197gat), .A2(G204gat), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(G197gat), .ZN(new_n274_));
  INV_X1    g073(.A(G204gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G197gat), .A2(G204gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n276_), .A2(KEYINPUT21), .A3(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G211gat), .B(G218gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n273_), .A2(new_n278_), .A3(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT80), .ZN(new_n281_));
  INV_X1    g080(.A(G218gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(G211gat), .ZN(new_n283_));
  INV_X1    g082(.A(G211gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(G218gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n286_), .A2(KEYINPUT21), .A3(new_n276_), .A4(new_n277_), .ZN(new_n287_));
  AND3_X1   g086(.A1(new_n280_), .A2(new_n281_), .A3(new_n287_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n281_), .B1(new_n280_), .B2(new_n287_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G169gat), .ZN(new_n291_));
  INV_X1    g090(.A(G176gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n292_), .A3(KEYINPUT73), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT73), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n294_), .B1(G169gat), .B2(G176gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT24), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT26), .B(G190gat), .ZN(new_n299_));
  INV_X1    g098(.A(G183gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT25), .B1(new_n300_), .B2(KEYINPUT72), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT25), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(new_n303_), .A3(G183gat), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n299_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n293_), .A2(new_n295_), .A3(KEYINPUT24), .A4(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n298_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT74), .B(KEYINPUT23), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT75), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n313_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT75), .B1(new_n311_), .B2(KEYINPUT23), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n312_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(G183gat), .A2(G190gat), .ZN(new_n321_));
  AOI211_X1 g120(.A(new_n320_), .B(new_n321_), .C1(new_n309_), .C2(new_n313_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n291_), .A2(KEYINPUT22), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n292_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G169gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n291_), .A2(KEYINPUT22), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT76), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n306_), .B1(new_n325_), .B2(new_n329_), .ZN(new_n330_));
  OAI22_X1  g129(.A1(new_n308_), .A2(new_n319_), .B1(new_n322_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT20), .B1(new_n290_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n280_), .A2(new_n287_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  AND2_X1   g133(.A1(KEYINPUT74), .A2(KEYINPUT23), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n313_), .B1(new_n335_), .B2(new_n314_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(KEYINPUT23), .B2(new_n313_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT24), .B1(new_n293_), .B2(new_n295_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT85), .B1(new_n337_), .B2(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n320_), .B1(new_n309_), .B2(new_n313_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT85), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n298_), .A3(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT25), .B(G183gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n299_), .A2(new_n343_), .ZN(new_n344_));
  AND2_X1   g143(.A1(new_n344_), .A2(new_n307_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n339_), .A2(new_n342_), .A3(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT22), .B(G169gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(new_n292_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n306_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT86), .ZN(new_n350_));
  INV_X1    g149(.A(new_n321_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n312_), .B(new_n351_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT86), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n348_), .A2(new_n353_), .A3(new_n306_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n350_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n334_), .B1(new_n346_), .B2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n269_), .B1(new_n332_), .B2(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G8gat), .B(G36gat), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT18), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G64gat), .B(G92gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n359_), .B(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n290_), .A2(new_n331_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n346_), .A2(new_n355_), .A3(new_n334_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n362_), .A2(new_n363_), .A3(KEYINPUT20), .A4(new_n267_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n357_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n361_), .B1(new_n357_), .B2(new_n364_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n248_), .A2(new_n252_), .A3(KEYINPUT89), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n257_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT89), .B1(new_n248_), .B2(new_n252_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n205_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT90), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n253_), .A2(new_n374_), .A3(new_n206_), .A4(new_n255_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n253_), .A2(new_n206_), .A3(new_n255_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT90), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n372_), .A2(new_n373_), .A3(new_n375_), .A4(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n262_), .A2(new_n264_), .A3(new_n368_), .A4(new_n378_), .ZN(new_n379_));
  OR3_X1    g178(.A1(new_n256_), .A2(new_n205_), .A3(new_n258_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(new_n259_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n361_), .A2(KEYINPUT32), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n357_), .A2(new_n382_), .A3(new_n364_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT91), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n362_), .A2(new_n363_), .A3(KEYINPUT20), .ZN(new_n385_));
  INV_X1    g184(.A(new_n267_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  OR2_X1    g186(.A1(new_n290_), .A2(new_n331_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n346_), .A2(new_n355_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n333_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n388_), .A2(new_n390_), .A3(KEYINPUT20), .A4(new_n268_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n387_), .A2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(KEYINPUT32), .A3(new_n361_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n381_), .A2(new_n384_), .A3(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n379_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n240_), .A2(KEYINPUT29), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n333_), .ZN(new_n397_));
  AND2_X1   g196(.A1(G228gat), .A2(G233gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n288_), .A2(new_n289_), .A3(new_n398_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n396_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G22gat), .B(G50gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT28), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT29), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(new_n251_), .B2(new_n406_), .ZN(new_n407_));
  AND4_X1   g206(.A1(new_n405_), .A2(new_n227_), .A3(new_n239_), .A4(new_n406_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n404_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G78gat), .B(G106gat), .Z(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT81), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n227_), .A2(new_n239_), .A3(new_n406_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT28), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n251_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n404_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n409_), .A2(new_n411_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n411_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n420_), .B1(new_n409_), .B2(new_n416_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n403_), .B1(new_n417_), .B2(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n415_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n419_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n409_), .A2(new_n411_), .A3(new_n416_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n402_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n422_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n395_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT27), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n365_), .A2(KEYINPUT92), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT92), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n357_), .A2(new_n434_), .A3(new_n364_), .A4(new_n361_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n361_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n430_), .B1(new_n392_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(KEYINPUT93), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT93), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n436_), .A2(new_n441_), .A3(new_n438_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n432_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n422_), .A2(new_n380_), .A3(new_n259_), .A4(new_n427_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n443_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n429_), .A2(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G71gat), .B(G99gat), .ZN(new_n448_));
  INV_X1    g247(.A(G43gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  OR2_X1    g249(.A1(new_n331_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n331_), .A2(new_n450_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n453_), .A2(new_n247_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n453_), .A2(new_n247_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G227gat), .A2(G233gat), .ZN(new_n456_));
  INV_X1    g255(.A(G15gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n458_), .B(KEYINPUT30), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT31), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  OR3_X1    g260(.A1(new_n454_), .A2(new_n455_), .A3(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n461_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n436_), .A2(new_n441_), .A3(new_n438_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n441_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n428_), .B(new_n431_), .C1(new_n465_), .C2(new_n466_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n464_), .A2(new_n381_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT94), .B1(new_n467_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT94), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n443_), .A2(new_n471_), .A3(new_n428_), .A4(new_n468_), .ZN(new_n472_));
  AOI22_X1  g271(.A1(new_n447_), .A2(new_n464_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G1gat), .B(G8gat), .Z(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G15gat), .B(G22gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT70), .ZN(new_n477_));
  INV_X1    g276(.A(G1gat), .ZN(new_n478_));
  INV_X1    g277(.A(G8gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT14), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n476_), .A2(new_n477_), .A3(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n477_), .B1(new_n476_), .B2(new_n480_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n475_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n483_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(new_n481_), .A3(new_n474_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G29gat), .B(G36gat), .Z(new_n487_));
  XOR2_X1   g286(.A(G43gat), .B(G50gat), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G29gat), .B(G36gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G43gat), .B(G50gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n484_), .A2(new_n486_), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G229gat), .A2(G233gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT15), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n493_), .B(new_n496_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n484_), .A2(new_n486_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n494_), .B(new_n495_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n495_), .ZN(new_n500_));
  AND3_X1   g299(.A1(new_n484_), .A2(new_n486_), .A3(new_n493_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n493_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n499_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G113gat), .B(G141gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G169gat), .B(G197gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(new_n505_), .B(new_n506_), .Z(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n504_), .A2(new_n508_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n499_), .A2(new_n503_), .A3(new_n507_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AND2_X1   g311(.A1(G230gat), .A2(G233gat), .ZN(new_n513_));
  INV_X1    g312(.A(G85gat), .ZN(new_n514_));
  INV_X1    g313(.A(G92gat), .ZN(new_n515_));
  OAI21_X1  g314(.A(KEYINPUT64), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  AOI22_X1  g315(.A1(new_n516_), .A2(KEYINPUT9), .B1(new_n514_), .B2(new_n515_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT9), .ZN(new_n518_));
  OAI211_X1 g317(.A(KEYINPUT64), .B(new_n518_), .C1(new_n514_), .C2(new_n515_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G99gat), .A2(G106gat), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT6), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT10), .B(G99gat), .Z(new_n526_));
  INV_X1    g325(.A(G106gat), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n520_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT7), .ZN(new_n530_));
  INV_X1    g329(.A(G99gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n527_), .ZN(new_n532_));
  OAI21_X1  g331(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n532_), .A2(new_n523_), .A3(new_n524_), .A4(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT8), .ZN(new_n535_));
  XOR2_X1   g334(.A(G85gat), .B(G92gat), .Z(new_n536_));
  NAND3_X1  g335(.A1(new_n534_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(new_n535_), .B1(new_n534_), .B2(new_n536_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n529_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G57gat), .B(G64gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G71gat), .B(G78gat), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n541_), .A2(new_n542_), .A3(KEYINPUT11), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n544_));
  INV_X1    g343(.A(new_n542_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n541_), .A2(KEYINPUT11), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n543_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT65), .B1(new_n540_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n534_), .A2(new_n536_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT8), .ZN(new_n552_));
  AOI22_X1  g351(.A1(new_n552_), .A2(new_n537_), .B1(new_n528_), .B2(new_n520_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT65), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n548_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n550_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n553_), .A2(new_n548_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n513_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n559_));
  NOR2_X1   g358(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n560_));
  OAI22_X1  g359(.A1(new_n553_), .A2(new_n548_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n513_), .B1(new_n553_), .B2(new_n548_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n560_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n540_), .A2(new_n549_), .A3(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n561_), .A2(new_n562_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n558_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G120gat), .B(G148gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT5), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G176gat), .B(G204gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n568_), .B(new_n569_), .Z(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n570_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n558_), .A2(new_n565_), .A3(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT13), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(KEYINPUT67), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(KEYINPUT67), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n473_), .A2(new_n512_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n553_), .A2(new_n493_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT34), .ZN(new_n583_));
  OAI221_X1 g382(.A(new_n581_), .B1(KEYINPUT35), .B2(new_n583_), .C1(new_n553_), .C2(new_n497_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n583_), .A2(KEYINPUT35), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n584_), .A2(new_n585_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G190gat), .B(G218gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(G134gat), .B(G162gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT68), .B(KEYINPUT69), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(new_n593_), .B(KEYINPUT36), .Z(new_n594_));
  NAND2_X1  g393(.A1(new_n588_), .A2(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(KEYINPUT36), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n586_), .A2(new_n596_), .A3(new_n587_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT37), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT37), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n595_), .A2(new_n600_), .A3(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n548_), .B(new_n604_), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(new_n498_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT17), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G183gat), .B(G211gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(KEYINPUT71), .B(KEYINPUT16), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  OR3_X1    g411(.A1(new_n606_), .A2(new_n607_), .A3(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(KEYINPUT17), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n606_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n603_), .A2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n580_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n478_), .A3(new_n381_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT38), .ZN(new_n620_));
  INV_X1    g419(.A(new_n381_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n598_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n473_), .A2(new_n622_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n579_), .A2(new_n616_), .A3(new_n512_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT95), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n623_), .A2(new_n624_), .A3(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n621_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n620_), .B1(new_n478_), .B2(new_n629_), .ZN(G1324gat));
  INV_X1    g429(.A(new_n443_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n618_), .A2(new_n479_), .A3(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(G8gat), .B1(new_n625_), .B2(new_n443_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(KEYINPUT39), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(KEYINPUT39), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n632_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT40), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(G1325gat));
  INV_X1    g437(.A(new_n464_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n618_), .A2(new_n457_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n626_), .A2(new_n628_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n457_), .B1(new_n641_), .B2(new_n639_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n642_), .A2(KEYINPUT41), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(KEYINPUT41), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n643_), .B2(new_n644_), .ZN(G1326gat));
  INV_X1    g444(.A(G22gat), .ZN(new_n646_));
  INV_X1    g445(.A(new_n428_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n618_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n428_), .B1(new_n626_), .B2(new_n628_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(new_n646_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n649_), .A2(KEYINPUT42), .A3(new_n646_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n648_), .B1(new_n652_), .B2(new_n653_), .ZN(G1327gat));
  INV_X1    g453(.A(new_n616_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n598_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT96), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n580_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(G29gat), .B1(new_n659_), .B2(new_n381_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n579_), .A2(new_n655_), .A3(new_n512_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT43), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n470_), .A2(new_n472_), .ZN(new_n663_));
  AOI211_X1 g462(.A(new_n432_), .B(new_n444_), .C1(new_n440_), .C2(new_n442_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n647_), .B1(new_n379_), .B2(new_n394_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n464_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n663_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n662_), .B1(new_n667_), .B2(new_n603_), .ZN(new_n668_));
  AOI211_X1 g467(.A(KEYINPUT43), .B(new_n602_), .C1(new_n663_), .C2(new_n666_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n661_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT43), .B1(new_n473_), .B2(new_n602_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n667_), .A2(new_n662_), .A3(new_n603_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(KEYINPUT44), .A3(new_n661_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n672_), .A2(new_n676_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n381_), .A2(G29gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n660_), .B1(new_n677_), .B2(new_n678_), .ZN(G1328gat));
  NAND3_X1  g478(.A1(new_n672_), .A2(new_n676_), .A3(new_n631_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G36gat), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n443_), .A2(G36gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n580_), .A2(new_n657_), .A3(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT45), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT46), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n681_), .A2(new_n684_), .A3(KEYINPUT46), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(G1329gat));
  NOR2_X1   g488(.A1(new_n464_), .A2(new_n449_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n672_), .A2(new_n676_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT97), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT97), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n672_), .A2(new_n676_), .A3(new_n693_), .A4(new_n690_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n449_), .B1(new_n658_), .B2(new_n464_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n692_), .A2(new_n694_), .A3(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT47), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT47), .ZN(new_n698_));
  NAND4_X1  g497(.A1(new_n692_), .A2(new_n698_), .A3(new_n694_), .A4(new_n695_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1330gat));
  OR3_X1    g499(.A1(new_n658_), .A2(G50gat), .A3(new_n428_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n672_), .A2(new_n676_), .A3(new_n647_), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n702_), .A2(KEYINPUT98), .A3(G50gat), .ZN(new_n703_));
  AOI21_X1  g502(.A(KEYINPUT98), .B1(new_n702_), .B2(G50gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n701_), .B1(new_n703_), .B2(new_n704_), .ZN(G1331gat));
  NOR2_X1   g504(.A1(new_n616_), .A2(new_n511_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n623_), .A2(new_n579_), .A3(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT100), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(G57gat), .A3(new_n381_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT101), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n579_), .A2(new_n617_), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT99), .Z(new_n712_));
  NOR2_X1   g511(.A1(new_n473_), .A2(new_n511_), .ZN(new_n713_));
  AND2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n381_), .ZN(new_n715_));
  INV_X1    g514(.A(G57gat), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n715_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT101), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n708_), .A2(new_n718_), .A3(G57gat), .A4(new_n381_), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n710_), .A2(new_n717_), .A3(new_n719_), .ZN(G1332gat));
  NOR2_X1   g519(.A1(new_n443_), .A2(G64gat), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT102), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n714_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n708_), .A2(new_n631_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n725_), .B2(G64gat), .ZN(new_n726_));
  INV_X1    g525(.A(G64gat), .ZN(new_n727_));
  AOI211_X1 g526(.A(KEYINPUT48), .B(new_n727_), .C1(new_n708_), .C2(new_n631_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n723_), .B1(new_n726_), .B2(new_n728_), .ZN(G1333gat));
  INV_X1    g528(.A(G71gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n714_), .A2(new_n730_), .A3(new_n639_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n708_), .A2(new_n639_), .ZN(new_n732_));
  XNOR2_X1  g531(.A(KEYINPUT103), .B(KEYINPUT49), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(G71gat), .A3(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n732_), .B2(G71gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n731_), .B1(new_n734_), .B2(new_n735_), .ZN(G1334gat));
  INV_X1    g535(.A(G78gat), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n647_), .A2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT104), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n714_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n708_), .A2(new_n647_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n741_), .B1(new_n742_), .B2(G78gat), .ZN(new_n743_));
  AOI211_X1 g542(.A(KEYINPUT50), .B(new_n737_), .C1(new_n708_), .C2(new_n647_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n743_), .B2(new_n744_), .ZN(G1335gat));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n616_), .A2(new_n512_), .ZN(new_n747_));
  OR3_X1    g546(.A1(new_n578_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n746_), .B1(new_n578_), .B2(new_n747_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n675_), .A2(new_n750_), .ZN(new_n751_));
  OAI21_X1  g550(.A(G85gat), .B1(new_n751_), .B2(new_n621_), .ZN(new_n752_));
  AND3_X1   g551(.A1(new_n713_), .A2(new_n579_), .A3(new_n657_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(new_n514_), .A3(new_n381_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1336gat));
  NAND4_X1  g554(.A1(new_n675_), .A2(G92gat), .A3(new_n631_), .A4(new_n750_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n631_), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n757_), .A2(KEYINPUT106), .A3(new_n515_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT106), .B1(new_n757_), .B2(new_n515_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n756_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT107), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT107), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n756_), .B(new_n762_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1337gat));
  NAND3_X1  g563(.A1(new_n753_), .A2(new_n526_), .A3(new_n639_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n751_), .A2(new_n464_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n531_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g567(.A1(new_n753_), .A2(new_n527_), .A3(new_n647_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n675_), .A2(new_n647_), .A3(new_n750_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(new_n771_), .A3(G106gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(G106gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(KEYINPUT108), .B(KEYINPUT53), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n769_), .B(new_n775_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1339gat));
  INV_X1    g578(.A(KEYINPUT111), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n561_), .A2(new_n564_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n513_), .B1(new_n781_), .B2(new_n556_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n565_), .A2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n561_), .A2(new_n562_), .A3(new_n564_), .A4(KEYINPUT55), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n784_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(new_n570_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n494_), .B(new_n500_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n495_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n792_), .A3(new_n508_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n510_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n510_), .A2(new_n793_), .A3(KEYINPUT110), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n786_), .A2(new_n789_), .A3(new_n570_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n573_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n780_), .B1(new_n790_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT58), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n780_), .B(new_n803_), .C1(new_n790_), .C2(new_n800_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n802_), .A2(new_n603_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n574_), .A2(new_n798_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(KEYINPUT109), .A2(KEYINPUT56), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n788_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n807_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n511_), .B(new_n573_), .C1(new_n787_), .C2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n806_), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n598_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT113), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n805_), .A2(new_n814_), .A3(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n811_), .A2(KEYINPUT57), .A3(new_n598_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT112), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n811_), .A2(new_n819_), .A3(KEYINPUT57), .A4(new_n598_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n816_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n815_), .B1(new_n805_), .B2(new_n814_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n616_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n602_), .A2(new_n575_), .A3(new_n706_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT54), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT54), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n602_), .A2(new_n827_), .A3(new_n575_), .A4(new_n706_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n824_), .A2(new_n829_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n467_), .A2(new_n621_), .A3(new_n464_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT59), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n830_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n602_), .B1(KEYINPUT58), .B2(new_n801_), .ZN(new_n836_));
  AOI22_X1  g635(.A1(new_n836_), .A2(new_n804_), .B1(new_n813_), .B2(new_n812_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n655_), .B1(new_n837_), .B2(new_n821_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n829_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n831_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n835_), .B1(new_n832_), .B2(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(G113gat), .B1(new_n842_), .B2(new_n512_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n512_), .A2(G113gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n843_), .B1(new_n840_), .B2(new_n844_), .ZN(G1340gat));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n842_), .B2(new_n578_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n830_), .A2(new_n834_), .B1(new_n840_), .B2(KEYINPUT59), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n848_), .A2(KEYINPUT114), .A3(new_n579_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n847_), .A2(G120gat), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(G120gat), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n578_), .B2(KEYINPUT60), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n841_), .B(new_n852_), .C1(KEYINPUT60), .C2(new_n851_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n850_), .A2(new_n853_), .ZN(G1341gat));
  AOI21_X1  g653(.A(G127gat), .B1(new_n841_), .B2(new_n655_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n655_), .A2(G127gat), .ZN(new_n856_));
  XOR2_X1   g655(.A(new_n856_), .B(KEYINPUT115), .Z(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n848_), .B2(new_n857_), .ZN(G1342gat));
  OAI21_X1  g657(.A(G134gat), .B1(new_n842_), .B2(new_n602_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n840_), .A2(G134gat), .A3(new_n598_), .ZN(new_n860_));
  INV_X1    g659(.A(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n859_), .A2(KEYINPUT116), .A3(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863_));
  INV_X1    g662(.A(G134gat), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n864_), .B1(new_n848_), .B2(new_n603_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n865_), .B2(new_n860_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n862_), .A2(new_n866_), .ZN(G1343gat));
  NAND2_X1  g666(.A1(new_n837_), .A2(new_n821_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n839_), .B1(new_n868_), .B2(new_n616_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n647_), .A2(new_n464_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n631_), .A2(new_n621_), .A3(new_n871_), .ZN(new_n872_));
  XOR2_X1   g671(.A(new_n872_), .B(KEYINPUT117), .Z(new_n873_));
  NAND2_X1  g672(.A1(new_n870_), .A2(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT118), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n870_), .A2(KEYINPUT118), .A3(new_n873_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G141gat), .B1(new_n879_), .B2(new_n512_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n878_), .A2(new_n208_), .A3(new_n511_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1344gat));
  OAI21_X1  g681(.A(G148gat), .B1(new_n879_), .B2(new_n578_), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n878_), .A2(new_n209_), .A3(new_n579_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1345gat));
  XNOR2_X1  g684(.A(KEYINPUT61), .B(G155gat), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n879_), .B2(new_n616_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n886_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n878_), .A2(new_n655_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n889_), .ZN(G1346gat));
  OAI21_X1  g689(.A(G162gat), .B1(new_n879_), .B2(new_n602_), .ZN(new_n891_));
  INV_X1    g690(.A(G162gat), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n878_), .A2(new_n892_), .A3(new_n622_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1347gat));
  INV_X1    g693(.A(KEYINPUT119), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n443_), .A2(new_n469_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n428_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n824_), .B2(new_n829_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n898_), .A2(new_n347_), .A3(new_n511_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n291_), .B1(new_n898_), .B2(new_n511_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(KEYINPUT62), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n902_));
  AOI211_X1 g701(.A(new_n902_), .B(new_n291_), .C1(new_n898_), .C2(new_n511_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n895_), .B1(new_n901_), .B2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n898_), .A2(new_n511_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(G169gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n902_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n900_), .A2(KEYINPUT62), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n907_), .A2(KEYINPUT119), .A3(new_n908_), .A4(new_n899_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n904_), .A2(new_n909_), .ZN(G1348gat));
  AOI21_X1  g709(.A(G176gat), .B1(new_n898_), .B2(new_n579_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n870_), .A2(new_n428_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n579_), .A2(G176gat), .A3(new_n896_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n911_), .A2(new_n914_), .ZN(G1349gat));
  NAND2_X1  g714(.A1(new_n896_), .A2(new_n655_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n300_), .B1(new_n912_), .B2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n898_), .ZN(new_n918_));
  OR2_X1    g717(.A1(new_n616_), .A2(new_n343_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n917_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT120), .ZN(G1350gat));
  OAI21_X1  g720(.A(G190gat), .B1(new_n918_), .B2(new_n602_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n898_), .A2(new_n622_), .A3(new_n299_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(G1351gat));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT121), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n443_), .A2(new_n381_), .A3(new_n871_), .ZN(new_n927_));
  INV_X1    g726(.A(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n926_), .B1(new_n869_), .B2(new_n928_), .ZN(new_n929_));
  OAI211_X1 g728(.A(KEYINPUT121), .B(new_n927_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n512_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n925_), .B1(new_n931_), .B2(G197gat), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(G197gat), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n931_), .A2(new_n925_), .A3(G197gat), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n934_), .A2(new_n935_), .ZN(G1352gat));
  NAND2_X1  g735(.A1(new_n929_), .A2(new_n930_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n937_), .A2(new_n579_), .ZN(new_n938_));
  XOR2_X1   g737(.A(KEYINPUT123), .B(G204gat), .Z(new_n939_));
  XNOR2_X1  g738(.A(new_n938_), .B(new_n939_), .ZN(G1353gat));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n616_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n937_), .B2(new_n942_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n942_), .ZN(new_n945_));
  AOI211_X1 g744(.A(KEYINPUT124), .B(new_n945_), .C1(new_n929_), .C2(new_n930_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  NOR2_X1   g746(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n944_), .A2(new_n947_), .A3(new_n948_), .ZN(new_n949_));
  OAI22_X1  g748(.A1(new_n943_), .A2(new_n946_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n949_), .A2(new_n950_), .ZN(G1354gat));
  AOI21_X1  g750(.A(new_n598_), .B1(new_n929_), .B2(new_n930_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(KEYINPUT125), .ZN(new_n953_));
  XOR2_X1   g752(.A(KEYINPUT126), .B(G218gat), .Z(new_n954_));
  NOR2_X1   g753(.A1(new_n602_), .A2(new_n954_), .ZN(new_n955_));
  XOR2_X1   g754(.A(new_n955_), .B(KEYINPUT127), .Z(new_n956_));
  AOI22_X1  g755(.A1(new_n953_), .A2(new_n954_), .B1(new_n937_), .B2(new_n956_), .ZN(G1355gat));
endmodule


