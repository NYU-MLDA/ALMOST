//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n861_, new_n862_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n902_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_;
  OR2_X1    g000(.A1(G169gat), .A2(G176gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G169gat), .A2(G176gat), .ZN(new_n203_));
  NAND3_X1  g002(.A1(new_n202_), .A2(KEYINPUT24), .A3(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT80), .Z(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT25), .B(G183gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT26), .B(G190gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n202_), .A2(KEYINPUT24), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT23), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT23), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G183gat), .A3(G190gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n209_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n205_), .A2(new_n208_), .A3(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(new_n212_), .B2(new_n210_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n217_), .B1(new_n212_), .B2(new_n210_), .ZN(new_n218_));
  OAI21_X1  g017(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n218_), .B(new_n219_), .C1(KEYINPUT22), .C2(new_n202_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G71gat), .B(G99gat), .Z(new_n222_));
  XNOR2_X1  g021(.A(G15gat), .B(G43gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n222_), .B(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n221_), .B(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n226_));
  XOR2_X1   g025(.A(new_n225_), .B(new_n226_), .Z(new_n227_));
  XNOR2_X1  g026(.A(G127gat), .B(G134gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G113gat), .B(G120gat), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT82), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(new_n229_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(new_n232_), .B(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(G227gat), .A2(G233gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT81), .ZN(new_n236_));
  XOR2_X1   g035(.A(new_n236_), .B(KEYINPUT30), .Z(new_n237_));
  XNOR2_X1  g036(.A(new_n234_), .B(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n227_), .B(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G155gat), .A2(G162gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(G155gat), .A2(G162gat), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT86), .ZN(new_n244_));
  OR3_X1    g043(.A1(new_n242_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n244_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(G141gat), .ZN(new_n248_));
  INV_X1    g047(.A(G148gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n248_), .A2(new_n249_), .A3(KEYINPUT3), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n251_), .B1(G141gat), .B2(G148gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  AND3_X1   g052(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT85), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n253_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n257_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n247_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT87), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  OAI211_X1 g061(.A(KEYINPUT87), .B(new_n247_), .C1(new_n258_), .C2(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(G141gat), .A2(G148gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n248_), .A2(new_n249_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n241_), .A2(KEYINPUT1), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n241_), .B1(new_n243_), .B2(KEYINPUT1), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT84), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  OAI211_X1 g069(.A(KEYINPUT84), .B(new_n241_), .C1(new_n243_), .C2(KEYINPUT1), .ZN(new_n271_));
  AOI211_X1 g070(.A(new_n265_), .B(new_n266_), .C1(new_n270_), .C2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n234_), .B1(new_n264_), .B2(new_n273_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n230_), .A2(new_n233_), .ZN(new_n275_));
  AOI211_X1 g074(.A(new_n272_), .B(new_n275_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n276_));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(G225gat), .A2(G233gat), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n253_), .A2(new_n256_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(KEYINPUT85), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n253_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT87), .B1(new_n283_), .B2(new_n247_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n263_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n273_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n234_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT4), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n277_), .A2(new_n279_), .A3(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n278_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G1gat), .B(G29gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(G85gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(KEYINPUT0), .B(G57gat), .ZN(new_n296_));
  XOR2_X1   g095(.A(new_n295_), .B(new_n296_), .Z(new_n297_));
  NAND2_X1  g096(.A1(new_n293_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n297_), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n291_), .A2(new_n299_), .A3(new_n292_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(KEYINPUT99), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT99), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n291_), .A2(new_n302_), .A3(new_n299_), .A4(new_n292_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n240_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT27), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT91), .ZN(new_n307_));
  INV_X1    g106(.A(G218gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G211gat), .ZN(new_n309_));
  INV_X1    g108(.A(G211gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(G218gat), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n309_), .A2(new_n311_), .A3(KEYINPUT90), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT90), .B1(new_n309_), .B2(new_n311_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n307_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT90), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n310_), .A2(G218gat), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n308_), .A2(G211gat), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n315_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n309_), .A2(new_n311_), .A3(KEYINPUT90), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n318_), .A2(KEYINPUT91), .A3(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G197gat), .B(G204gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT21), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n314_), .A2(new_n320_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT92), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT92), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n314_), .A2(new_n320_), .A3(new_n326_), .A4(new_n323_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n321_), .A2(new_n322_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT89), .ZN(new_n331_));
  INV_X1    g130(.A(G197gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(G204gat), .ZN(new_n333_));
  INV_X1    g132(.A(G204gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(G197gat), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n333_), .A2(new_n335_), .A3(KEYINPUT88), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT21), .B1(new_n333_), .B2(KEYINPUT88), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n331_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n321_), .A2(KEYINPUT88), .ZN(new_n339_));
  OR2_X1    g138(.A1(new_n333_), .A2(KEYINPUT88), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n339_), .A2(KEYINPUT89), .A3(new_n340_), .A4(KEYINPUT21), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n330_), .B1(new_n338_), .B2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n328_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT93), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n342_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT93), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n346_), .A2(new_n348_), .A3(new_n221_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(G226gat), .A2(G233gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT19), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT22), .B(G169gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n353_), .A2(G176gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n203_), .B(KEYINPUT98), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n354_), .A2(new_n218_), .A3(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT97), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n214_), .B(new_n357_), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n208_), .A2(new_n204_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n356_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n351_), .B1(new_n360_), .B2(new_n347_), .ZN(new_n361_));
  AND3_X1   g160(.A1(new_n349_), .A2(KEYINPUT20), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n351_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n221_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n347_), .A2(KEYINPUT93), .ZN(new_n365_));
  AOI211_X1 g164(.A(new_n345_), .B(new_n342_), .C1(new_n325_), .C2(new_n327_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n360_), .A2(new_n347_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n363_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n362_), .A2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G8gat), .B(G36gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT18), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G64gat), .B(G92gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  AOI21_X1  g175(.A(new_n306_), .B1(new_n372_), .B2(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n376_), .B(KEYINPUT100), .Z(new_n378_));
  NOR2_X1   g177(.A1(new_n365_), .A2(new_n366_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n369_), .B1(new_n379_), .B2(new_n221_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT94), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n344_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n347_), .A2(KEYINPUT94), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n382_), .A2(new_n360_), .A3(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n363_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n367_), .A2(new_n370_), .A3(new_n363_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n378_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n377_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n376_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(new_n362_), .B2(new_n371_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n349_), .A2(KEYINPUT20), .A3(new_n361_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n367_), .A2(new_n370_), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n376_), .B(new_n391_), .C1(new_n392_), .C2(new_n363_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(KEYINPUT101), .B(KEYINPUT27), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n388_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n286_), .A2(KEYINPUT29), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n347_), .A2(KEYINPUT94), .ZN(new_n399_));
  AOI211_X1 g198(.A(new_n381_), .B(new_n342_), .C1(new_n325_), .C2(new_n327_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n398_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(G228gat), .ZN(new_n402_));
  INV_X1    g201(.A(G233gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n404_), .B1(new_n286_), .B2(KEYINPUT29), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n379_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G78gat), .B(G106gat), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n405_), .A2(KEYINPUT95), .A3(new_n407_), .A4(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G22gat), .B(G50gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n272_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT28), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n414_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n412_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n418_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(new_n416_), .A3(new_n411_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  AND2_X1   g221(.A1(new_n410_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n404_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n382_), .A2(new_n383_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n424_), .B1(new_n425_), .B2(new_n398_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n406_), .A2(new_n346_), .A3(new_n348_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n408_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT95), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n405_), .A2(new_n409_), .A3(new_n407_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n423_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(KEYINPUT96), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT96), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n405_), .A2(new_n434_), .A3(new_n407_), .A4(new_n409_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n422_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n433_), .A2(new_n435_), .A3(new_n428_), .A4(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n432_), .A2(new_n437_), .ZN(new_n438_));
  NOR3_X1   g237(.A1(new_n305_), .A2(new_n397_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n376_), .A2(KEYINPUT32), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n440_), .B(new_n391_), .C1(new_n392_), .C2(new_n363_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n380_), .A2(new_n384_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n386_), .B1(new_n442_), .B2(new_n351_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n441_), .B1(new_n443_), .B2(new_n440_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT33), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n445_), .B1(new_n293_), .B2(new_n297_), .ZN(new_n446_));
  AOI211_X1 g245(.A(KEYINPUT33), .B(new_n299_), .C1(new_n291_), .C2(new_n292_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n288_), .B(new_n279_), .C1(new_n286_), .C2(new_n275_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n277_), .A2(new_n290_), .ZN(new_n450_));
  OAI211_X1 g249(.A(new_n299_), .B(new_n449_), .C1(new_n450_), .C2(new_n279_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(new_n390_), .A3(new_n393_), .ZN(new_n452_));
  OAI22_X1  g251(.A1(new_n304_), .A2(new_n444_), .B1(new_n448_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n438_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n432_), .A2(new_n437_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n456_));
  AOI22_X1  g255(.A1(new_n387_), .A2(new_n377_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n455_), .A2(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n439_), .B1(new_n459_), .B2(new_n239_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G229gat), .A2(G233gat), .ZN(new_n461_));
  XOR2_X1   g260(.A(new_n461_), .B(KEYINPUT77), .Z(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT74), .B(G8gat), .ZN(new_n464_));
  INV_X1    g263(.A(G1gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT14), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT75), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G15gat), .B(G22gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G1gat), .B(G8gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n469_), .B(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G29gat), .B(G36gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G43gat), .B(G50gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n463_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n475_), .B(KEYINPUT15), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n471_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n476_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n471_), .B(new_n475_), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n479_), .B1(new_n480_), .B2(new_n461_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G113gat), .B(G141gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G169gat), .B(G197gat), .ZN(new_n483_));
  XOR2_X1   g282(.A(new_n482_), .B(new_n483_), .Z(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n481_), .A2(KEYINPUT78), .A3(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(KEYINPUT78), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n479_), .B(new_n487_), .C1(new_n480_), .C2(new_n461_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT79), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n460_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G57gat), .B(G64gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT11), .ZN(new_n493_));
  XOR2_X1   g292(.A(G71gat), .B(G78gat), .Z(new_n494_));
  OR2_X1    g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n492_), .A2(KEYINPUT11), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n494_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n495_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n498_), .A2(KEYINPUT68), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(KEYINPUT68), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(KEYINPUT12), .A3(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n502_));
  NAND2_X1  g301(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G99gat), .ZN(new_n505_));
  INV_X1    g304(.A(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G99gat), .A2(G106gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT6), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n503_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT65), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT8), .ZN(new_n514_));
  XOR2_X1   g313(.A(G85gat), .B(G92gat), .Z(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(new_n514_), .A3(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n508_), .A2(KEYINPUT66), .A3(new_n511_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT66), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n502_), .A2(new_n503_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n511_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n517_), .A2(new_n521_), .A3(new_n510_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT67), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n523_), .A3(new_n515_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(KEYINPUT8), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n523_), .B1(new_n522_), .B2(new_n515_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n516_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(KEYINPUT10), .B(G99gat), .Z(new_n528_));
  NAND2_X1  g327(.A1(new_n528_), .A2(new_n506_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n515_), .A2(KEYINPUT9), .ZN(new_n530_));
  INV_X1    g329(.A(G85gat), .ZN(new_n531_));
  INV_X1    g330(.A(G92gat), .ZN(new_n532_));
  OR3_X1    g331(.A1(new_n531_), .A2(new_n532_), .A3(KEYINPUT9), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n529_), .A2(new_n530_), .A3(new_n510_), .A4(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n501_), .B1(new_n527_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT69), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n534_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n522_), .A2(new_n515_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT67), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(KEYINPUT8), .A3(new_n524_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n538_), .B1(new_n541_), .B2(new_n516_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT69), .B1(new_n542_), .B2(new_n501_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT12), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(new_n542_), .B2(new_n498_), .ZN(new_n545_));
  AND2_X1   g344(.A1(G230gat), .A2(G233gat), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n542_), .B2(new_n498_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n537_), .A2(new_n543_), .A3(new_n545_), .A4(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n527_), .A2(new_n534_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n498_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n542_), .A2(new_n498_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n546_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G120gat), .B(G148gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT5), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G176gat), .B(G204gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n548_), .A2(new_n554_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n559_), .B1(new_n548_), .B2(new_n554_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(G190gat), .B(G218gat), .Z(new_n567_));
  XNOR2_X1  g366(.A(G134gat), .B(G162gat), .ZN(new_n568_));
  OR2_X1    g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n568_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT36), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n527_), .A2(new_n475_), .A3(new_n534_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G232gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT34), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(KEYINPUT35), .ZN(new_n576_));
  INV_X1    g375(.A(new_n477_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n573_), .B(new_n576_), .C1(new_n577_), .C2(new_n542_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(KEYINPUT35), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT70), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n579_), .B1(new_n573_), .B2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n578_), .A2(new_n581_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n572_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  AND2_X1   g383(.A1(new_n573_), .A2(new_n576_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n549_), .A2(new_n477_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT70), .B1(new_n542_), .B2(new_n475_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n585_), .B(new_n586_), .C1(new_n587_), .C2(new_n579_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n578_), .A2(new_n581_), .ZN(new_n589_));
  AOI21_X1  g388(.A(KEYINPUT36), .B1(new_n569_), .B2(new_n570_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT71), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n591_), .B(KEYINPUT72), .Z(new_n592_));
  NAND3_X1  g391(.A1(new_n588_), .A2(new_n589_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n584_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT73), .ZN(new_n595_));
  INV_X1    g394(.A(new_n572_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n594_), .B(KEYINPUT37), .C1(new_n595_), .C2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599_));
  OAI211_X1 g398(.A(new_n584_), .B(new_n593_), .C1(KEYINPUT73), .C2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G127gat), .B(G155gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G183gat), .B(G211gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT17), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n606_), .A2(new_n607_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G231gat), .A2(G233gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n471_), .B(new_n610_), .Z(new_n611_));
  AOI211_X1 g410(.A(new_n608_), .B(new_n609_), .C1(new_n611_), .C2(new_n498_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n498_), .B2(new_n611_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n499_), .A2(new_n500_), .ZN(new_n614_));
  OR2_X1    g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n611_), .A2(new_n614_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(new_n616_), .A3(new_n608_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n613_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n601_), .A2(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n566_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n491_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n304_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(new_n465_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT38), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n454_), .A2(new_n457_), .A3(new_n304_), .A4(new_n240_), .ZN(new_n628_));
  AOI22_X1  g427(.A1(new_n453_), .A2(new_n454_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n628_), .B1(new_n629_), .B2(new_n240_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n584_), .A2(new_n593_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n618_), .A2(new_n631_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n489_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n566_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G1gat), .B1(new_n636_), .B2(new_n304_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n625_), .A2(new_n626_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n627_), .A2(new_n637_), .A3(new_n638_), .ZN(G1324gat));
  OAI21_X1  g438(.A(G8gat), .B1(new_n636_), .B2(new_n457_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT39), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n623_), .A2(new_n397_), .A3(new_n464_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g443(.A(G15gat), .B1(new_n636_), .B2(new_n239_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT41), .ZN(new_n646_));
  NOR3_X1   g445(.A1(new_n622_), .A2(G15gat), .A3(new_n239_), .ZN(new_n647_));
  OR2_X1    g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1326gat));
  OAI21_X1  g447(.A(G22gat), .B1(new_n636_), .B2(new_n454_), .ZN(new_n649_));
  XOR2_X1   g448(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  OR2_X1    g450(.A1(new_n454_), .A2(G22gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n651_), .B1(new_n622_), .B2(new_n652_), .ZN(G1327gat));
  NOR3_X1   g452(.A1(new_n566_), .A2(new_n619_), .A3(new_n594_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n491_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G29gat), .B1(new_n656_), .B2(new_n624_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n566_), .A2(new_n634_), .A3(new_n619_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n598_), .A2(KEYINPUT103), .A3(new_n600_), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT103), .B1(new_n598_), .B2(new_n600_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(KEYINPUT43), .B1(new_n460_), .B2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(KEYINPUT37), .B1(new_n597_), .B2(new_n595_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n631_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n600_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(new_n630_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n659_), .B1(new_n663_), .B2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT104), .B1(new_n672_), .B2(KEYINPUT44), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n674_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n598_), .A2(KEYINPUT103), .A3(new_n600_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n668_), .B1(new_n630_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n458_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n448_), .A2(new_n452_), .ZN(new_n680_));
  OAI211_X1 g479(.A(KEYINPUT32), .B(new_n376_), .C1(new_n385_), .C2(new_n386_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n301_), .A2(new_n681_), .A3(new_n303_), .A4(new_n441_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n438_), .B1(new_n680_), .B2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n239_), .B1(new_n679_), .B2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n669_), .B1(new_n684_), .B2(new_n628_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n658_), .B1(new_n678_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n686_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n673_), .A2(new_n689_), .ZN(new_n690_));
  OAI211_X1 g489(.A(KEYINPUT44), .B(new_n658_), .C1(new_n678_), .C2(new_n685_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n624_), .A2(G29gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n657_), .B1(new_n692_), .B2(new_n693_), .ZN(G1328gat));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n397_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n457_), .A2(KEYINPUT106), .ZN(new_n697_));
  AND2_X1   g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n655_), .A2(G36gat), .A3(new_n698_), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT45), .Z(new_n700_));
  AOI21_X1  g499(.A(new_n457_), .B1(new_n672_), .B2(KEYINPUT44), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n686_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n687_), .B1(new_n686_), .B2(new_n688_), .ZN(new_n703_));
  OAI211_X1 g502(.A(KEYINPUT105), .B(new_n701_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G36gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT105), .B1(new_n690_), .B2(new_n701_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n700_), .B1(new_n705_), .B2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT46), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT46), .B(new_n700_), .C1(new_n705_), .C2(new_n706_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1329gat));
  NAND4_X1  g510(.A1(new_n690_), .A2(G43gat), .A3(new_n240_), .A4(new_n691_), .ZN(new_n712_));
  INV_X1    g511(.A(G43gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n713_), .B1(new_n655_), .B2(new_n239_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g515(.A(G50gat), .B1(new_n656_), .B2(new_n438_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n438_), .A2(G50gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n692_), .B2(new_n718_), .ZN(G1331gat));
  AND3_X1   g518(.A1(new_n633_), .A2(new_n490_), .A3(new_n566_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(G57gat), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n721_), .A2(new_n722_), .A3(new_n304_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n630_), .A2(new_n634_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT107), .Z(new_n725_));
  NOR2_X1   g524(.A1(new_n620_), .A2(new_n565_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n304_), .B1(new_n727_), .B2(KEYINPUT108), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n728_), .B1(KEYINPUT108), .B2(new_n727_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n723_), .B1(new_n729_), .B2(new_n722_), .ZN(G1332gat));
  INV_X1    g529(.A(G64gat), .ZN(new_n731_));
  INV_X1    g530(.A(new_n698_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n720_), .B2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT110), .ZN(new_n734_));
  XNOR2_X1  g533(.A(KEYINPUT109), .B(KEYINPUT48), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n727_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(new_n731_), .A3(new_n732_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n736_), .A2(new_n738_), .ZN(G1333gat));
  INV_X1    g538(.A(G71gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n720_), .B2(new_n240_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT49), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n737_), .A2(new_n740_), .A3(new_n240_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1334gat));
  OAI21_X1  g543(.A(G78gat), .B1(new_n721_), .B2(new_n454_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT50), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n454_), .A2(G78gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n727_), .B2(new_n747_), .ZN(G1335gat));
  NAND3_X1  g547(.A1(new_n566_), .A2(new_n634_), .A3(new_n618_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n663_), .B2(new_n671_), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n750_), .A2(KEYINPUT111), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(KEYINPUT111), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(G85gat), .B1(new_n753_), .B2(new_n304_), .ZN(new_n754_));
  AND4_X1   g553(.A1(new_n566_), .A2(new_n725_), .A3(new_n618_), .A4(new_n631_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n531_), .A3(new_n624_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1336gat));
  OAI21_X1  g556(.A(G92gat), .B1(new_n753_), .B2(new_n698_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n755_), .A2(new_n532_), .A3(new_n397_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(G1337gat));
  NAND3_X1  g559(.A1(new_n755_), .A2(new_n240_), .A3(new_n528_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n239_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(new_n505_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT51), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT51), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n761_), .B(new_n765_), .C1(new_n762_), .C2(new_n505_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1338gat));
  NAND3_X1  g566(.A1(new_n755_), .A2(new_n506_), .A3(new_n438_), .ZN(new_n768_));
  AOI211_X1 g567(.A(KEYINPUT52), .B(new_n506_), .C1(new_n750_), .C2(new_n438_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n750_), .A2(new_n438_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(G106gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n768_), .B1(new_n769_), .B2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT53), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT53), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n768_), .B(new_n775_), .C1(new_n772_), .C2(new_n769_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(G1339gat));
  NAND2_X1  g576(.A1(new_n548_), .A2(KEYINPUT55), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n551_), .A2(new_n544_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT55), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n779_), .A2(new_n780_), .A3(new_n543_), .A4(new_n547_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n778_), .A2(new_n781_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n537_), .A2(new_n543_), .A3(new_n545_), .A4(new_n552_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n546_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT56), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n559_), .A2(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(KEYINPUT112), .A3(new_n787_), .ZN(new_n788_));
  AOI22_X1  g587(.A1(new_n778_), .A2(new_n781_), .B1(new_n546_), .B2(new_n783_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n786_), .B1(new_n789_), .B2(new_n559_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT112), .ZN(new_n791_));
  INV_X1    g590(.A(new_n787_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n791_), .B1(new_n789_), .B2(new_n792_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n788_), .A2(new_n790_), .A3(new_n793_), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n480_), .A2(new_n463_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n472_), .A2(new_n475_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(new_n478_), .A3(new_n463_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n484_), .B1(new_n795_), .B2(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n798_), .B1(new_n484_), .B2(new_n481_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n799_), .A2(new_n561_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n794_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT58), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n794_), .A2(KEYINPUT58), .A3(new_n800_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n803_), .A2(new_n667_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n489_), .A2(new_n560_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n785_), .A2(new_n787_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n790_), .B2(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n799_), .A2(new_n563_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n594_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT57), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(KEYINPUT57), .B(new_n594_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n805_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n618_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n565_), .A2(new_n490_), .A3(new_n601_), .A4(new_n619_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT54), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n815_), .A2(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n397_), .A2(new_n438_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n821_), .A2(new_n624_), .A3(new_n240_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n820_), .A2(KEYINPUT59), .A3(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n818_), .B1(new_n814_), .B2(new_n618_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n822_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n824_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G113gat), .B1(new_n829_), .B2(new_n490_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n820_), .A2(new_n831_), .A3(new_n823_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT113), .B1(new_n826_), .B2(new_n822_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(G113gat), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n835_), .A3(new_n489_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n830_), .A2(new_n836_), .ZN(G1340gat));
  OAI21_X1  g636(.A(G120gat), .B1(new_n829_), .B2(new_n565_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n565_), .A2(KEYINPUT60), .ZN(new_n839_));
  MUX2_X1   g638(.A(new_n839_), .B(KEYINPUT60), .S(G120gat), .Z(new_n840_));
  NAND2_X1  g639(.A1(new_n834_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n841_), .ZN(G1341gat));
  NAND3_X1  g641(.A1(new_n832_), .A2(new_n619_), .A3(new_n833_), .ZN(new_n843_));
  INV_X1    g642(.A(G127gat), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT114), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT114), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n843_), .A2(new_n847_), .A3(new_n844_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n618_), .A2(new_n844_), .ZN(new_n849_));
  AOI22_X1  g648(.A1(new_n846_), .A2(new_n848_), .B1(new_n828_), .B2(new_n849_), .ZN(G1342gat));
  AOI21_X1  g649(.A(G134gat), .B1(new_n834_), .B2(new_n631_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n667_), .A2(G134gat), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT115), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n828_), .B2(new_n853_), .ZN(G1343gat));
  NAND4_X1  g653(.A1(new_n698_), .A2(new_n624_), .A3(new_n438_), .A4(new_n239_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT116), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n815_), .B2(new_n819_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n489_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT117), .B(G141gat), .Z(new_n859_));
  XNOR2_X1  g658(.A(new_n858_), .B(new_n859_), .ZN(G1344gat));
  NAND2_X1  g659(.A1(new_n857_), .A2(new_n566_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(KEYINPUT118), .B(G148gat), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1345gat));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n856_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n812_), .A2(new_n813_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n619_), .B1(new_n867_), .B2(new_n805_), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n619_), .B(new_n866_), .C1(new_n868_), .C2(new_n818_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(KEYINPUT119), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n857_), .A2(new_n871_), .A3(new_n619_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873_));
  AND3_X1   g672(.A1(new_n870_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n865_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n870_), .A2(new_n872_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(KEYINPUT120), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n870_), .A2(new_n872_), .A3(new_n873_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n878_), .A2(new_n864_), .A3(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n876_), .A2(new_n880_), .ZN(G1346gat));
  INV_X1    g680(.A(new_n857_), .ZN(new_n882_));
  INV_X1    g681(.A(G162gat), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n882_), .A2(new_n883_), .A3(new_n662_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n882_), .B2(new_n594_), .ZN(new_n885_));
  OR2_X1    g684(.A1(new_n885_), .A2(KEYINPUT121), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(KEYINPUT121), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n884_), .B1(new_n886_), .B2(new_n887_), .ZN(G1347gat));
  NOR3_X1   g687(.A1(new_n698_), .A2(new_n438_), .A3(new_n305_), .ZN(new_n889_));
  AND2_X1   g688(.A1(new_n820_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n489_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(G169gat), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n891_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n895_));
  OAI211_X1 g694(.A(new_n894_), .B(new_n895_), .C1(new_n353_), .C2(new_n891_), .ZN(G1348gat));
  XOR2_X1   g695(.A(KEYINPUT122), .B(G176gat), .Z(new_n897_));
  NOR2_X1   g696(.A1(KEYINPUT122), .A2(G176gat), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n820_), .A2(new_n889_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n899_), .A2(new_n565_), .ZN(new_n900_));
  MUX2_X1   g699(.A(new_n897_), .B(new_n898_), .S(new_n900_), .Z(G1349gat));
  NOR2_X1   g700(.A1(new_n899_), .A2(new_n618_), .ZN(new_n902_));
  MUX2_X1   g701(.A(G183gat), .B(new_n206_), .S(new_n902_), .Z(G1350gat));
  NAND3_X1  g702(.A1(new_n890_), .A2(new_n207_), .A3(new_n631_), .ZN(new_n904_));
  OAI21_X1  g703(.A(G190gat), .B1(new_n899_), .B2(new_n601_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1351gat));
  AOI21_X1  g705(.A(new_n634_), .B1(KEYINPUT124), .B2(new_n332_), .ZN(new_n907_));
  NOR4_X1   g706(.A1(new_n698_), .A2(new_n624_), .A3(new_n454_), .A4(new_n240_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n820_), .A2(new_n908_), .ZN(new_n909_));
  AND2_X1   g708(.A1(new_n909_), .A2(KEYINPUT123), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n909_), .A2(KEYINPUT123), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n907_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n332_), .A2(KEYINPUT124), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n913_), .B(KEYINPUT125), .Z(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n912_), .A2(new_n915_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n907_), .B(new_n914_), .C1(new_n910_), .C2(new_n911_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1352gat));
  NOR2_X1   g717(.A1(new_n910_), .A2(new_n911_), .ZN(new_n919_));
  OAI21_X1  g718(.A(G204gat), .B1(new_n919_), .B2(new_n565_), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n334_), .B(new_n566_), .C1(new_n910_), .C2(new_n911_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(G1353gat));
  NOR3_X1   g721(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n923_));
  AOI211_X1 g722(.A(new_n923_), .B(new_n618_), .C1(KEYINPUT63), .C2(G211gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n924_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n925_));
  OAI21_X1  g724(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n925_), .A2(new_n927_), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n926_), .B(new_n924_), .C1(new_n910_), .C2(new_n911_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1354gat));
  INV_X1    g729(.A(new_n911_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n909_), .A2(KEYINPUT123), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n601_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n631_), .A2(new_n308_), .ZN(new_n934_));
  OAI22_X1  g733(.A1(new_n933_), .A2(new_n308_), .B1(new_n919_), .B2(new_n934_), .ZN(G1355gat));
endmodule


