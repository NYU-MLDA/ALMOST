//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n951_, new_n952_, new_n953_, new_n955_,
    new_n956_, new_n958_, new_n959_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n966_, new_n967_, new_n968_, new_n969_;
  INV_X1    g000(.A(KEYINPUT82), .ZN(new_n202_));
  INV_X1    g001(.A(G183gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT25), .ZN(new_n204_));
  OR2_X1    g003(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  OR2_X1    g006(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n208_));
  NAND2_X1  g007(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n203_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT81), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n204_), .B(new_n207_), .C1(new_n210_), .C2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(new_n209_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(KEYINPUT80), .A2(KEYINPUT25), .ZN(new_n214_));
  OAI211_X1 g013(.A(new_n211_), .B(G183gat), .C1(new_n213_), .C2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n202_), .B1(new_n212_), .B2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(G183gat), .B1(new_n213_), .B2(new_n214_), .ZN(new_n218_));
  AOI22_X1  g017(.A1(new_n218_), .A2(KEYINPUT81), .B1(new_n205_), .B2(new_n206_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n219_), .A2(KEYINPUT82), .A3(new_n204_), .A4(new_n215_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n221_));
  AND3_X1   g020(.A1(KEYINPUT83), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT83), .B1(G183gat), .B2(G190gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n227_), .A2(KEYINPUT24), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n227_), .A2(KEYINPUT24), .A3(new_n230_), .ZN(new_n231_));
  AND4_X1   g030(.A1(new_n224_), .A2(new_n228_), .A3(new_n229_), .A4(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n217_), .A2(new_n220_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT84), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n234_), .B1(new_n225_), .B2(KEYINPUT22), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT22), .B(G169gat), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n226_), .B(new_n235_), .C1(new_n236_), .C2(new_n234_), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT23), .B1(new_n222_), .B2(new_n223_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n221_), .A2(G183gat), .A3(G190gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT85), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT85), .ZN(new_n244_));
  AOI211_X1 g043(.A(new_n244_), .B(new_n241_), .C1(new_n238_), .C2(new_n239_), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n230_), .B(new_n237_), .C1(new_n243_), .C2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n233_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT30), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n233_), .A2(new_n246_), .A3(KEYINPUT30), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT86), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT86), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n249_), .A2(new_n253_), .A3(new_n250_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G71gat), .B(G99gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G227gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G15gat), .B(G43gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n257_), .B(new_n258_), .Z(new_n259_));
  NAND3_X1  g058(.A1(new_n252_), .A2(new_n254_), .A3(new_n259_), .ZN(new_n260_));
  OR3_X1    g059(.A1(new_n251_), .A2(KEYINPUT86), .A3(new_n259_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT87), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT31), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT31), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .A4(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G127gat), .B(G134gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G113gat), .B(G120gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n264_), .A2(new_n270_), .A3(new_n266_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G64gat), .B(G92gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(G8gat), .B(G36gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT102), .B(KEYINPUT18), .ZN(new_n278_));
  XOR2_X1   g077(.A(new_n277_), .B(new_n278_), .Z(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G226gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT19), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n282_), .B(KEYINPUT97), .Z(new_n283_));
  INV_X1    g082(.A(KEYINPUT98), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n205_), .A2(new_n284_), .A3(new_n206_), .ZN(new_n285_));
  AND2_X1   g084(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT98), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT25), .B(G183gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n285_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n231_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT99), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n240_), .A2(new_n228_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT99), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n290_), .A2(new_n295_), .A3(new_n231_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n294_), .A3(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT100), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n224_), .A2(new_n242_), .A3(new_n229_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n236_), .A2(new_n226_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n230_), .B(KEYINPUT101), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n300_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT100), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n292_), .A2(new_n303_), .A3(new_n294_), .A4(new_n296_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n298_), .A2(new_n302_), .A3(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G211gat), .A2(G218gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G211gat), .A2(G218gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n307_), .A2(KEYINPUT93), .A3(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT93), .ZN(new_n310_));
  INV_X1    g109(.A(new_n308_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n310_), .B1(new_n311_), .B2(new_n306_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(KEYINPUT92), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G197gat), .B(G204gat), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT21), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n313_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n315_), .A2(new_n316_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n314_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n313_), .B(new_n317_), .C1(KEYINPUT92), .C2(new_n319_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n305_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n233_), .A2(new_n323_), .A3(new_n246_), .ZN(new_n326_));
  AND2_X1   g125(.A1(new_n326_), .A2(KEYINPUT20), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n283_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT20), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n247_), .B2(new_n324_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n298_), .A2(new_n323_), .A3(new_n302_), .A4(new_n304_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n282_), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n280_), .B1(new_n328_), .B2(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n326_), .A2(KEYINPUT20), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n336_), .B1(new_n324_), .B2(new_n305_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n335_), .B(new_n279_), .C1(new_n337_), .C2(new_n283_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(KEYINPUT103), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT27), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT103), .ZN(new_n341_));
  OAI211_X1 g140(.A(new_n341_), .B(new_n280_), .C1(new_n328_), .C2(new_n333_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT107), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n290_), .A2(new_n295_), .A3(new_n231_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n295_), .B1(new_n290_), .B2(new_n231_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n345_), .A2(new_n346_), .A3(new_n293_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n302_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n344_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n297_), .A2(KEYINPUT107), .A3(new_n302_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n323_), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n351_), .A2(new_n330_), .ZN(new_n352_));
  AOI22_X1  g151(.A1(new_n337_), .A2(new_n283_), .B1(new_n352_), .B2(new_n282_), .ZN(new_n353_));
  OAI211_X1 g152(.A(KEYINPUT27), .B(new_n338_), .C1(new_n353_), .C2(new_n279_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n343_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT4), .ZN(new_n358_));
  AND3_X1   g157(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n359_));
  AOI21_X1  g158(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT1), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT88), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT1), .ZN(new_n365_));
  NAND3_X1  g164(.A1(KEYINPUT88), .A2(G155gat), .A3(G162gat), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  OR2_X1    g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n361_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  XOR2_X1   g168(.A(G141gat), .B(G148gat), .Z(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n368_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT89), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT89), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n374_), .B(new_n368_), .C1(new_n359_), .C2(new_n360_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT2), .ZN(new_n376_));
  INV_X1    g175(.A(G141gat), .ZN(new_n377_));
  INV_X1    g176(.A(G148gat), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n376_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT3), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n380_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n379_), .A2(new_n381_), .A3(new_n382_), .A4(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n373_), .A2(new_n375_), .A3(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n371_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n271_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n371_), .A2(new_n385_), .A3(new_n270_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n387_), .A2(KEYINPUT104), .A3(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT104), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n386_), .A2(new_n390_), .A3(new_n271_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n358_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n387_), .A2(KEYINPUT4), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n357_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G57gat), .B(G85gat), .Z(new_n395_));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT105), .B(KEYINPUT0), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n389_), .A2(new_n391_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(new_n356_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n394_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n400_), .B1(new_n394_), .B2(new_n402_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n323_), .B1(KEYINPUT29), .B2(new_n386_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(G228gat), .A2(G233gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT91), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT94), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n408_), .B1(new_n323_), .B2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n406_), .B(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G78gat), .B(G106gat), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n406_), .A2(new_n410_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n406_), .A2(new_n410_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n415_), .A2(new_n416_), .A3(new_n412_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n414_), .A2(KEYINPUT95), .A3(new_n417_), .ZN(new_n418_));
  OR3_X1    g217(.A1(new_n411_), .A2(KEYINPUT95), .A3(new_n413_), .ZN(new_n419_));
  OR3_X1    g218(.A1(new_n386_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT28), .B1(new_n386_), .B2(KEYINPUT29), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G22gat), .B(G50gat), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n422_), .A2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n422_), .A2(new_n424_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(KEYINPUT90), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n430_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n418_), .A2(new_n419_), .A3(new_n429_), .A4(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT96), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n417_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n414_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n411_), .A2(new_n433_), .A3(new_n413_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n435_), .A2(new_n428_), .A3(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n432_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n274_), .A2(new_n355_), .A3(new_n405_), .A4(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n279_), .A2(KEYINPUT32), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n335_), .B(new_n441_), .C1(new_n337_), .C2(new_n283_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n442_), .B1(new_n353_), .B2(new_n441_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT108), .B1(new_n443_), .B2(new_n405_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n394_), .A2(new_n402_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(new_n399_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n394_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT108), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n325_), .A2(new_n327_), .A3(new_n283_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n332_), .B1(new_n351_), .B2(new_n330_), .ZN(new_n451_));
  OAI211_X1 g250(.A(KEYINPUT32), .B(new_n279_), .C1(new_n450_), .C2(new_n451_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n448_), .A2(new_n449_), .A3(new_n442_), .A4(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n339_), .A2(new_n342_), .ZN(new_n454_));
  OR3_X1    g253(.A1(new_n392_), .A2(new_n357_), .A3(new_n393_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT106), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n401_), .B(new_n456_), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n400_), .B(new_n455_), .C1(new_n457_), .C2(new_n356_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT33), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n404_), .A2(new_n459_), .ZN(new_n460_));
  AOI211_X1 g259(.A(KEYINPUT33), .B(new_n400_), .C1(new_n394_), .C2(new_n402_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n458_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n444_), .B(new_n453_), .C1(new_n454_), .C2(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n448_), .B1(new_n432_), .B2(new_n437_), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n463_), .A2(new_n439_), .B1(new_n355_), .B2(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n440_), .B1(new_n465_), .B2(new_n274_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G230gat), .A2(G233gat), .ZN(new_n467_));
  XOR2_X1   g266(.A(new_n467_), .B(KEYINPUT64), .Z(new_n468_));
  OR3_X1    g267(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G99gat), .A2(G106gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n469_), .A2(new_n472_), .A3(new_n473_), .A4(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G85gat), .ZN(new_n476_));
  INV_X1    g275(.A(G92gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G85gat), .A2(G92gat), .ZN(new_n479_));
  AND3_X1   g278(.A1(new_n478_), .A2(KEYINPUT68), .A3(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n475_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT8), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT8), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n482_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT67), .ZN(new_n486_));
  INV_X1    g285(.A(G99gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT10), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT10), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(G99gat), .ZN(new_n490_));
  AOI21_X1  g289(.A(G106gat), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n472_), .A2(new_n473_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT65), .ZN(new_n494_));
  AND3_X1   g293(.A1(new_n479_), .A2(new_n494_), .A3(KEYINPUT9), .ZN(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT9), .B1(new_n479_), .B2(new_n494_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n479_), .A2(KEYINPUT66), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n495_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT9), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n479_), .A2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n500_), .B1(KEYINPUT66), .B2(new_n478_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n486_), .B(new_n493_), .C1(new_n498_), .C2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n479_), .A2(new_n494_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n499_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n479_), .A2(KEYINPUT66), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n479_), .A2(new_n494_), .A3(KEYINPUT9), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n505_), .A2(new_n506_), .A3(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n478_), .A2(KEYINPUT66), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n509_), .B1(new_n499_), .B2(new_n479_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n486_), .B1(new_n511_), .B2(new_n493_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n485_), .B1(new_n503_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G57gat), .A2(G64gat), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(G57gat), .A2(G64gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT69), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(G57gat), .A2(G64gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT69), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n518_), .A2(new_n519_), .A3(new_n514_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(KEYINPUT11), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT11), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n517_), .A2(new_n520_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G71gat), .B(G78gat), .Z(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n523_), .B1(new_n517_), .B2(new_n520_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(new_n526_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n513_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n529_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n533_), .B(new_n485_), .C1(new_n512_), .C2(new_n503_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n534_), .A3(KEYINPUT12), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT12), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n513_), .A2(new_n536_), .A3(new_n531_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n468_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT70), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n532_), .A2(new_n534_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(new_n468_), .ZN(new_n542_));
  XOR2_X1   g341(.A(G176gat), .B(G204gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(G120gat), .B(G148gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n540_), .A2(KEYINPUT72), .A3(new_n542_), .A4(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n535_), .A2(new_n537_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n468_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n539_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n551_));
  AOI211_X1 g350(.A(KEYINPUT70), .B(new_n468_), .C1(new_n535_), .C2(new_n537_), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n542_), .B(new_n547_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT72), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n548_), .A2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n540_), .A2(new_n542_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n547_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n556_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n562_));
  AOI21_X1  g361(.A(new_n562_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT15), .ZN(new_n565_));
  XNOR2_X1  g364(.A(G43gat), .B(G50gat), .ZN(new_n566_));
  INV_X1    g365(.A(G36gat), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n567_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(KEYINPUT75), .B(G29gat), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n570_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n565_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G15gat), .B(G22gat), .ZN(new_n575_));
  INV_X1    g374(.A(G1gat), .ZN(new_n576_));
  INV_X1    g375(.A(G8gat), .ZN(new_n577_));
  OAI21_X1  g376(.A(KEYINPUT14), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G1gat), .B(G8gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n566_), .B(new_n567_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n570_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(KEYINPUT15), .A3(new_n571_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n574_), .A2(new_n581_), .A3(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(G229gat), .A2(G233gat), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n571_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n581_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n586_), .A2(new_n587_), .A3(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n581_), .A2(new_n584_), .A3(new_n571_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n587_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n591_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT78), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT78), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n595_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT79), .B(G113gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n601_), .B(G141gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G169gat), .B(G197gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n602_), .B(new_n603_), .Z(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n604_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n597_), .A2(new_n599_), .A3(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n564_), .A2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n466_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT77), .ZN(new_n612_));
  NAND2_X1  g411(.A1(G232gat), .A2(G233gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT34), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n614_), .A2(KEYINPUT35), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n511_), .A2(new_n493_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT67), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n617_), .A2(new_n502_), .B1(new_n484_), .B2(new_n482_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n615_), .B1(new_n618_), .B2(new_n588_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n513_), .A2(new_n585_), .A3(new_n574_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n614_), .A2(KEYINPUT35), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT74), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n621_), .A2(KEYINPUT76), .A3(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G190gat), .B(G218gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G134gat), .B(G162gat), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n625_), .B(new_n626_), .Z(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT36), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(KEYINPUT76), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n623_), .A2(KEYINPUT76), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n619_), .A2(new_n629_), .A3(new_n630_), .A4(new_n620_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n624_), .A2(new_n628_), .A3(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n627_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n633_), .A2(KEYINPUT36), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n635_), .B1(new_n624_), .B2(new_n631_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n612_), .B1(new_n632_), .B2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT37), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n624_), .A2(new_n628_), .A3(new_n631_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT77), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n637_), .A2(new_n638_), .A3(new_n640_), .ZN(new_n641_));
  OAI21_X1  g440(.A(KEYINPUT37), .B1(new_n632_), .B2(new_n636_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(G231gat), .A2(G233gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n581_), .B(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(new_n533_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(G127gat), .B(G155gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(G211gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT16), .B(G183gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n647_), .B1(KEYINPUT17), .B2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(KEYINPUT17), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n647_), .A2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n644_), .A2(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n611_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n576_), .A3(new_n448_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT38), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT109), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n637_), .A2(new_n660_), .A3(new_n640_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n637_), .B2(new_n640_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(new_n655_), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n611_), .A2(new_n664_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n665_), .A2(new_n448_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n659_), .B1(new_n576_), .B2(new_n666_), .ZN(G1324gat));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT111), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n343_), .A2(new_n354_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n466_), .A2(new_n610_), .A3(new_n664_), .A4(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(G8gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n669_), .B1(new_n672_), .B2(KEYINPUT39), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n671_), .A2(KEYINPUT111), .A3(new_n674_), .A4(G8gat), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  AOI211_X1 g475(.A(KEYINPUT110), .B(new_n674_), .C1(new_n671_), .C2(G8gat), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT110), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n672_), .B2(KEYINPUT39), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n676_), .A2(new_n677_), .A3(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n657_), .A2(new_n577_), .A3(new_n670_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n668_), .B1(new_n680_), .B2(new_n682_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n679_), .A2(new_n677_), .ZN(new_n684_));
  OAI211_X1 g483(.A(KEYINPUT40), .B(new_n681_), .C1(new_n684_), .C2(new_n676_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n683_), .A2(new_n685_), .ZN(G1325gat));
  INV_X1    g485(.A(G15gat), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n687_), .B1(new_n665_), .B2(new_n274_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT41), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n657_), .A2(new_n687_), .A3(new_n274_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT112), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1326gat));
  INV_X1    g491(.A(G22gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n693_), .B1(new_n665_), .B2(new_n438_), .ZN(new_n694_));
  XOR2_X1   g493(.A(new_n694_), .B(KEYINPUT42), .Z(new_n695_));
  NAND3_X1  g494(.A1(new_n657_), .A2(new_n693_), .A3(new_n438_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(G1327gat));
  INV_X1    g496(.A(new_n663_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n655_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n611_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(G29gat), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(new_n448_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT116), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n655_), .B(new_n608_), .C1(new_n561_), .C2(new_n563_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT113), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  AOI22_X1  g506(.A1(new_n548_), .A2(new_n555_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n560_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n709_), .B1(new_n708_), .B2(new_n562_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n710_), .A2(KEYINPUT113), .A3(new_n655_), .A4(new_n608_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n707_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n713_));
  XNOR2_X1  g512(.A(new_n643_), .B(KEYINPUT114), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n713_), .B1(new_n466_), .B2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n644_), .A2(new_n713_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n274_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n444_), .A2(new_n453_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n339_), .A2(new_n342_), .ZN(new_n720_));
  OAI211_X1 g519(.A(new_n720_), .B(new_n458_), .C1(new_n460_), .C2(new_n461_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n438_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n464_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n723_), .A2(new_n670_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n718_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n717_), .B1(new_n725_), .B2(new_n440_), .ZN(new_n726_));
  OAI211_X1 g525(.A(KEYINPUT44), .B(new_n712_), .C1(new_n716_), .C2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(KEYINPUT115), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n466_), .A2(new_n713_), .A3(new_n644_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n714_), .B1(new_n725_), .B2(new_n440_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n729_), .B1(new_n730_), .B2(new_n713_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT115), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n731_), .A2(new_n732_), .A3(KEYINPUT44), .A4(new_n712_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n728_), .A2(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n712_), .B1(new_n716_), .B2(new_n726_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n405_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n737_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n704_), .B1(new_n738_), .B2(G29gat), .ZN(new_n739_));
  AOI211_X1 g538(.A(KEYINPUT116), .B(new_n702_), .C1(new_n734_), .C2(new_n737_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n703_), .B1(new_n739_), .B2(new_n740_), .ZN(G1328gat));
  NAND3_X1  g540(.A1(new_n611_), .A2(new_n567_), .A3(new_n700_), .ZN(new_n742_));
  XNOR2_X1  g541(.A(new_n670_), .B(KEYINPUT117), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  OR3_X1    g543(.A1(new_n742_), .A2(KEYINPUT45), .A3(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT45), .B1(new_n742_), .B2(new_n744_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n735_), .A2(new_n736_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(new_n670_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n728_), .B2(new_n733_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT46), .B(new_n747_), .C1(new_n750_), .C2(new_n567_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT46), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n355_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n567_), .B1(new_n734_), .B2(new_n753_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n745_), .A2(new_n746_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n752_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n751_), .A2(new_n756_), .ZN(G1329gat));
  INV_X1    g556(.A(G43gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n734_), .A2(new_n274_), .A3(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n701_), .A2(new_n274_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT47), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n760_), .A2(new_n765_), .A3(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1330gat));
  AOI21_X1  g566(.A(new_n439_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n734_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT118), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n734_), .A2(KEYINPUT118), .A3(new_n768_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(G50gat), .A3(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(G50gat), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n701_), .A2(new_n774_), .A3(new_n438_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n773_), .A2(new_n775_), .ZN(G1331gat));
  NOR2_X1   g575(.A1(new_n710_), .A2(new_n608_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n466_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n656_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT119), .Z(new_n780_));
  AOI21_X1  g579(.A(G57gat), .B1(new_n780_), .B2(new_n448_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n778_), .A2(new_n664_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n782_), .A2(new_n448_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n781_), .B1(G57gat), .B2(new_n783_), .ZN(G1332gat));
  NOR2_X1   g583(.A1(new_n744_), .A2(G64gat), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT120), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n780_), .A2(new_n786_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n782_), .A2(new_n743_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(G64gat), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n789_), .A2(KEYINPUT48), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(KEYINPUT48), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n787_), .B1(new_n790_), .B2(new_n791_), .ZN(G1333gat));
  INV_X1    g591(.A(G71gat), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n780_), .A2(new_n793_), .A3(new_n274_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n782_), .A2(new_n274_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(G71gat), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n796_), .A2(KEYINPUT49), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n796_), .A2(KEYINPUT49), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(G1334gat));
  INV_X1    g598(.A(G78gat), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n780_), .A2(new_n800_), .A3(new_n438_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n782_), .A2(new_n438_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(G78gat), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n803_), .A2(KEYINPUT50), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n803_), .A2(KEYINPUT50), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n801_), .B1(new_n804_), .B2(new_n805_), .ZN(G1335gat));
  OAI211_X1 g605(.A(new_n655_), .B(new_n777_), .C1(new_n716_), .C2(new_n726_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n807_), .A2(new_n476_), .A3(new_n405_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n778_), .A2(new_n700_), .ZN(new_n809_));
  AOI21_X1  g608(.A(G85gat), .B1(new_n809_), .B2(new_n448_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n808_), .A2(new_n810_), .ZN(G1336gat));
  NOR3_X1   g610(.A1(new_n807_), .A2(new_n477_), .A3(new_n744_), .ZN(new_n812_));
  AOI21_X1  g611(.A(G92gat), .B1(new_n809_), .B2(new_n670_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(G1337gat));
  OAI21_X1  g613(.A(G99gat), .B1(new_n807_), .B2(new_n718_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT51), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n718_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n809_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n815_), .A2(new_n817_), .A3(new_n819_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n816_), .A2(KEYINPUT51), .ZN(new_n821_));
  XOR2_X1   g620(.A(new_n820_), .B(new_n821_), .Z(G1338gat));
  INV_X1    g621(.A(G106gat), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n809_), .A2(new_n823_), .A3(new_n438_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n825_), .B(G106gat), .C1(new_n807_), .C2(new_n439_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n731_), .A2(new_n655_), .A3(new_n438_), .A4(new_n777_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n825_), .B1(new_n828_), .B2(G106gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n824_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT53), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT53), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n832_), .B(new_n824_), .C1(new_n827_), .C2(new_n829_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1339gat));
  NAND3_X1  g633(.A1(new_n710_), .A2(new_n656_), .A3(new_n609_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n835_), .B(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT122), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n586_), .A2(new_n594_), .A3(new_n590_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n593_), .A2(new_n587_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n839_), .A2(new_n840_), .A3(new_n604_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n607_), .A2(new_n838_), .A3(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n838_), .B1(new_n607_), .B2(new_n841_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n844_), .B1(new_n555_), .B2(new_n548_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n538_), .A2(KEYINPUT55), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n847_), .B(new_n848_), .C1(new_n550_), .C2(new_n549_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n849_), .A2(KEYINPUT56), .A3(new_n558_), .ZN(new_n850_));
  AOI21_X1  g649(.A(KEYINPUT56), .B1(new_n849_), .B2(new_n558_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n845_), .B1(new_n850_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(new_n845_), .B(KEYINPUT58), .C1(new_n850_), .C2(new_n851_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n644_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT123), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n849_), .A2(new_n558_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT56), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n849_), .A2(KEYINPUT56), .A3(new_n558_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n609_), .B1(new_n548_), .B2(new_n555_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n708_), .A2(new_n844_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT57), .B(new_n698_), .C1(new_n865_), .C2(new_n866_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n854_), .A2(KEYINPUT123), .A3(new_n644_), .A4(new_n855_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869_));
  INV_X1    g668(.A(new_n708_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n844_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n863_), .A2(new_n864_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n869_), .B1(new_n872_), .B2(new_n663_), .ZN(new_n873_));
  NAND4_X1  g672(.A1(new_n858_), .A2(new_n867_), .A3(new_n868_), .A4(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n837_), .B1(new_n874_), .B2(new_n655_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n355_), .A2(new_n448_), .A3(new_n439_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n718_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n875_), .A2(new_n878_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G113gat), .B1(new_n879_), .B2(new_n608_), .ZN(new_n880_));
  OAI21_X1  g679(.A(KEYINPUT59), .B1(new_n875_), .B2(new_n878_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n867_), .A2(new_n873_), .A3(new_n856_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n655_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n837_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT59), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n885_), .A2(new_n886_), .A3(new_n877_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n881_), .A2(new_n608_), .A3(new_n887_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n880_), .B1(new_n888_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g688(.A(G120gat), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n890_), .B1(new_n710_), .B2(KEYINPUT60), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n879_), .B(new_n891_), .C1(KEYINPUT60), .C2(new_n890_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n881_), .A2(new_n564_), .A3(new_n887_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n890_), .ZN(G1341gat));
  AOI21_X1  g693(.A(G127gat), .B1(new_n879_), .B2(new_n699_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT124), .ZN(new_n896_));
  OAI21_X1  g695(.A(G127gat), .B1(new_n655_), .B2(new_n896_), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n881_), .A2(new_n887_), .A3(new_n897_), .ZN(new_n898_));
  INV_X1    g697(.A(G127gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(KEYINPUT124), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n895_), .B1(new_n898_), .B2(new_n900_), .ZN(G1342gat));
  AOI21_X1  g700(.A(G134gat), .B1(new_n879_), .B2(new_n663_), .ZN(new_n902_));
  AND3_X1   g701(.A1(new_n881_), .A2(G134gat), .A3(new_n887_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(new_n644_), .ZN(G1343gat));
  NOR3_X1   g703(.A1(new_n875_), .A2(new_n439_), .A3(new_n274_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n743_), .A2(new_n405_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n905_), .A2(new_n608_), .A3(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G141gat), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n905_), .A2(new_n377_), .A3(new_n608_), .A4(new_n906_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1344gat));
  NAND3_X1  g709(.A1(new_n905_), .A2(new_n564_), .A3(new_n906_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(G148gat), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n905_), .A2(new_n378_), .A3(new_n564_), .A4(new_n906_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1345gat));
  NAND2_X1  g713(.A1(new_n874_), .A2(new_n655_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n274_), .B1(new_n915_), .B2(new_n884_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n916_), .A2(new_n699_), .A3(new_n438_), .A4(new_n906_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT61), .B(G155gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n917_), .B(new_n918_), .ZN(G1346gat));
  INV_X1    g718(.A(G162gat), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n905_), .A2(new_n663_), .A3(new_n906_), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n916_), .A2(new_n438_), .A3(new_n906_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n714_), .A2(new_n920_), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n920_), .A2(new_n921_), .B1(new_n922_), .B2(new_n923_), .ZN(G1347gat));
  INV_X1    g723(.A(KEYINPUT62), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n743_), .A2(new_n405_), .A3(new_n274_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n926_), .ZN(new_n927_));
  NAND4_X1  g726(.A1(new_n885_), .A2(new_n608_), .A3(new_n439_), .A4(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n925_), .B1(new_n929_), .B2(new_n225_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n236_), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n928_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n930_), .A2(new_n931_), .A3(new_n932_), .ZN(G1348gat));
  AOI21_X1  g732(.A(new_n837_), .B1(new_n655_), .B2(new_n882_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n934_), .A2(new_n438_), .A3(new_n926_), .ZN(new_n935_));
  AOI21_X1  g734(.A(G176gat), .B1(new_n935_), .B2(new_n564_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n927_), .A2(new_n564_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n915_), .A2(new_n884_), .ZN(new_n938_));
  INV_X1    g737(.A(KEYINPUT125), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n938_), .A2(new_n939_), .A3(new_n439_), .ZN(new_n940_));
  OAI21_X1  g739(.A(KEYINPUT125), .B1(new_n875_), .B2(new_n438_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n937_), .B1(new_n940_), .B2(new_n941_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n936_), .B1(new_n942_), .B2(G176gat), .ZN(G1349gat));
  NOR2_X1   g742(.A1(new_n655_), .A2(new_n289_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n935_), .A2(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n926_), .A2(new_n655_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n939_), .B1(new_n938_), .B2(new_n439_), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n875_), .A2(KEYINPUT125), .A3(new_n438_), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n946_), .B1(new_n947_), .B2(new_n948_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n945_), .B1(new_n949_), .B2(new_n203_), .ZN(G1350gat));
  NAND4_X1  g749(.A1(new_n935_), .A2(new_n663_), .A3(new_n288_), .A4(new_n285_), .ZN(new_n951_));
  AND2_X1   g750(.A1(new_n935_), .A2(new_n644_), .ZN(new_n952_));
  INV_X1    g751(.A(G190gat), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n951_), .B1(new_n952_), .B2(new_n953_), .ZN(G1351gat));
  NOR2_X1   g753(.A1(new_n744_), .A2(new_n723_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n916_), .A2(new_n608_), .A3(new_n955_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g756(.A1(new_n916_), .A2(new_n564_), .A3(new_n955_), .ZN(new_n958_));
  XOR2_X1   g757(.A(KEYINPUT126), .B(G204gat), .Z(new_n959_));
  XNOR2_X1  g758(.A(new_n958_), .B(new_n959_), .ZN(G1353gat));
  NAND2_X1  g759(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n961_));
  NAND4_X1  g760(.A1(new_n916_), .A2(new_n699_), .A3(new_n955_), .A4(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n963_));
  XOR2_X1   g762(.A(new_n963_), .B(KEYINPUT127), .Z(new_n964_));
  XNOR2_X1  g763(.A(new_n962_), .B(new_n964_), .ZN(G1354gat));
  NOR4_X1   g764(.A1(new_n875_), .A2(new_n723_), .A3(new_n274_), .A4(new_n744_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n966_), .A2(new_n663_), .ZN(new_n967_));
  INV_X1    g766(.A(G218gat), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n643_), .A2(new_n968_), .ZN(new_n969_));
  AOI22_X1  g768(.A1(new_n967_), .A2(new_n968_), .B1(new_n966_), .B2(new_n969_), .ZN(G1355gat));
endmodule


