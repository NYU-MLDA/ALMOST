//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n848_, new_n849_, new_n850_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_;
  INV_X1    g000(.A(KEYINPUT105), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G190gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT73), .ZN(new_n204_));
  XOR2_X1   g003(.A(G134gat), .B(G162gat), .Z(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT36), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT71), .B(KEYINPUT34), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G232gat), .A2(G233gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n209_), .B(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT72), .B(KEYINPUT35), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n214_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n218_), .B(KEYINPUT65), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n220_), .B1(new_n217_), .B2(KEYINPUT9), .ZN(new_n221_));
  AND2_X1   g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G99gat), .A2(G106gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT6), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT10), .B(G99gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n224_), .B1(G106gat), .B2(new_n225_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n222_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT7), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT66), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(new_n224_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n224_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT66), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n217_), .A2(new_n220_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT8), .ZN(new_n240_));
  INV_X1    g039(.A(new_n236_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n241_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n240_), .B1(new_n242_), .B2(KEYINPUT67), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n239_), .A2(new_n243_), .ZN(new_n244_));
  OAI211_X1 g043(.A(new_n240_), .B(new_n236_), .C1(new_n233_), .C2(new_n230_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n227_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G29gat), .B(G36gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G43gat), .B(G50gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT74), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n251_), .B1(new_n211_), .B2(new_n212_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n249_), .B(KEYINPUT15), .Z(new_n254_));
  NOR2_X1   g053(.A1(new_n246_), .A2(new_n254_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n213_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n207_), .A2(KEYINPUT36), .ZN(new_n257_));
  OR2_X1    g056(.A1(new_n246_), .A2(new_n254_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n213_), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n258_), .A2(new_n259_), .A3(new_n250_), .A4(new_n252_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n256_), .A2(new_n257_), .A3(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n257_), .B1(new_n256_), .B2(new_n260_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n208_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT75), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n261_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT37), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n264_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G57gat), .B(G64gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT11), .ZN(new_n270_));
  XOR2_X1   g069(.A(G71gat), .B(G78gat), .Z(new_n271_));
  OR2_X1    g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n269_), .A2(KEYINPUT11), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n270_), .A2(new_n271_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n272_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G231gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT76), .B(G15gat), .ZN(new_n279_));
  INV_X1    g078(.A(G22gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(G1gat), .ZN(new_n282_));
  INV_X1    g081(.A(G8gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT14), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G1gat), .B(G8gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT77), .ZN(new_n287_));
  OR2_X1    g086(.A1(new_n285_), .A2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n285_), .A2(new_n287_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n278_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G127gat), .B(G155gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT16), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G183gat), .B(G211gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT17), .ZN(new_n296_));
  INV_X1    g095(.A(new_n290_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(new_n277_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n291_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT17), .ZN(new_n300_));
  AOI211_X1 g099(.A(new_n300_), .B(new_n295_), .C1(new_n291_), .C2(new_n298_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n299_), .B1(new_n301_), .B2(KEYINPUT78), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n299_), .A2(KEYINPUT78), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n304_), .A2(KEYINPUT79), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(KEYINPUT79), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n268_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT70), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT13), .ZN(new_n310_));
  NOR2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(KEYINPUT70), .A2(KEYINPUT13), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XOR2_X1   g112(.A(G120gat), .B(G148gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(G176gat), .B(G204gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n316_), .B(new_n317_), .Z(new_n318_));
  XNOR2_X1  g117(.A(new_n246_), .B(new_n275_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n275_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT12), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n235_), .A2(KEYINPUT67), .A3(new_n236_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT8), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n242_), .A2(KEYINPUT67), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n245_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n227_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n275_), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT68), .B1(new_n328_), .B2(KEYINPUT12), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT68), .ZN(new_n330_));
  OAI211_X1 g129(.A(new_n330_), .B(new_n321_), .C1(new_n246_), .C2(new_n275_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n319_), .A2(new_n322_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G230gat), .A2(G233gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n333_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n319_), .A2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n318_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n336_), .A3(new_n318_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n313_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n339_), .ZN(new_n341_));
  NOR3_X1   g140(.A1(new_n341_), .A2(new_n337_), .A3(new_n311_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n308_), .A2(new_n343_), .ZN(new_n344_));
  OR3_X1    g143(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n345_));
  INV_X1    g144(.A(G169gat), .ZN(new_n346_));
  INV_X1    g145(.A(G176gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n345_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G183gat), .A2(G190gat), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT23), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n350_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT25), .B(G183gat), .ZN(new_n357_));
  INV_X1    g156(.A(G190gat), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT26), .B1(new_n358_), .B2(KEYINPUT80), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n358_), .A2(KEYINPUT26), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n357_), .B(new_n359_), .C1(new_n360_), .C2(KEYINPUT80), .ZN(new_n361_));
  INV_X1    g160(.A(G183gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n358_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n353_), .A2(new_n354_), .A3(new_n363_), .ZN(new_n364_));
  OAI21_X1  g163(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n356_), .A2(new_n361_), .B1(new_n364_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G227gat), .A2(G233gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G71gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(G99gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n369_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G15gat), .B(G43gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT81), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT30), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n373_), .B(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT82), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G127gat), .B(G134gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G113gat), .B(G120gat), .ZN(new_n381_));
  OR2_X1    g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n381_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(new_n384_), .B(KEYINPUT31), .Z(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n379_), .A2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n385_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n387_), .B1(new_n388_), .B2(new_n379_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n384_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT95), .ZN(new_n391_));
  OR2_X1    g190(.A1(G155gat), .A2(G162gat), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT1), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G155gat), .A2(G162gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n393_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G141gat), .A2(G148gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G141gat), .A2(G148gat), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n396_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT3), .ZN(new_n401_));
  INV_X1    g200(.A(G141gat), .ZN(new_n402_));
  INV_X1    g201(.A(G148gat), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT2), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n397_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n404_), .A2(new_n406_), .A3(new_n407_), .A4(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n392_), .A2(new_n394_), .ZN(new_n410_));
  AOI22_X1  g209(.A1(new_n395_), .A2(new_n400_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n390_), .B1(new_n391_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n409_), .A2(new_n410_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n396_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n398_), .A2(new_n399_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n395_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(new_n416_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n417_), .A2(new_n384_), .A3(KEYINPUT95), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n412_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G225gat), .A2(G233gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n411_), .A2(new_n384_), .A3(KEYINPUT4), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n411_), .A2(new_n391_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(new_n384_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n422_), .B1(new_n424_), .B2(KEYINPUT4), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n421_), .B1(new_n425_), .B2(new_n420_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G1gat), .B(G29gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(new_n215_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT0), .B(G57gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n428_), .B(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  OAI21_X1  g230(.A(KEYINPUT4), .B1(new_n412_), .B2(new_n418_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n422_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n420_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n420_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n424_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n430_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n431_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n389_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n442_));
  NAND2_X1  g241(.A1(G226gat), .A2(G233gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT93), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n364_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n367_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n448_), .A2(KEYINPUT92), .A3(new_n365_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n353_), .A2(new_n363_), .A3(KEYINPUT93), .A4(new_n354_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT92), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n451_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n447_), .A2(new_n449_), .A3(new_n450_), .A4(new_n452_), .ZN(new_n453_));
  OR2_X1    g252(.A1(new_n348_), .A2(new_n349_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT26), .B(G190gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n357_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n355_), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n454_), .A2(new_n456_), .A3(new_n457_), .A4(new_n345_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n453_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(G197gat), .ZN(new_n461_));
  INV_X1    g260(.A(G204gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT83), .B(G204gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n463_), .B1(new_n464_), .B2(new_n461_), .ZN(new_n465_));
  INV_X1    g264(.A(G218gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(G211gat), .ZN(new_n467_));
  INV_X1    g266(.A(G211gat), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(G218gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT21), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT84), .B1(new_n465_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n462_), .A2(KEYINPUT83), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT83), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n474_), .A2(G204gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(G197gat), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT84), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT21), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n479_), .B1(new_n467_), .B2(new_n469_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n477_), .A2(new_n478_), .A3(new_n463_), .A4(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n465_), .A2(new_n479_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n473_), .A2(new_n475_), .A3(new_n461_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n479_), .B1(G197gat), .B2(G204gat), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n470_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  AOI22_X1  g284(.A1(new_n472_), .A2(new_n481_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(KEYINPUT20), .B1(new_n460_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n472_), .A2(new_n481_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n482_), .A2(new_n485_), .ZN(new_n489_));
  AND3_X1   g288(.A1(new_n369_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n445_), .B1(new_n487_), .B2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(G8gat), .B(G36gat), .Z(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT18), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G64gat), .B(G92gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT20), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n496_), .B1(new_n460_), .B2(new_n486_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n488_), .A2(new_n489_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n369_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n497_), .A2(new_n444_), .A3(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n491_), .A2(new_n495_), .A3(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT27), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n497_), .A2(new_n500_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n445_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n496_), .B1(new_n498_), .B2(new_n459_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n486_), .A2(new_n369_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n444_), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n495_), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(KEYINPUT99), .B1(new_n503_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n495_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n508_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n444_), .B1(new_n497_), .B2(new_n500_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n511_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT99), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n514_), .A2(new_n515_), .A3(KEYINPUT27), .A4(new_n502_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n510_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n501_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n444_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n511_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n520_), .A2(KEYINPUT94), .A3(new_n502_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT27), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n518_), .A2(new_n519_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT94), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(new_n495_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n521_), .A2(new_n522_), .A3(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n517_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(G228gat), .ZN(new_n528_));
  INV_X1    g327(.A(G233gat), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT29), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n498_), .B(new_n531_), .C1(new_n532_), .C2(new_n411_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G78gat), .B(G106gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT87), .Z(new_n535_));
  XOR2_X1   g334(.A(new_n535_), .B(KEYINPUT88), .Z(new_n536_));
  INV_X1    g335(.A(KEYINPUT85), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n417_), .A2(new_n537_), .A3(KEYINPUT29), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT85), .B1(new_n411_), .B2(new_n532_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n498_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n540_), .A2(KEYINPUT86), .A3(new_n530_), .ZN(new_n541_));
  AOI21_X1  g340(.A(KEYINPUT86), .B1(new_n540_), .B2(new_n530_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n533_), .B(new_n536_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n411_), .A2(new_n532_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT28), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G22gat), .B(G50gat), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n546_), .A2(new_n547_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n543_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT86), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n537_), .B1(new_n417_), .B2(KEYINPUT29), .ZN(new_n553_));
  AOI211_X1 g352(.A(KEYINPUT85), .B(new_n532_), .C1(new_n413_), .C2(new_n416_), .ZN(new_n554_));
  NOR3_X1   g353(.A1(new_n486_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n552_), .B1(new_n555_), .B2(new_n531_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n540_), .A2(KEYINPUT86), .A3(new_n530_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n535_), .B1(new_n558_), .B2(new_n533_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT90), .B1(new_n551_), .B2(new_n559_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n533_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n535_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT90), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n563_), .A2(new_n564_), .A3(new_n550_), .A4(new_n543_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n543_), .A2(KEYINPUT89), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT89), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n558_), .A2(new_n567_), .A3(new_n533_), .A4(new_n536_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n536_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n561_), .A2(new_n569_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n566_), .A2(new_n568_), .A3(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n550_), .ZN(new_n572_));
  AOI22_X1  g371(.A1(new_n560_), .A2(new_n565_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n441_), .A2(new_n527_), .A3(new_n573_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n517_), .A2(new_n526_), .A3(new_n439_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n560_), .A2(new_n565_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n571_), .A2(new_n572_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n575_), .A2(new_n578_), .A3(KEYINPUT100), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT100), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n517_), .A2(new_n526_), .A3(new_n439_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n573_), .B2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT33), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT96), .B1(new_n437_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT96), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n426_), .A2(new_n585_), .A3(KEYINPUT33), .A4(new_n430_), .ZN(new_n586_));
  XOR2_X1   g385(.A(KEYINPUT97), .B(KEYINPUT33), .Z(new_n587_));
  NAND2_X1  g386(.A1(new_n437_), .A2(new_n587_), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n419_), .A2(new_n420_), .ZN(new_n589_));
  OAI21_X1  g388(.A(KEYINPUT98), .B1(new_n589_), .B2(new_n430_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n425_), .A2(new_n420_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n430_), .B1(new_n424_), .B2(new_n435_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT98), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n590_), .A2(new_n591_), .A3(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n584_), .A2(new_n586_), .A3(new_n588_), .A4(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n521_), .A2(new_n525_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n505_), .A2(new_n508_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n495_), .A2(KEYINPUT32), .ZN(new_n599_));
  MUX2_X1   g398(.A(new_n598_), .B(new_n523_), .S(new_n599_), .Z(new_n600_));
  OAI22_X1  g399(.A1(new_n596_), .A2(new_n597_), .B1(new_n439_), .B2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n573_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n579_), .A2(new_n582_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n574_), .B1(new_n603_), .B2(new_n389_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n290_), .B(new_n249_), .Z(new_n605_));
  NAND2_X1  g404(.A1(G229gat), .A2(G233gat), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n605_), .A2(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n297_), .A2(new_n249_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n609_), .B(new_n606_), .C1(new_n297_), .C2(new_n254_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G113gat), .B(G141gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G169gat), .B(G197gat), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n612_), .B(new_n613_), .Z(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n611_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n608_), .A2(new_n610_), .A3(new_n614_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  NOR2_X1   g418(.A1(new_n604_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n344_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT101), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n344_), .A2(KEYINPUT101), .A3(new_n620_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n439_), .A2(G1gat), .ZN(new_n625_));
  NAND4_X1  g424(.A1(new_n623_), .A2(KEYINPUT38), .A3(new_n624_), .A4(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n626_), .B(new_n627_), .ZN(new_n628_));
  OAI22_X1  g427(.A1(new_n341_), .A2(new_n337_), .B1(new_n312_), .B2(new_n311_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n338_), .A2(new_n339_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(new_n311_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n631_), .A2(new_n618_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n632_), .A2(new_n304_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n604_), .A2(new_n264_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT103), .ZN(new_n636_));
  OAI21_X1  g435(.A(G1gat), .B1(new_n636_), .B2(new_n439_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n628_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT38), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n639_), .A2(KEYINPUT104), .A3(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT104), .B1(new_n639_), .B2(new_n640_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n202_), .B1(new_n638_), .B2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n643_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n645_), .A2(KEYINPUT105), .A3(new_n628_), .A4(new_n637_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(G1324gat));
  INV_X1    g446(.A(new_n527_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n623_), .A2(new_n283_), .A3(new_n648_), .A4(new_n624_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n633_), .A2(new_n648_), .A3(new_n634_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT106), .B(KEYINPUT39), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n650_), .A2(G8gat), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n650_), .B2(G8gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  XOR2_X1   g453(.A(new_n654_), .B(KEYINPUT40), .Z(G1325gat));
  NOR3_X1   g454(.A1(new_n621_), .A2(G15gat), .A3(new_n389_), .ZN(new_n656_));
  INV_X1    g455(.A(G15gat), .ZN(new_n657_));
  INV_X1    g456(.A(new_n636_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n389_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n657_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  XOR2_X1   g459(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n661_));
  AOI21_X1  g460(.A(new_n656_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n662_), .B1(new_n660_), .B2(new_n661_), .ZN(G1326gat));
  OAI21_X1  g462(.A(G22gat), .B1(new_n636_), .B2(new_n573_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT42), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n578_), .A2(new_n280_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n621_), .B2(new_n666_), .ZN(G1327gat));
  NAND2_X1  g466(.A1(new_n603_), .A2(new_n389_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n574_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT43), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n264_), .B(new_n267_), .Z(new_n672_));
  NAND3_X1  g471(.A1(new_n670_), .A2(new_n671_), .A3(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(KEYINPUT43), .B1(new_n604_), .B2(new_n268_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n307_), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n618_), .B(new_n676_), .C1(new_n340_), .C2(new_n342_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n675_), .A2(KEYINPUT44), .A3(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(KEYINPUT109), .B(KEYINPUT44), .Z(new_n680_));
  INV_X1    g479(.A(KEYINPUT108), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n681_), .B1(new_n675_), .B2(new_n678_), .ZN(new_n682_));
  AOI211_X1 g481(.A(KEYINPUT108), .B(new_n677_), .C1(new_n673_), .C2(new_n674_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n680_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT110), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT110), .B(new_n680_), .C1(new_n682_), .C2(new_n683_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n679_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n688_), .A2(new_n440_), .ZN(new_n689_));
  INV_X1    g488(.A(G29gat), .ZN(new_n690_));
  INV_X1    g489(.A(new_n264_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n307_), .A2(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n631_), .A2(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n693_), .A2(new_n620_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n440_), .A2(new_n690_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT111), .ZN(new_n697_));
  OAI22_X1  g496(.A1(new_n689_), .A2(new_n690_), .B1(new_n695_), .B2(new_n697_), .ZN(G1328gat));
  INV_X1    g497(.A(G36gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n694_), .A2(new_n699_), .A3(new_n648_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT45), .ZN(new_n701_));
  OR2_X1    g500(.A1(new_n679_), .A2(new_n527_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n701_), .B1(new_n703_), .B2(new_n699_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(KEYINPUT46), .B(new_n701_), .C1(new_n703_), .C2(new_n699_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1329gat));
  NAND2_X1  g507(.A1(new_n659_), .A2(G43gat), .ZN(new_n709_));
  AOI211_X1 g508(.A(new_n679_), .B(new_n709_), .C1(new_n686_), .C2(new_n687_), .ZN(new_n710_));
  AOI21_X1  g509(.A(G43gat), .B1(new_n694_), .B2(new_n659_), .ZN(new_n711_));
  OAI21_X1  g510(.A(KEYINPUT47), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n688_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715_));
  INV_X1    g514(.A(new_n711_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n714_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n712_), .A2(new_n717_), .ZN(G1330gat));
  AOI21_X1  g517(.A(G50gat), .B1(new_n694_), .B2(new_n578_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n578_), .A2(G50gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n688_), .B2(new_n720_), .ZN(G1331gat));
  NOR2_X1   g520(.A1(new_n308_), .A2(new_n631_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n604_), .A2(new_n618_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(G57gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n725_), .A2(new_n726_), .A3(new_n440_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n619_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n728_));
  NOR4_X1   g527(.A1(new_n631_), .A2(new_n604_), .A3(new_n264_), .A4(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(new_n440_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n727_), .B1(new_n730_), .B2(new_n726_), .ZN(G1332gat));
  INV_X1    g530(.A(G64gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n729_), .B2(new_n648_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT48), .Z(new_n734_));
  NAND3_X1  g533(.A1(new_n725_), .A2(new_n732_), .A3(new_n648_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n734_), .A2(new_n735_), .ZN(G1333gat));
  INV_X1    g535(.A(G71gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n729_), .B2(new_n659_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT49), .Z(new_n739_));
  NAND2_X1  g538(.A1(new_n659_), .A2(new_n737_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n739_), .B1(new_n724_), .B2(new_n740_), .ZN(G1334gat));
  INV_X1    g540(.A(G78gat), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n742_), .B1(new_n729_), .B2(new_n578_), .ZN(new_n743_));
  XOR2_X1   g542(.A(new_n743_), .B(KEYINPUT50), .Z(new_n744_));
  NAND3_X1  g543(.A1(new_n725_), .A2(new_n742_), .A3(new_n578_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT112), .ZN(G1335gat));
  NAND3_X1  g546(.A1(new_n723_), .A2(new_n343_), .A3(new_n692_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n215_), .B1(new_n748_), .B2(new_n439_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT113), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n343_), .A2(new_n619_), .A3(new_n676_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n673_), .B2(new_n674_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n439_), .A2(new_n215_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n750_), .B1(new_n752_), .B2(new_n753_), .ZN(G1336gat));
  OAI21_X1  g553(.A(new_n216_), .B1(new_n748_), .B2(new_n527_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT114), .Z(new_n756_));
  NOR2_X1   g555(.A1(new_n527_), .A2(new_n216_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n752_), .B2(new_n757_), .ZN(G1337gat));
  OR2_X1    g557(.A1(new_n389_), .A2(new_n225_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT51), .ZN(new_n760_));
  OAI22_X1  g559(.A1(new_n748_), .A2(new_n759_), .B1(KEYINPUT115), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n752_), .A2(new_n659_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(G99gat), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n760_), .A2(KEYINPUT115), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n763_), .B(new_n764_), .Z(G1338gat));
  OR3_X1    g564(.A1(new_n748_), .A2(G106gat), .A3(new_n573_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n752_), .A2(new_n578_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT52), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n767_), .A2(new_n768_), .A3(G106gat), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n768_), .B1(new_n767_), .B2(G106gat), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n766_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g571(.A1(new_n307_), .A2(KEYINPUT116), .A3(new_n619_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n728_), .A2(new_n774_), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n268_), .A2(new_n773_), .A3(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT54), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n631_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(new_n631_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n329_), .A2(new_n331_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n326_), .A2(new_n327_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n782_), .A2(new_n320_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n322_), .B1(new_n783_), .B2(new_n328_), .ZN(new_n784_));
  OAI21_X1  g583(.A(KEYINPUT55), .B1(new_n333_), .B2(KEYINPUT117), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(new_n335_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n781_), .A2(new_n784_), .A3(new_n788_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n785_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n790_));
  OAI21_X1  g589(.A(KEYINPUT118), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n318_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n781_), .A2(new_n784_), .A3(new_n788_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT118), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n793_), .B(new_n794_), .C1(new_n332_), .C2(new_n785_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n791_), .A2(new_n792_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT56), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n605_), .A2(new_n606_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n297_), .A2(new_n254_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n609_), .A2(new_n607_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n798_), .B(new_n615_), .C1(new_n799_), .C2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n801_), .A2(new_n802_), .ZN(new_n804_));
  AND4_X1   g603(.A1(new_n617_), .A2(new_n339_), .A3(new_n803_), .A4(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n793_), .B1(new_n332_), .B2(new_n785_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n318_), .B1(new_n806_), .B2(KEYINPUT118), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n795_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n797_), .A2(new_n805_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT58), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n268_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n811_), .B2(new_n810_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT57), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT119), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n807_), .A2(new_n815_), .A3(new_n808_), .A4(new_n795_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n796_), .A2(KEYINPUT119), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n341_), .A2(new_n619_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n816_), .A2(new_n797_), .A3(new_n817_), .A4(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n630_), .A2(new_n617_), .A3(new_n803_), .A4(new_n804_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n814_), .B1(new_n821_), .B2(new_n691_), .ZN(new_n822_));
  AOI211_X1 g621(.A(KEYINPUT57), .B(new_n264_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n813_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n780_), .B1(new_n824_), .B2(new_n676_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n648_), .A2(new_n578_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n389_), .A2(new_n439_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OR3_X1    g627(.A1(new_n825_), .A2(KEYINPUT59), .A3(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n780_), .B1(new_n824_), .B2(new_n304_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT59), .B1(new_n830_), .B2(new_n828_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n829_), .A2(new_n831_), .A3(new_n618_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(G113gat), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n830_), .A2(new_n828_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  OR3_X1    g634(.A1(new_n835_), .A2(G113gat), .A3(new_n619_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n836_), .ZN(G1340gat));
  XOR2_X1   g636(.A(KEYINPUT121), .B(G120gat), .Z(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n631_), .B2(KEYINPUT60), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n834_), .B(new_n839_), .C1(KEYINPUT60), .C2(new_n838_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n829_), .A2(new_n343_), .A3(new_n831_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n841_), .B2(new_n838_), .ZN(G1341gat));
  INV_X1    g641(.A(new_n304_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n829_), .A2(new_n831_), .A3(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(G127gat), .ZN(new_n845_));
  OR3_X1    g644(.A1(new_n835_), .A2(G127gat), .A3(new_n676_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(G1342gat));
  NAND3_X1  g646(.A1(new_n829_), .A2(new_n831_), .A3(new_n672_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G134gat), .ZN(new_n849_));
  OR3_X1    g648(.A1(new_n835_), .A2(G134gat), .A3(new_n691_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1343gat));
  NOR3_X1   g650(.A1(new_n648_), .A2(new_n439_), .A3(new_n659_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n578_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n824_), .A2(new_n304_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n780_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n853_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n618_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n343_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g659(.A(KEYINPUT122), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n856_), .B2(new_n307_), .ZN(new_n862_));
  NOR4_X1   g661(.A1(new_n830_), .A2(KEYINPUT122), .A3(new_n676_), .A4(new_n853_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(KEYINPUT61), .B(G155gat), .ZN(new_n864_));
  INV_X1    g663(.A(new_n864_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n862_), .A2(new_n863_), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n853_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n264_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(new_n814_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n843_), .B1(new_n869_), .B2(new_n813_), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n307_), .B(new_n867_), .C1(new_n870_), .C2(new_n780_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT122), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n856_), .A2(new_n861_), .A3(new_n307_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n864_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n866_), .A2(new_n874_), .ZN(G1346gat));
  INV_X1    g674(.A(new_n856_), .ZN(new_n876_));
  OR3_X1    g675(.A1(new_n876_), .A2(G162gat), .A3(new_n691_), .ZN(new_n877_));
  OAI21_X1  g676(.A(G162gat), .B1(new_n876_), .B2(new_n268_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(G1347gat));
  NAND2_X1  g678(.A1(new_n824_), .A2(new_n676_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n855_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT22), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n648_), .A2(new_n441_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n578_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n881_), .A2(new_n882_), .A3(new_n618_), .A4(new_n884_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n885_), .A2(new_n346_), .A3(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n884_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n825_), .A2(new_n619_), .A3(new_n889_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n886_), .B1(new_n890_), .B2(new_n882_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n881_), .A2(new_n618_), .A3(new_n886_), .A4(new_n884_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(G169gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n888_), .B1(new_n891_), .B2(new_n893_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(G1348gat));
  NOR3_X1   g694(.A1(new_n825_), .A2(new_n631_), .A3(new_n889_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT124), .ZN(new_n897_));
  OR3_X1    g696(.A1(new_n896_), .A2(new_n897_), .A3(G176gat), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n896_), .B2(G176gat), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n830_), .A2(new_n578_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n631_), .A2(new_n347_), .A3(new_n883_), .ZN(new_n901_));
  AOI22_X1  g700(.A1(new_n898_), .A2(new_n899_), .B1(new_n900_), .B2(new_n901_), .ZN(G1349gat));
  NAND4_X1  g701(.A1(new_n900_), .A2(new_n648_), .A3(new_n441_), .A4(new_n307_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n825_), .A2(new_n889_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n304_), .A2(new_n357_), .ZN(new_n905_));
  AOI22_X1  g704(.A1(new_n903_), .A2(new_n362_), .B1(new_n904_), .B2(new_n905_), .ZN(G1350gat));
  NAND4_X1  g705(.A1(new_n881_), .A2(new_n455_), .A3(new_n264_), .A4(new_n884_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n825_), .A2(new_n268_), .A3(new_n889_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n908_), .B2(new_n358_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n907_), .B(KEYINPUT125), .C1(new_n908_), .C2(new_n358_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1351gat));
  NOR3_X1   g712(.A1(new_n573_), .A2(new_n659_), .A3(new_n440_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n527_), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(new_n915_), .B2(new_n914_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n830_), .A2(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n618_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g719(.A1(new_n918_), .A2(new_n343_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n464_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n462_), .B2(new_n921_), .ZN(G1353gat));
  NOR2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(KEYINPUT127), .ZN(new_n925_));
  NAND2_X1  g724(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n918_), .A2(new_n843_), .A3(new_n925_), .A4(new_n926_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n924_), .A2(KEYINPUT127), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n927_), .B(new_n928_), .ZN(G1354gat));
  NAND3_X1  g728(.A1(new_n918_), .A2(new_n466_), .A3(new_n264_), .ZN(new_n930_));
  NOR3_X1   g729(.A1(new_n830_), .A2(new_n268_), .A3(new_n917_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n931_), .B2(new_n466_), .ZN(G1355gat));
endmodule


