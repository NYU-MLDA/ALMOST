//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n846_, new_n847_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n908_, new_n909_, new_n911_, new_n912_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_;
  AND2_X1   g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G85gat), .B(G92gat), .Z(new_n203_));
  AOI21_X1  g002(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT66), .ZN(new_n206_));
  OAI211_X1 g005(.A(new_n206_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n205_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G99gat), .ZN(new_n210_));
  INV_X1    g009(.A(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT7), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n210_), .B(new_n211_), .C1(new_n212_), .C2(KEYINPUT66), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(KEYINPUT66), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n203_), .B1(new_n209_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT8), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT8), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n218_), .B(new_n203_), .C1(new_n209_), .C2(new_n215_), .ZN(new_n219_));
  XOR2_X1   g018(.A(KEYINPUT10), .B(G99gat), .Z(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT64), .B(G106gat), .Z(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT9), .ZN(new_n223_));
  INV_X1    g022(.A(G85gat), .ZN(new_n224_));
  INV_X1    g023(.A(G92gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n223_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n224_), .A2(new_n225_), .ZN(new_n230_));
  NAND4_X1  g029(.A1(KEYINPUT65), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n226_), .A2(new_n229_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n232_));
  AND3_X1   g031(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(new_n204_), .ZN(new_n234_));
  AND2_X1   g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  AOI22_X1  g034(.A1(new_n217_), .A2(new_n219_), .B1(new_n222_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G57gat), .A2(G64gat), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(G57gat), .A2(G64gat), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT11), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G57gat), .ZN(new_n241_));
  INV_X1    g040(.A(G64gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT11), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(new_n237_), .ZN(new_n245_));
  INV_X1    g044(.A(G78gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G71gat), .ZN(new_n247_));
  INV_X1    g046(.A(G71gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(G78gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n240_), .A2(new_n245_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n243_), .A2(new_n237_), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n252_), .A2(KEYINPUT11), .A3(new_n247_), .A4(new_n249_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n254_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n202_), .B1(new_n236_), .B2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n222_), .A2(new_n232_), .A3(new_n234_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n260_), .A2(KEYINPUT69), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(KEYINPUT69), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n234_), .A2(new_n207_), .A3(new_n214_), .A4(new_n213_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n218_), .B1(new_n263_), .B2(new_n203_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n219_), .ZN(new_n265_));
  OAI22_X1  g064(.A1(new_n261_), .A2(new_n262_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n251_), .A2(new_n253_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n254_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n255_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n266_), .A2(KEYINPUT12), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n260_), .B1(new_n265_), .B2(new_n264_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n270_), .ZN(new_n274_));
  XOR2_X1   g073(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n272_), .B1(new_n274_), .B2(new_n276_), .ZN(new_n277_));
  AOI211_X1 g076(.A(KEYINPUT71), .B(new_n275_), .C1(new_n273_), .C2(new_n270_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n259_), .B(new_n271_), .C1(new_n277_), .C2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n236_), .A2(new_n258_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n274_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n202_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT5), .B(G176gat), .ZN(new_n284_));
  INV_X1    g083(.A(G204gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G120gat), .B(G148gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n286_), .B(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n283_), .B(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n289_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G113gat), .B(G141gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G169gat), .B(G197gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G29gat), .B(G36gat), .ZN(new_n300_));
  INV_X1    g099(.A(G50gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT73), .B(G43gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n300_), .B(G50gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n306_), .A2(new_n303_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G1gat), .B(G8gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT79), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(G1gat), .ZN(new_n312_));
  INV_X1    g111(.A(G8gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT14), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT78), .B(G15gat), .ZN(new_n315_));
  INV_X1    g114(.A(G22gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n311_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n314_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n319_), .A2(new_n310_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n308_), .B1(new_n318_), .B2(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n310_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n311_), .A2(new_n314_), .A3(new_n317_), .ZN(new_n323_));
  OAI211_X1 g122(.A(new_n322_), .B(new_n323_), .C1(new_n305_), .C2(new_n307_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n321_), .A2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(G229gat), .A3(G233gat), .ZN(new_n326_));
  XOR2_X1   g125(.A(KEYINPUT74), .B(KEYINPUT15), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n328_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n302_), .A2(new_n304_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n306_), .A2(new_n303_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n330_), .A2(new_n331_), .A3(new_n327_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n329_), .A2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n318_), .A2(new_n320_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G229gat), .A2(G233gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n335_), .A2(new_n336_), .A3(new_n321_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n326_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n299_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  AOI211_X1 g139(.A(KEYINPUT82), .B(new_n298_), .C1(new_n326_), .C2(new_n337_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n295_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT98), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT29), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G155gat), .A2(G162gat), .ZN(new_n352_));
  AND3_X1   g151(.A1(new_n352_), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n353_));
  AOI21_X1  g152(.A(KEYINPUT89), .B1(new_n352_), .B2(KEYINPUT1), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G155gat), .A2(G162gat), .ZN(new_n356_));
  AND2_X1   g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n356_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n351_), .B1(new_n355_), .B2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n357_), .A2(new_n356_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT2), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n347_), .B1(new_n363_), .B2(KEYINPUT90), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT90), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n365_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n366_));
  AND2_X1   g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(G141gat), .ZN(new_n368_));
  INV_X1    g167(.A(G148gat), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n369_), .A3(KEYINPUT3), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT3), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n371_), .B1(G141gat), .B2(G148gat), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n370_), .A2(new_n372_), .B1(KEYINPUT90), .B2(new_n363_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n362_), .B1(new_n367_), .B2(new_n373_), .ZN(new_n374_));
  OAI21_X1  g173(.A(KEYINPUT91), .B1(new_n360_), .B2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n370_), .A2(new_n372_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n363_), .A2(KEYINPUT90), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n364_), .A2(new_n366_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n361_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT89), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n381_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n352_), .A2(KEYINPUT89), .A3(KEYINPUT1), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n359_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n350_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT91), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n380_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n346_), .B1(new_n375_), .B2(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G211gat), .B(G218gat), .Z(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G197gat), .B(G204gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT21), .ZN(new_n392_));
  NOR3_X1   g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT93), .ZN(new_n394_));
  INV_X1    g193(.A(G197gat), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(G204gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n285_), .A2(G197gat), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n396_), .A2(new_n397_), .A3(KEYINPUT92), .ZN(new_n398_));
  OAI21_X1  g197(.A(KEYINPUT21), .B1(new_n396_), .B2(KEYINPUT92), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n394_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n285_), .A2(G197gat), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT92), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n392_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n396_), .A2(new_n397_), .A3(KEYINPUT92), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n403_), .A2(KEYINPUT93), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n389_), .B1(new_n400_), .B2(new_n405_), .ZN(new_n406_));
  OR2_X1    g205(.A1(KEYINPUT94), .A2(KEYINPUT21), .ZN(new_n407_));
  NAND2_X1  g206(.A1(KEYINPUT94), .A2(KEYINPUT21), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n407_), .A2(new_n396_), .A3(new_n397_), .A4(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT95), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n391_), .A2(KEYINPUT95), .A3(new_n408_), .A4(new_n407_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n393_), .B1(new_n406_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G228gat), .A2(G233gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n388_), .A2(new_n414_), .A3(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n405_), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT93), .B1(new_n403_), .B2(new_n404_), .ZN(new_n419_));
  OAI211_X1 g218(.A(new_n413_), .B(new_n390_), .C1(new_n418_), .C2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n393_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT97), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT97), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n420_), .A2(new_n424_), .A3(new_n421_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n380_), .A2(new_n385_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT29), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT96), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT96), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n426_), .A2(new_n429_), .A3(KEYINPUT29), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n423_), .A2(new_n425_), .A3(new_n428_), .A4(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n417_), .B1(new_n431_), .B2(new_n416_), .ZN(new_n432_));
  XOR2_X1   g231(.A(G78gat), .B(G106gat), .Z(new_n433_));
  AOI21_X1  g232(.A(new_n345_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n375_), .A2(new_n346_), .A3(new_n387_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(G22gat), .B(G50gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT28), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n435_), .B(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n433_), .ZN(new_n440_));
  AOI211_X1 g239(.A(new_n440_), .B(new_n417_), .C1(new_n416_), .C2(new_n431_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n431_), .A2(new_n416_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n417_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n433_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  OAI22_X1  g243(.A1(new_n434_), .A2(new_n439_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n442_), .A2(new_n443_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n440_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n432_), .A2(new_n433_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n447_), .A2(new_n345_), .A3(new_n448_), .A4(new_n438_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n445_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G8gat), .B(G36gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(new_n225_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT18), .B(G64gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G226gat), .A2(G233gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT19), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  XNOR2_X1  g257(.A(KEYINPUT99), .B(KEYINPUT24), .ZN(new_n459_));
  OR2_X1    g258(.A1(G169gat), .A2(G176gat), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G183gat), .A2(G190gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT23), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT23), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(G183gat), .A3(G190gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G169gat), .A2(G176gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n459_), .A2(new_n467_), .A3(new_n460_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n461_), .A2(new_n466_), .A3(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT25), .B(G183gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT26), .B(G190gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n462_), .A2(new_n473_), .A3(KEYINPUT23), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n473_), .B1(new_n462_), .B2(KEYINPUT23), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n465_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(G183gat), .A2(G190gat), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n476_), .A2(new_n477_), .B1(G169gat), .B2(G176gat), .ZN(new_n478_));
  XNOR2_X1  g277(.A(KEYINPUT22), .B(G169gat), .ZN(new_n479_));
  INV_X1    g278(.A(G176gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n469_), .A2(new_n472_), .B1(new_n478_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT104), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n478_), .A2(new_n481_), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n461_), .A2(new_n468_), .A3(new_n466_), .A4(new_n472_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT104), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  AOI211_X1 g287(.A(KEYINPUT97), .B(new_n393_), .C1(new_n406_), .C2(new_n413_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n424_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n483_), .B(new_n488_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT20), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT26), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n493_), .A2(KEYINPUT84), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(KEYINPUT84), .ZN(new_n495_));
  OAI21_X1  g294(.A(G190gat), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT83), .B(G190gat), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n496_), .B(new_n470_), .C1(new_n493_), .C2(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n460_), .A2(KEYINPUT24), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n460_), .A2(KEYINPUT24), .A3(new_n467_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n498_), .A2(new_n499_), .A3(new_n500_), .A4(new_n476_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n466_), .B1(new_n497_), .B2(G183gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(KEYINPUT86), .A2(G169gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT22), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n502_), .B(new_n467_), .C1(G176gat), .C2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n492_), .B1(new_n422_), .B2(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n458_), .B1(new_n491_), .B2(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT20), .B1(new_n414_), .B2(new_n482_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n422_), .A2(new_n506_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n509_), .A2(new_n510_), .A3(new_n457_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n455_), .B1(new_n508_), .B2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT100), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n501_), .A2(new_n505_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT20), .B1(new_n514_), .B2(new_n414_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n458_), .B1(new_n422_), .B2(new_n486_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n513_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n457_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n457_), .B1(new_n414_), .B2(new_n482_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n519_), .A2(new_n507_), .A3(KEYINPUT100), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n517_), .A2(new_n518_), .A3(new_n454_), .A4(new_n520_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n512_), .A2(KEYINPUT27), .A3(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n517_), .A2(new_n518_), .A3(new_n520_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(new_n455_), .ZN(new_n524_));
  AOI21_X1  g323(.A(KEYINPUT27), .B1(new_n524_), .B2(new_n521_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G225gat), .A2(G233gat), .ZN(new_n527_));
  XOR2_X1   g326(.A(new_n527_), .B(KEYINPUT101), .Z(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G127gat), .B(G134gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G113gat), .B(G120gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n360_), .A2(new_n374_), .A3(KEYINPUT91), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n386_), .B1(new_n380_), .B2(new_n385_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n426_), .A2(new_n533_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(KEYINPUT4), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n532_), .B1(new_n375_), .B2(new_n387_), .ZN(new_n540_));
  XOR2_X1   g339(.A(KEYINPUT102), .B(KEYINPUT4), .Z(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n529_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n528_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n544_));
  XOR2_X1   g343(.A(G57gat), .B(G85gat), .Z(new_n545_));
  XNOR2_X1  g344(.A(G1gat), .B(G29gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT103), .B(KEYINPUT0), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NOR3_X1   g349(.A1(new_n543_), .A2(new_n544_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n550_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n501_), .A2(new_n556_), .A3(new_n505_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n556_), .B1(new_n501_), .B2(new_n505_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n533_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n506_), .A2(KEYINPUT30), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n561_), .A2(new_n532_), .A3(new_n557_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G71gat), .B(G99gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT31), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G227gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n563_), .A2(new_n568_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G15gat), .B(G43gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT87), .B(KEYINPUT88), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n570_), .B(new_n571_), .Z(new_n572_));
  NAND3_X1  g371(.A1(new_n560_), .A2(new_n562_), .A3(new_n567_), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n569_), .A2(new_n572_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n572_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND4_X1  g375(.A1(new_n450_), .A2(new_n526_), .A3(new_n555_), .A4(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n454_), .A2(KEYINPUT32), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n508_), .B2(new_n511_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n517_), .A2(new_n518_), .A3(new_n578_), .A4(new_n520_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n542_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT4), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n540_), .A2(new_n583_), .A3(new_n537_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n528_), .B1(new_n582_), .B2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n544_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n549_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  OAI211_X1 g386(.A(new_n580_), .B(new_n581_), .C1(new_n587_), .C2(new_n551_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT33), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n553_), .A2(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(KEYINPUT33), .B(new_n550_), .C1(new_n543_), .C2(new_n544_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n539_), .A2(new_n529_), .A3(new_n542_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n536_), .A2(new_n528_), .A3(new_n538_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(new_n549_), .A3(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n524_), .A2(new_n521_), .A3(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n588_), .B1(new_n592_), .B2(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n554_), .B1(new_n445_), .B2(new_n449_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n450_), .A2(new_n597_), .B1(new_n598_), .B2(new_n526_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n577_), .B1(new_n599_), .B2(new_n576_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n344_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n270_), .B(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(new_n334_), .Z(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G183gat), .B(G211gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n610_), .A2(KEYINPUT17), .ZN(new_n611_));
  AOI21_X1  g410(.A(KEYINPUT81), .B1(new_n605_), .B2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n610_), .A2(KEYINPUT17), .ZN(new_n613_));
  OR3_X1    g412(.A1(new_n605_), .A2(new_n611_), .A3(new_n613_), .ZN(new_n614_));
  MUX2_X1   g413(.A(KEYINPUT81), .B(new_n612_), .S(new_n614_), .Z(new_n615_));
  XNOR2_X1  g414(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n616_));
  NAND2_X1  g415(.A1(G232gat), .A2(G233gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT34), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n308_), .A2(new_n236_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT75), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n333_), .A2(new_n266_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  OAI211_X1 g421(.A(KEYINPUT35), .B(new_n618_), .C1(new_n620_), .C2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT75), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n619_), .B(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n618_), .A2(KEYINPUT35), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n618_), .A2(KEYINPUT35), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .A4(new_n621_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n623_), .A2(KEYINPUT76), .A3(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G190gat), .B(G218gat), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G134gat), .B(G162gat), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n630_), .B(new_n631_), .Z(new_n632_));
  INV_X1    g431(.A(KEYINPUT36), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n629_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n634_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n623_), .A2(new_n628_), .A3(KEYINPUT76), .A4(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n632_), .A2(new_n633_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n623_), .B2(new_n628_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n616_), .B1(new_n638_), .B2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n616_), .ZN(new_n644_));
  AOI211_X1 g443(.A(new_n641_), .B(new_n644_), .C1(new_n635_), .C2(new_n637_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n601_), .A2(new_n615_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n554_), .B(KEYINPUT105), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n649_), .A2(new_n312_), .A3(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT38), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n638_), .A2(new_n642_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT106), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n525_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n512_), .A2(KEYINPUT27), .A3(new_n521_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n576_), .A2(new_n445_), .A3(new_n449_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n658_), .A2(new_n659_), .A3(new_n554_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n450_), .A2(new_n597_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n445_), .A2(new_n449_), .ZN(new_n662_));
  NAND4_X1  g461(.A1(new_n662_), .A2(new_n555_), .A3(new_n656_), .A4(new_n657_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n661_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n576_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n660_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n655_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n667_), .A2(new_n615_), .A3(new_n344_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G1gat), .B1(new_n668_), .B2(new_n555_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n652_), .A2(new_n669_), .ZN(G1324gat));
  OAI21_X1  g469(.A(G8gat), .B1(new_n668_), .B2(new_n526_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT39), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n649_), .A2(new_n313_), .A3(new_n658_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT107), .B(KEYINPUT40), .Z(new_n675_));
  XNOR2_X1  g474(.A(new_n674_), .B(new_n675_), .ZN(G1325gat));
  OAI21_X1  g475(.A(G15gat), .B1(new_n668_), .B2(new_n665_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT41), .ZN(new_n678_));
  NOR3_X1   g477(.A1(new_n648_), .A2(G15gat), .A3(new_n665_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT108), .ZN(G1326gat));
  OAI21_X1  g480(.A(G22gat), .B1(new_n668_), .B2(new_n450_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT42), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n649_), .A2(new_n316_), .A3(new_n662_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1327gat));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n576_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n686_), .B(new_n646_), .C1(new_n687_), .C2(new_n660_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT109), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT43), .B1(new_n666_), .B2(new_n647_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT109), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n600_), .A2(new_n691_), .A3(new_n686_), .A4(new_n646_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n689_), .A2(new_n690_), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n615_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n693_), .A2(new_n694_), .A3(new_n344_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n693_), .A2(KEYINPUT44), .A3(new_n694_), .A4(new_n344_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n650_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G29gat), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n653_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n615_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n601_), .A2(new_n703_), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n704_), .A2(G29gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n555_), .B2(new_n705_), .ZN(G1328gat));
  NAND3_X1  g505(.A1(new_n697_), .A2(new_n658_), .A3(new_n698_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n697_), .A2(KEYINPUT110), .A3(new_n658_), .A4(new_n698_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n709_), .A2(G36gat), .A3(new_n710_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n704_), .A2(G36gat), .A3(new_n526_), .ZN(new_n712_));
  XOR2_X1   g511(.A(new_n712_), .B(KEYINPUT45), .Z(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n711_), .A2(KEYINPUT46), .A3(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1329gat));
  INV_X1    g517(.A(G43gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n719_), .B1(new_n704_), .B2(new_n665_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n697_), .A2(G43gat), .A3(new_n576_), .A4(new_n698_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n721_), .A2(new_n722_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT47), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT47), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n727_), .B(new_n720_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1330gat));
  OAI21_X1  g528(.A(G50gat), .B1(new_n699_), .B2(new_n450_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n662_), .A2(new_n301_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT112), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n730_), .B1(new_n704_), .B2(new_n732_), .ZN(G1331gat));
  NOR2_X1   g532(.A1(new_n294_), .A2(new_n342_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n600_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n615_), .A3(new_n647_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT113), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n737_), .B(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G57gat), .B1(new_n739_), .B2(new_n650_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT114), .Z(new_n741_));
  NAND3_X1  g540(.A1(new_n667_), .A2(new_n615_), .A3(new_n734_), .ZN(new_n742_));
  NOR3_X1   g541(.A1(new_n742_), .A2(new_n241_), .A3(new_n555_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1332gat));
  OAI21_X1  g543(.A(G64gat), .B1(new_n742_), .B2(new_n526_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT48), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n739_), .A2(new_n242_), .A3(new_n658_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1333gat));
  OAI21_X1  g547(.A(G71gat), .B1(new_n742_), .B2(new_n665_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT49), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n739_), .A2(new_n248_), .A3(new_n576_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1334gat));
  OAI21_X1  g551(.A(G78gat), .B1(new_n742_), .B2(new_n450_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT50), .ZN(new_n754_));
  INV_X1    g553(.A(new_n739_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n662_), .A2(new_n246_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT115), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n754_), .B1(new_n755_), .B2(new_n757_), .ZN(G1335gat));
  NAND2_X1  g557(.A1(new_n736_), .A2(new_n703_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n650_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n693_), .A2(new_n694_), .A3(new_n734_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n762_), .A2(new_n555_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n763_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g563(.A(G92gat), .B1(new_n760_), .B2(new_n658_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n762_), .A2(new_n526_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G92gat), .ZN(G1337gat));
  INV_X1    g566(.A(new_n762_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n210_), .B1(new_n768_), .B2(new_n576_), .ZN(new_n769_));
  AND2_X1   g568(.A1(new_n576_), .A2(new_n220_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n760_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(KEYINPUT51), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(KEYINPUT51), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n775_), .A2(KEYINPUT117), .ZN(new_n776_));
  AOI22_X1  g575(.A1(new_n773_), .A2(new_n775_), .B1(new_n771_), .B2(new_n776_), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n760_), .A2(new_n662_), .A3(new_n221_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n768_), .A2(new_n662_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n780_), .B2(G106gat), .ZN(new_n781_));
  AOI211_X1 g580(.A(KEYINPUT52), .B(new_n211_), .C1(new_n768_), .C2(new_n662_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g583(.A1(new_n647_), .A2(new_n615_), .A3(new_n343_), .A4(new_n294_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT54), .ZN(new_n786_));
  OR2_X1    g585(.A1(new_n283_), .A2(new_n288_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n336_), .B1(new_n335_), .B2(new_n321_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n321_), .A2(new_n324_), .A3(new_n336_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n298_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n326_), .A2(new_n337_), .A3(new_n299_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n787_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT118), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n787_), .A2(new_n792_), .A3(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n280_), .B(new_n271_), .C1(new_n277_), .C2(new_n278_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n202_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n279_), .A2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n276_), .B1(new_n236_), .B2(new_n258_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT71), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n274_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n805_), .A2(KEYINPUT55), .A3(new_n259_), .A4(new_n271_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n799_), .A2(new_n801_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT56), .B1(new_n807_), .B2(new_n288_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n807_), .A2(KEYINPUT56), .A3(new_n288_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n808_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  AOI211_X1 g610(.A(KEYINPUT119), .B(KEYINPUT56), .C1(new_n807_), .C2(new_n288_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n797_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT58), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n797_), .B(KEYINPUT58), .C1(new_n811_), .C2(new_n812_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n646_), .A3(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n807_), .A2(KEYINPUT56), .A3(new_n288_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n342_), .B(new_n787_), .C1(new_n819_), .C2(new_n808_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n289_), .A2(new_n792_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n818_), .B1(new_n822_), .B2(new_n702_), .ZN(new_n823_));
  AOI211_X1 g622(.A(KEYINPUT57), .B(new_n653_), .C1(new_n820_), .C2(new_n821_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n817_), .B(KEYINPUT120), .C1(new_n823_), .C2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n694_), .ZN(new_n826_));
  OR2_X1    g625(.A1(new_n823_), .A2(new_n824_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT120), .B1(new_n827_), .B2(new_n817_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n786_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n700_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(G113gat), .B1(new_n831_), .B2(new_n342_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(G113gat), .ZN(new_n835_));
  INV_X1    g634(.A(new_n817_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n823_), .A2(new_n824_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n694_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n786_), .A2(new_n838_), .ZN(new_n839_));
  XOR2_X1   g638(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n840_));
  AND3_X1   g639(.A1(new_n839_), .A2(new_n830_), .A3(new_n840_), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n834_), .A2(new_n835_), .A3(new_n841_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n832_), .B1(new_n842_), .B2(new_n342_), .ZN(G1340gat));
  INV_X1    g642(.A(G120gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n844_), .B1(new_n294_), .B2(KEYINPUT60), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n831_), .B(new_n845_), .C1(KEYINPUT60), .C2(new_n844_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n834_), .A2(new_n294_), .A3(new_n841_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n844_), .ZN(G1341gat));
  AOI21_X1  g647(.A(G127gat), .B1(new_n831_), .B2(new_n615_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n834_), .A2(new_n841_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n615_), .A2(G127gat), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT122), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n849_), .B1(new_n850_), .B2(new_n852_), .ZN(G1342gat));
  AOI21_X1  g652(.A(G134gat), .B1(new_n831_), .B2(new_n655_), .ZN(new_n854_));
  INV_X1    g653(.A(G134gat), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n834_), .A2(new_n855_), .A3(new_n841_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n854_), .B1(new_n856_), .B2(new_n646_), .ZN(G1343gat));
  NOR2_X1   g656(.A1(new_n658_), .A2(new_n450_), .ZN(new_n858_));
  NAND4_X1  g657(.A1(new_n829_), .A2(new_n665_), .A3(new_n650_), .A4(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT123), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n862_), .A2(new_n694_), .A3(new_n825_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n576_), .B1(new_n863_), .B2(new_n786_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n864_), .A2(new_n865_), .A3(new_n650_), .A4(new_n858_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n860_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n342_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n868_), .A2(G141gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n867_), .A2(new_n368_), .A3(new_n342_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1344gat));
  NAND2_X1  g670(.A1(new_n867_), .A2(new_n295_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G148gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n867_), .A2(new_n369_), .A3(new_n295_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1345gat));
  XNOR2_X1  g674(.A(KEYINPUT61), .B(G155gat), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n876_), .B1(new_n867_), .B2(new_n615_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n876_), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n694_), .B(new_n878_), .C1(new_n860_), .C2(new_n866_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n877_), .A2(new_n879_), .ZN(G1346gat));
  AOI21_X1  g679(.A(G162gat), .B1(new_n867_), .B2(new_n655_), .ZN(new_n881_));
  INV_X1    g680(.A(G162gat), .ZN(new_n882_));
  AOI211_X1 g681(.A(new_n882_), .B(new_n647_), .C1(new_n860_), .C2(new_n866_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n881_), .A2(new_n883_), .ZN(G1347gat));
  NOR3_X1   g683(.A1(new_n650_), .A2(new_n526_), .A3(new_n659_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n839_), .A2(new_n342_), .A3(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(KEYINPUT124), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n839_), .A2(new_n888_), .A3(new_n342_), .A4(new_n885_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n887_), .A2(G169gat), .A3(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT125), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT125), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n887_), .A2(new_n892_), .A3(G169gat), .A4(new_n889_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n891_), .A2(KEYINPUT62), .A3(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n839_), .A2(new_n885_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n479_), .A3(new_n342_), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n890_), .A2(KEYINPUT125), .A3(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n894_), .A2(new_n897_), .A3(new_n899_), .ZN(G1348gat));
  AND3_X1   g699(.A1(new_n829_), .A2(new_n295_), .A3(new_n885_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n295_), .A2(new_n480_), .ZN(new_n902_));
  OAI22_X1  g701(.A1(new_n901_), .A2(new_n480_), .B1(new_n895_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT126), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1349gat));
  NOR2_X1   g704(.A1(new_n895_), .A2(new_n694_), .ZN(new_n906_));
  MUX2_X1   g705(.A(G183gat), .B(new_n470_), .S(new_n906_), .Z(G1350gat));
  OAI21_X1  g706(.A(G190gat), .B1(new_n895_), .B2(new_n647_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n655_), .A2(new_n471_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n895_), .B2(new_n909_), .ZN(G1351gat));
  AND2_X1   g709(.A1(new_n864_), .A2(new_n598_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(new_n658_), .A3(new_n342_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g712(.A1(new_n911_), .A2(new_n658_), .A3(new_n295_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g714(.A(new_n694_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n911_), .A2(new_n658_), .A3(new_n916_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT127), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n917_), .B(new_n919_), .ZN(G1354gat));
  AND3_X1   g719(.A1(new_n911_), .A2(G218gat), .A3(new_n658_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n911_), .A2(new_n658_), .A3(new_n655_), .ZN(new_n922_));
  INV_X1    g721(.A(G218gat), .ZN(new_n923_));
  AOI22_X1  g722(.A1(new_n921_), .A2(new_n646_), .B1(new_n922_), .B2(new_n923_), .ZN(G1355gat));
endmodule


