//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 0 0 0 1 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n766_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n921_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_;
  INV_X1    g000(.A(KEYINPUT12), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT10), .B(G99gat), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n203_), .B1(new_n204_), .B2(G106gat), .ZN(new_n205_));
  INV_X1    g004(.A(G85gat), .ZN(new_n206_));
  INV_X1    g005(.A(G92gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G85gat), .A2(G92gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n208_), .A2(KEYINPUT9), .A3(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT9), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G85gat), .A3(G92gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n216_));
  AND3_X1   g015(.A1(new_n213_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n218_));
  INV_X1    g017(.A(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n218_), .A2(KEYINPUT65), .A3(new_n219_), .A4(new_n220_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n205_), .A2(new_n210_), .A3(new_n217_), .A4(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT7), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n224_), .A3(new_n219_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n225_), .A2(new_n213_), .A3(new_n216_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n208_), .A2(new_n209_), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n228_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n222_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n202_), .B1(new_n232_), .B2(KEYINPUT66), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G57gat), .B(G64gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G71gat), .B(G78gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(KEYINPUT11), .ZN(new_n236_));
  XOR2_X1   g035(.A(G71gat), .B(G78gat), .Z(new_n237_));
  INV_X1    g036(.A(G64gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G57gat), .ZN(new_n239_));
  INV_X1    g038(.A(G57gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G64gat), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n241_), .A3(KEYINPUT11), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n234_), .A2(KEYINPUT11), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n236_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n227_), .A2(new_n229_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT8), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n245_), .B1(new_n249_), .B2(new_n222_), .ZN(new_n250_));
  OAI211_X1 g049(.A(new_n245_), .B(new_n222_), .C1(new_n230_), .C2(new_n231_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n233_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n245_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n232_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT66), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n256_), .B1(new_n249_), .B2(new_n222_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n255_), .B1(new_n257_), .B2(new_n202_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G230gat), .A2(G233gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT64), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n253_), .A2(new_n258_), .A3(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n260_), .B1(new_n250_), .B2(new_n252_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G120gat), .B(G148gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(G176gat), .B(G204gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n264_), .A2(new_n270_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n262_), .A2(new_n263_), .A3(new_n269_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(KEYINPUT13), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n274_), .A2(KEYINPUT68), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(KEYINPUT68), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(G183gat), .ZN(new_n280_));
  INV_X1    g079(.A(G190gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT23), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n280_), .A2(KEYINPUT23), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT79), .B1(new_n283_), .B2(G190gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT23), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n285_), .A2(KEYINPUT79), .A3(G183gat), .A4(G190gat), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n282_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  NOR3_X1   g087(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(KEYINPUT80), .A3(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT80), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n285_), .B1(G183gat), .B2(G190gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n285_), .A2(G183gat), .A3(G190gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT79), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n293_), .B1(new_n296_), .B2(new_n286_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n292_), .B1(new_n297_), .B2(new_n289_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT25), .B(G183gat), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT77), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(new_n281_), .B2(KEYINPUT26), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n281_), .A2(KEYINPUT26), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n281_), .A2(KEYINPUT26), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT77), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT78), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  OR2_X1    g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT24), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AOI22_X1  g110(.A1(new_n302_), .A2(new_n305_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n291_), .A2(new_n298_), .A3(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT22), .B(G169gat), .ZN(new_n314_));
  INV_X1    g113(.A(G176gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n308_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT81), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n282_), .A2(new_n294_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT81), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n316_), .A2(new_n308_), .A3(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n318_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n313_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G197gat), .B(G204gat), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT21), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G211gat), .B(G218gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n327_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n330_), .B1(new_n333_), .B2(KEYINPUT21), .ZN(new_n334_));
  INV_X1    g133(.A(G197gat), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n335_), .A2(KEYINPUT87), .A3(G204gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT21), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT87), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n337_), .B1(new_n338_), .B2(new_n327_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n332_), .B1(new_n334_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n326_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G226gat), .A2(G233gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT19), .ZN(new_n343_));
  INV_X1    g142(.A(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT20), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n288_), .A2(new_n321_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n317_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n289_), .B1(new_n282_), .B2(new_n294_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT26), .B(G190gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(new_n299_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n306_), .A2(KEYINPUT24), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT89), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n306_), .A2(KEYINPUT89), .A3(KEYINPUT24), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n309_), .A3(new_n355_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n346_), .A2(new_n347_), .B1(new_n351_), .B2(new_n356_), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n331_), .B1(new_n328_), .B2(new_n327_), .ZN(new_n358_));
  OAI211_X1 g157(.A(KEYINPUT21), .B(new_n336_), .C1(new_n333_), .C2(KEYINPUT87), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n358_), .A2(new_n359_), .B1(new_n331_), .B2(new_n329_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n345_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n341_), .A2(new_n344_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT90), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND4_X1  g163(.A1(new_n341_), .A2(KEYINPUT90), .A3(new_n344_), .A4(new_n361_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n343_), .B(KEYINPUT88), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n313_), .A2(new_n360_), .A3(new_n325_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n356_), .A2(new_n350_), .A3(new_n348_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n297_), .A2(new_n320_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(new_n317_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n345_), .B1(new_n370_), .B2(new_n340_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n366_), .B1(new_n367_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n364_), .A2(new_n365_), .A3(new_n373_), .ZN(new_n374_));
  XOR2_X1   g173(.A(G8gat), .B(G36gat), .Z(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n379_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n364_), .A2(new_n365_), .A3(new_n381_), .A4(new_n373_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT27), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n360_), .B1(new_n313_), .B2(new_n325_), .ZN(new_n384_));
  OAI21_X1  g183(.A(KEYINPUT20), .B1(new_n370_), .B2(new_n340_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n343_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT96), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  OAI211_X1 g187(.A(KEYINPUT96), .B(new_n343_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n367_), .A2(new_n371_), .A3(new_n366_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n388_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT98), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n391_), .A2(new_n392_), .A3(new_n379_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n382_), .A2(KEYINPUT27), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n392_), .B1(new_n391_), .B2(new_n379_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n383_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT99), .ZN(new_n399_));
  INV_X1    g198(.A(G141gat), .ZN(new_n400_));
  INV_X1    g199(.A(G148gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G141gat), .A2(G148gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NOR2_X1   g203(.A1(G155gat), .A2(G162gat), .ZN(new_n405_));
  AND2_X1   g204(.A1(G155gat), .A2(G162gat), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT1), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n405_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(G155gat), .ZN(new_n409_));
  INV_X1    g208(.A(G162gat), .ZN(new_n410_));
  OAI21_X1  g209(.A(KEYINPUT1), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n404_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n402_), .B2(KEYINPUT3), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n403_), .A2(KEYINPUT2), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT2), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(G141gat), .A3(G148gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n415_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n402_), .A2(KEYINPUT3), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT3), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n420_), .A2(new_n400_), .A3(new_n401_), .A4(KEYINPUT84), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n414_), .A2(new_n418_), .A3(new_n419_), .A4(new_n421_), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n406_), .A2(new_n405_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n412_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT28), .B1(new_n425_), .B2(KEYINPUT29), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT28), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT29), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G22gat), .B(G50gat), .ZN(new_n431_));
  AND2_X1   g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n430_), .A2(new_n431_), .ZN(new_n433_));
  OR2_X1    g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G228gat), .A2(G233gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(KEYINPUT86), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n435_), .A2(KEYINPUT86), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n436_), .B(new_n437_), .C1(new_n360_), .C2(KEYINPUT85), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n340_), .B1(new_n424_), .B2(new_n428_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(G78gat), .ZN(new_n440_));
  INV_X1    g239(.A(G78gat), .ZN(new_n441_));
  OAI211_X1 g240(.A(new_n340_), .B(new_n441_), .C1(new_n424_), .C2(new_n428_), .ZN(new_n442_));
  AOI21_X1  g241(.A(G106gat), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n440_), .A2(G106gat), .A3(new_n442_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n438_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n445_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n438_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n447_), .A2(new_n443_), .A3(new_n448_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n434_), .B1(new_n446_), .B2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n432_), .A2(new_n433_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n448_), .B1(new_n447_), .B2(new_n443_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n444_), .A2(new_n445_), .A3(new_n438_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n451_), .A2(new_n452_), .A3(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n450_), .A2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(G71gat), .B(G99gat), .Z(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(G43gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT30), .ZN(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G227gat), .A2(G233gat), .ZN(new_n460_));
  INV_X1    g259(.A(G15gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n326_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n326_), .A2(new_n462_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n459_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n465_), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n468_), .A2(new_n458_), .A3(new_n463_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G127gat), .B(G134gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G113gat), .B(G120gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT31), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT82), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n471_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n467_), .A2(new_n470_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n477_), .B1(new_n471_), .B2(new_n475_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n466_), .B2(new_n469_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G1gat), .B(G29gat), .Z(new_n482_));
  XNOR2_X1  g281(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G57gat), .B(G85gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n474_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n422_), .A2(new_n423_), .ZN(new_n488_));
  OAI211_X1 g287(.A(KEYINPUT92), .B(new_n487_), .C1(new_n488_), .C2(new_n412_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT92), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n490_), .B1(new_n424_), .B2(new_n474_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT93), .B1(new_n425_), .B2(new_n487_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT93), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n424_), .A2(new_n494_), .A3(new_n474_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n492_), .A2(KEYINPUT4), .A3(new_n493_), .A4(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G225gat), .A2(G233gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n424_), .A2(new_n474_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT4), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n497_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n493_), .A2(new_n495_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n502_), .A2(new_n497_), .A3(new_n492_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n486_), .B1(new_n501_), .B2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n501_), .A2(new_n503_), .A3(new_n486_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n481_), .A2(new_n507_), .ZN(new_n508_));
  NAND4_X1  g307(.A1(new_n398_), .A2(new_n399_), .A3(new_n455_), .A4(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT27), .ZN(new_n510_));
  AND4_X1   g309(.A1(new_n381_), .A2(new_n364_), .A3(new_n365_), .A4(new_n373_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n372_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n381_), .B1(new_n512_), .B2(new_n365_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n510_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n391_), .A2(new_n392_), .A3(new_n379_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n515_), .A2(KEYINPUT27), .A3(new_n382_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n514_), .B(new_n455_), .C1(new_n516_), .C2(new_n396_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n481_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n507_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(KEYINPUT99), .B1(new_n517_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n509_), .A2(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n511_), .A2(new_n513_), .ZN(new_n523_));
  AND3_X1   g322(.A1(new_n501_), .A2(new_n503_), .A3(new_n486_), .ZN(new_n524_));
  OAI21_X1  g323(.A(KEYINPUT95), .B1(new_n524_), .B2(KEYINPUT33), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT95), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT33), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n506_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n501_), .A2(new_n503_), .A3(KEYINPUT33), .A4(new_n486_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n497_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n496_), .A2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n502_), .A2(new_n530_), .A3(new_n492_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n486_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n532_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  AND2_X1   g334(.A1(new_n529_), .A2(new_n535_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n523_), .A2(new_n525_), .A3(new_n528_), .A4(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n381_), .A2(KEYINPUT32), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n512_), .A2(new_n365_), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n539_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n391_), .A2(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n507_), .A2(new_n538_), .A3(new_n540_), .A4(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(new_n542_), .B(new_n540_), .C1(new_n524_), .C2(new_n504_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n544_), .A2(KEYINPUT97), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n537_), .A2(new_n543_), .A3(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n455_), .A2(new_n507_), .ZN(new_n547_));
  AOI22_X1  g346(.A1(new_n546_), .A2(new_n455_), .B1(new_n398_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n522_), .B1(new_n548_), .B2(new_n518_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G1gat), .B(G8gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(KEYINPUT71), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G15gat), .B(G22gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G1gat), .A2(G8gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT14), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n552_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n550_), .A2(KEYINPUT71), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n550_), .A2(KEYINPUT71), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n557_), .A2(new_n554_), .A3(new_n552_), .A4(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n556_), .A2(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G29gat), .B(G36gat), .Z(new_n561_));
  XOR2_X1   g360(.A(G43gat), .B(G50gat), .Z(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G29gat), .B(G36gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G43gat), .B(G50gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n560_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT74), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT74), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n560_), .A2(new_n570_), .A3(new_n567_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n560_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n567_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n572_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G229gat), .A2(G233gat), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(KEYINPUT75), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT75), .ZN(new_n580_));
  AOI22_X1  g379(.A1(new_n569_), .A2(new_n571_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n581_), .B2(new_n577_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n567_), .B(KEYINPUT15), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n573_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n572_), .A2(new_n577_), .A3(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n579_), .A2(new_n582_), .A3(new_n585_), .ZN(new_n586_));
  XOR2_X1   g385(.A(G113gat), .B(G141gat), .Z(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT76), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G169gat), .B(G197gat), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n588_), .B(new_n589_), .Z(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n579_), .A2(new_n582_), .A3(new_n585_), .A4(new_n590_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n549_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT100), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n549_), .A2(KEYINPUT100), .A3(new_n594_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n279_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(KEYINPUT35), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n583_), .B2(new_n232_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n249_), .A2(new_n567_), .A3(new_n222_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n603_), .A2(KEYINPUT35), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT70), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n608_), .A2(KEYINPUT70), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G134gat), .B(G162gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n615_), .A2(KEYINPUT36), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n612_), .A2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n615_), .B(KEYINPUT36), .Z(new_n619_));
  NAND2_X1  g418(.A1(new_n612_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n621_), .A2(KEYINPUT37), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT37), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n618_), .A2(new_n623_), .A3(new_n620_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT72), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n560_), .B(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(new_n254_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(G127gat), .B(G155gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G183gat), .B(G211gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT17), .ZN(new_n636_));
  OR3_X1    g435(.A1(new_n635_), .A2(KEYINPUT66), .A3(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n636_), .ZN(new_n638_));
  AND2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n630_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n630_), .A2(new_n637_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n626_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n599_), .A2(new_n643_), .ZN(new_n644_));
  OR3_X1    g443(.A1(new_n644_), .A2(G1gat), .A3(new_n519_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT38), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n642_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n278_), .A2(new_n648_), .A3(new_n594_), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n649_), .A2(KEYINPUT101), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n612_), .A2(new_n617_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n651_), .B1(new_n612_), .B2(new_n619_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT102), .ZN(new_n653_));
  AND2_X1   g452(.A1(new_n549_), .A2(new_n653_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n649_), .A2(KEYINPUT101), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n650_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT103), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n507_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(G1gat), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n645_), .A2(new_n646_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n647_), .A2(new_n659_), .A3(new_n660_), .ZN(G1324gat));
  OAI21_X1  g460(.A(G8gat), .B1(new_n656_), .B2(new_n398_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT39), .ZN(new_n663_));
  OR3_X1    g462(.A1(new_n644_), .A2(G8gat), .A3(new_n398_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n663_), .A2(new_n664_), .A3(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1325gat));
  INV_X1    g467(.A(new_n644_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n669_), .A2(new_n461_), .A3(new_n518_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n657_), .A2(new_n518_), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n671_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(KEYINPUT41), .B1(new_n671_), .B2(G15gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n672_), .B2(new_n673_), .ZN(G1326gat));
  INV_X1    g473(.A(G22gat), .ZN(new_n675_));
  INV_X1    g474(.A(new_n455_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n669_), .A2(new_n675_), .A3(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n657_), .A2(new_n676_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(G22gat), .ZN(new_n680_));
  AOI211_X1 g479(.A(KEYINPUT42), .B(new_n675_), .C1(new_n657_), .C2(new_n676_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n677_), .B1(new_n680_), .B2(new_n681_), .ZN(G1327gat));
  NOR2_X1   g481(.A1(new_n621_), .A2(new_n648_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n599_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G29gat), .B1(new_n685_), .B2(new_n507_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n278_), .A2(new_n642_), .A3(new_n594_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT43), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n625_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n622_), .A2(KEYINPUT106), .A3(new_n624_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT105), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n549_), .B2(new_n694_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n522_), .B(KEYINPUT105), .C1(new_n548_), .C2(new_n518_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n689_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n549_), .A2(new_n689_), .A3(new_n626_), .ZN(new_n698_));
  OAI211_X1 g497(.A(KEYINPUT44), .B(new_n688_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n699_), .A2(G29gat), .A3(new_n507_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n688_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n686_), .B1(new_n700_), .B2(new_n703_), .ZN(G1328gat));
  INV_X1    g503(.A(KEYINPUT46), .ZN(new_n705_));
  INV_X1    g504(.A(G36gat), .ZN(new_n706_));
  INV_X1    g505(.A(new_n398_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n699_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n706_), .B1(new_n709_), .B2(new_n703_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n398_), .A2(G36gat), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT45), .B1(new_n684_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n599_), .A2(new_n714_), .A3(new_n683_), .A4(new_n711_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n705_), .B1(new_n710_), .B2(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n703_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G36gat), .B1(new_n719_), .B2(new_n708_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(KEYINPUT46), .A3(new_n716_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n718_), .A2(new_n721_), .ZN(G1329gat));
  XNOR2_X1  g521(.A(KEYINPUT107), .B(G43gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n723_), .B1(new_n684_), .B2(new_n481_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n699_), .A2(G43gat), .A3(new_n518_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n724_), .B1(new_n719_), .B2(new_n725_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g526(.A(G50gat), .B1(new_n685_), .B2(new_n676_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n699_), .A2(G50gat), .A3(new_n676_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n729_), .B2(new_n703_), .ZN(G1331gat));
  INV_X1    g529(.A(new_n594_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n549_), .A2(new_n279_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n643_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n519_), .B1(new_n734_), .B2(KEYINPUT108), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n735_), .B1(KEYINPUT108), .B2(new_n734_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n594_), .A2(new_n642_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n654_), .A2(new_n279_), .A3(new_n737_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n519_), .A2(new_n240_), .ZN(new_n739_));
  AOI22_X1  g538(.A1(new_n736_), .A2(new_n240_), .B1(new_n738_), .B2(new_n739_), .ZN(G1332gat));
  AOI21_X1  g539(.A(new_n238_), .B1(new_n738_), .B2(new_n707_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT48), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n734_), .A2(new_n238_), .A3(new_n707_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n738_), .B2(new_n518_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT49), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n734_), .A2(new_n745_), .A3(new_n518_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1334gat));
  AOI21_X1  g548(.A(new_n441_), .B1(new_n738_), .B2(new_n676_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT50), .Z(new_n751_));
  NAND3_X1  g550(.A1(new_n734_), .A2(new_n441_), .A3(new_n676_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(G1335gat));
  NOR2_X1   g552(.A1(new_n697_), .A2(new_n698_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n276_), .A2(new_n642_), .A3(new_n277_), .A4(new_n731_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT109), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n754_), .A2(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n206_), .B1(new_n758_), .B2(new_n507_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n732_), .A2(new_n683_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n761_), .A2(G85gat), .A3(new_n519_), .ZN(new_n762_));
  OR3_X1    g561(.A1(new_n759_), .A2(new_n760_), .A3(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n760_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(G1336gat));
  INV_X1    g564(.A(new_n761_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(new_n207_), .A3(new_n707_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n754_), .A2(new_n398_), .A3(new_n757_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(new_n207_), .ZN(G1337gat));
  XNOR2_X1  g568(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n518_), .B(new_n756_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(G99gat), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n481_), .A2(new_n204_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n732_), .A2(new_n683_), .A3(new_n777_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT112), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n770_), .B1(new_n776_), .B2(new_n779_), .ZN(new_n780_));
  AND3_X1   g579(.A1(new_n771_), .A2(KEYINPUT111), .A3(G99gat), .ZN(new_n781_));
  AOI21_X1  g580(.A(KEYINPUT111), .B1(new_n771_), .B2(G99gat), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n779_), .B(new_n770_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n780_), .A2(new_n784_), .ZN(G1338gat));
  NAND3_X1  g584(.A1(new_n766_), .A2(new_n219_), .A3(new_n676_), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n676_), .B(new_n756_), .C1(new_n697_), .C2(new_n698_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n787_), .A2(new_n788_), .A3(G106gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n787_), .B2(G106gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT53), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n793_), .B(new_n786_), .C1(new_n789_), .C2(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1339gat));
  NAND3_X1  g594(.A1(new_n625_), .A2(new_n274_), .A3(new_n737_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n796_), .B(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n262_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n262_), .B2(new_n800_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n261_), .B1(new_n253_), .B2(new_n258_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n802_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(KEYINPUT56), .B1(new_n805_), .B2(new_n269_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n262_), .A2(new_n800_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT55), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n262_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n804_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n808_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n270_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n806_), .A2(new_n272_), .A3(new_n594_), .A4(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n572_), .A2(new_n578_), .A3(new_n584_), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n815_), .B(new_n591_), .C1(new_n578_), .C2(new_n581_), .ZN(new_n816_));
  AND2_X1   g615(.A1(new_n593_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n273_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n652_), .B1(new_n814_), .B2(new_n818_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(KEYINPUT57), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n821_), .B(new_n652_), .C1(new_n814_), .C2(new_n818_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n820_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n272_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n811_), .A2(new_n270_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(KEYINPUT56), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n826_), .A2(KEYINPUT116), .A3(new_n817_), .A4(new_n813_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT58), .B1(new_n827_), .B2(KEYINPUT117), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n826_), .A2(new_n817_), .A3(new_n813_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(KEYINPUT117), .A2(KEYINPUT58), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT116), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n626_), .B1(new_n828_), .B2(new_n832_), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n823_), .A2(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n799_), .B1(new_n834_), .B2(new_n648_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT59), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n517_), .A2(new_n519_), .A3(new_n481_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n835_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(KEYINPUT115), .B1(new_n820_), .B2(new_n822_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n819_), .B2(KEYINPUT57), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n841_), .A3(new_n833_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n642_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n799_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n844_), .A2(new_n837_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n838_), .B1(new_n845_), .B2(new_n836_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n594_), .A2(G113gat), .ZN(new_n847_));
  XOR2_X1   g646(.A(new_n847_), .B(KEYINPUT118), .Z(new_n848_));
  NOR2_X1   g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(G113gat), .B1(new_n845_), .B2(new_n594_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1340gat));
  INV_X1    g650(.A(KEYINPUT60), .ZN(new_n852_));
  AOI21_X1  g651(.A(G120gat), .B1(new_n279_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n852_), .B2(G120gat), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n845_), .A2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n855_), .B(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(G120gat), .B1(new_n846_), .B2(new_n278_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(G1341gat));
  NAND2_X1  g658(.A1(new_n648_), .A2(G127gat), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(KEYINPUT120), .Z(new_n861_));
  NOR2_X1   g660(.A1(new_n846_), .A2(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(G127gat), .B1(new_n845_), .B2(new_n648_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n862_), .A2(new_n863_), .ZN(G1342gat));
  OAI21_X1  g663(.A(G134gat), .B1(new_n846_), .B2(new_n625_), .ZN(new_n865_));
  INV_X1    g664(.A(G134gat), .ZN(new_n866_));
  INV_X1    g665(.A(new_n653_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n845_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n865_), .A2(new_n868_), .ZN(G1343gat));
  NOR2_X1   g668(.A1(new_n518_), .A2(new_n455_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n844_), .A2(new_n870_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n871_), .A2(new_n707_), .A3(new_n519_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n594_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n279_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g675(.A1(new_n872_), .A2(new_n648_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT61), .B(G155gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  AOI21_X1  g678(.A(G162gat), .B1(new_n872_), .B2(new_n867_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n693_), .A2(new_n410_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n880_), .B1(new_n872_), .B2(new_n881_), .ZN(G1347gat));
  NOR2_X1   g681(.A1(new_n398_), .A2(new_n520_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n676_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n835_), .A2(new_n885_), .ZN(new_n886_));
  OAI21_X1  g685(.A(G169gat), .B1(new_n886_), .B2(new_n731_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n888_));
  OR2_X1    g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n886_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n890_), .A2(new_n594_), .A3(new_n314_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n887_), .A2(new_n888_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n889_), .A2(new_n891_), .A3(new_n892_), .ZN(G1348gat));
  AOI21_X1  g692(.A(G176gat), .B1(new_n890_), .B2(new_n279_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n798_), .B1(new_n842_), .B2(new_n642_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n676_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n278_), .A2(new_n884_), .A3(new_n315_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n894_), .B1(new_n896_), .B2(new_n897_), .ZN(G1349gat));
  NAND3_X1  g697(.A1(new_n896_), .A2(new_n648_), .A3(new_n883_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n642_), .A2(new_n299_), .ZN(new_n900_));
  AOI22_X1  g699(.A1(new_n899_), .A2(new_n280_), .B1(new_n890_), .B2(new_n900_), .ZN(G1350gat));
  NAND3_X1  g700(.A1(new_n890_), .A2(new_n349_), .A3(new_n867_), .ZN(new_n902_));
  OAI21_X1  g701(.A(G190gat), .B1(new_n886_), .B2(new_n625_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n903_), .A2(KEYINPUT121), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n903_), .A2(KEYINPUT121), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n902_), .B1(new_n904_), .B2(new_n905_), .ZN(G1351gat));
  INV_X1    g705(.A(new_n870_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n398_), .A2(new_n507_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NOR4_X1   g708(.A1(new_n895_), .A2(new_n731_), .A3(new_n907_), .A4(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911_));
  OAI21_X1  g710(.A(KEYINPUT123), .B1(new_n910_), .B2(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G197gat), .B1(new_n910_), .B2(new_n911_), .ZN(new_n913_));
  NAND4_X1  g712(.A1(new_n844_), .A2(new_n594_), .A3(new_n870_), .A4(new_n908_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n914_), .A2(KEYINPUT122), .A3(new_n915_), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n912_), .A2(new_n913_), .A3(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(new_n913_), .B1(new_n916_), .B2(new_n912_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1352gat));
  NOR2_X1   g718(.A1(new_n871_), .A2(new_n909_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n279_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g721(.A1(new_n895_), .A2(new_n907_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n642_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n926_));
  XOR2_X1   g725(.A(new_n926_), .B(KEYINPUT124), .Z(new_n927_));
  NAND4_X1  g726(.A1(new_n923_), .A2(new_n908_), .A3(new_n925_), .A4(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n928_), .A2(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n925_), .B1(new_n920_), .B2(new_n927_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n928_), .A2(new_n929_), .ZN(new_n932_));
  NOR3_X1   g731(.A1(new_n930_), .A2(new_n931_), .A3(new_n932_), .ZN(G1354gat));
  NAND3_X1  g732(.A1(new_n923_), .A2(new_n867_), .A3(new_n908_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(KEYINPUT126), .ZN(new_n935_));
  XOR2_X1   g734(.A(KEYINPUT127), .B(G218gat), .Z(new_n936_));
  NOR2_X1   g735(.A1(new_n625_), .A2(new_n936_), .ZN(new_n937_));
  AOI22_X1  g736(.A1(new_n935_), .A2(new_n936_), .B1(new_n920_), .B2(new_n937_), .ZN(G1355gat));
endmodule


