//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n756_, new_n757_, new_n758_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n867_, new_n868_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n906_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_,
    new_n941_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT23), .ZN(new_n203_));
  NOR2_X1   g002(.A1(G169gat), .A2(G176gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT81), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(new_n203_), .B1(new_n206_), .B2(KEYINPUT24), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G169gat), .A2(G176gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n208_), .B(KEYINPUT82), .Z(new_n209_));
  INV_X1    g008(.A(new_n204_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(new_n205_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n204_), .A2(KEYINPUT81), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n211_), .A2(KEYINPUT24), .A3(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n207_), .B1(new_n209_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT79), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT26), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n215_), .B1(new_n216_), .B2(G190gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT25), .B(G183gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT26), .B(G190gat), .ZN(new_n219_));
  OAI211_X1 g018(.A(new_n217_), .B(new_n218_), .C1(new_n219_), .C2(new_n215_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT80), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n214_), .A2(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(KEYINPUT83), .B(G176gat), .Z(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT22), .B(G169gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n226_), .A2(new_n209_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n203_), .B1(G183gat), .B2(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n223_), .A2(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n230_), .B(KEYINPUT30), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT84), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT87), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G127gat), .B(G134gat), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n236_), .A2(KEYINPUT86), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(KEYINPUT86), .ZN(new_n238_));
  XOR2_X1   g037(.A(G113gat), .B(G120gat), .Z(new_n239_));
  OR3_X1    g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n239_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT31), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n243_), .A2(KEYINPUT85), .ZN(new_n244_));
  INV_X1    g043(.A(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n231_), .A2(new_n232_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G71gat), .B(G99gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(G43gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G227gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n249_), .B(G15gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n248_), .B(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n245_), .B1(new_n246_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n246_), .A2(new_n245_), .A3(new_n251_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n235_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n254_), .ZN(new_n256_));
  NOR3_X1   g055(.A1(new_n256_), .A2(KEYINPUT87), .A3(new_n252_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n234_), .B1(new_n255_), .B2(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT87), .B1(new_n256_), .B2(new_n252_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n253_), .A2(new_n235_), .A3(new_n254_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n259_), .A2(new_n260_), .A3(new_n233_), .ZN(new_n261_));
  AND2_X1   g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G225gat), .A2(G233gat), .ZN(new_n263_));
  NOR2_X1   g062(.A1(G141gat), .A2(G148gat), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT89), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(KEYINPUT3), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT3), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n265_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G141gat), .A2(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT2), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n267_), .A2(new_n269_), .A3(new_n272_), .A4(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(G155gat), .ZN(new_n275_));
  INV_X1    g074(.A(G162gat), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(KEYINPUT88), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT88), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(G155gat), .B2(G162gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G155gat), .A2(G162gat), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(KEYINPUT1), .ZN(new_n283_));
  OR2_X1    g082(.A1(new_n281_), .A2(KEYINPUT1), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n280_), .A2(new_n283_), .A3(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n270_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n286_), .A2(new_n264_), .ZN(new_n287_));
  AOI22_X1  g086(.A1(new_n274_), .A2(new_n282_), .B1(new_n285_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n242_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(KEYINPUT4), .A3(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT4), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n242_), .A2(new_n293_), .A3(new_n289_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n263_), .B1(new_n292_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  XOR2_X1   g095(.A(G1gat), .B(G29gat), .Z(new_n297_));
  XNOR2_X1  g096(.A(G57gat), .B(G85gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n300_));
  XOR2_X1   g099(.A(new_n299_), .B(new_n300_), .Z(new_n301_));
  INV_X1    g100(.A(new_n263_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n296_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n301_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n306_), .B1(new_n295_), .B2(new_n303_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(G197gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT91), .B1(new_n309_), .B2(G204gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT91), .ZN(new_n311_));
  INV_X1    g110(.A(G204gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n311_), .A2(new_n312_), .A3(G197gat), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n309_), .A2(G204gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n310_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT93), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G211gat), .B(G218gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT92), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT21), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n319_), .B1(new_n318_), .B2(new_n317_), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n315_), .A2(KEYINPUT21), .ZN(new_n321_));
  INV_X1    g120(.A(new_n314_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n309_), .A2(G204gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT21), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  AND2_X1   g123(.A1(new_n324_), .A2(new_n317_), .ZN(new_n325_));
  AOI22_X1  g124(.A1(new_n316_), .A2(new_n320_), .B1(new_n321_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n289_), .A2(KEYINPUT29), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(G228gat), .A3(G233gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G228gat), .A2(G233gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(new_n331_), .A3(new_n328_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(KEYINPUT28), .B(G22gat), .Z(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n274_), .A2(new_n282_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n285_), .A2(new_n287_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT29), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT90), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n288_), .A2(KEYINPUT90), .A3(new_n338_), .ZN(new_n342_));
  INV_X1    g141(.A(G50gat), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n343_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n335_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n341_), .A2(new_n342_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(G50gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n341_), .A2(new_n342_), .A3(new_n343_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(new_n334_), .A3(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n333_), .A2(new_n346_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT94), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n346_), .A2(new_n350_), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n330_), .A2(new_n332_), .ZN(new_n355_));
  XOR2_X1   g154(.A(G78gat), .B(G106gat), .Z(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n357_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n353_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n354_), .A2(new_n355_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n356_), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n363_), .A2(new_n352_), .A3(new_n351_), .A4(new_n358_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT19), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n223_), .A2(new_n326_), .A3(new_n229_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n210_), .A2(KEYINPUT24), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n203_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n371_), .B1(new_n213_), .B2(new_n208_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n219_), .B(KEYINPUT95), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n218_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n372_), .A2(new_n374_), .B1(new_n228_), .B2(new_n227_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT20), .B1(new_n375_), .B2(new_n326_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n367_), .B1(new_n369_), .B2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G8gat), .B(G36gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT18), .ZN(new_n379_));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  NAND2_X1  g180(.A1(new_n230_), .A2(new_n327_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n367_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT20), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n384_), .B1(new_n375_), .B2(new_n326_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n382_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n377_), .A2(new_n381_), .A3(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n387_), .A2(KEYINPUT27), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n372_), .A2(new_n374_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(new_n229_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n384_), .B1(new_n390_), .B2(new_n327_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(new_n383_), .A3(new_n368_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n382_), .A2(new_n385_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n392_), .B1(new_n393_), .B2(new_n383_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n381_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n382_), .A2(new_n383_), .A3(new_n385_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n383_), .B1(new_n391_), .B2(new_n368_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n395_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n387_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT99), .B(KEYINPUT27), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  AOI22_X1  g201(.A1(new_n388_), .A2(new_n396_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NOR4_X1   g203(.A1(new_n262_), .A2(new_n308_), .A3(new_n365_), .A4(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n308_), .ZN(new_n406_));
  NOR3_X1   g205(.A1(new_n359_), .A2(new_n353_), .A3(new_n360_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n363_), .A2(new_n358_), .B1(new_n352_), .B2(new_n351_), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n403_), .B(new_n406_), .C1(new_n407_), .C2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT100), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT100), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n365_), .A2(new_n411_), .A3(new_n406_), .A4(new_n403_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n365_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n381_), .A2(KEYINPUT32), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n392_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n383_), .B1(new_n382_), .B2(new_n385_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT98), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT98), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n394_), .A2(new_n420_), .A3(new_n415_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n377_), .A2(new_n386_), .A3(new_n414_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n419_), .A2(new_n421_), .A3(new_n308_), .A4(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT33), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n307_), .A2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n290_), .A2(new_n302_), .A3(new_n291_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n292_), .A2(new_n294_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n301_), .B(new_n426_), .C1(new_n427_), .C2(new_n302_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n425_), .A2(new_n399_), .A3(new_n387_), .A4(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(KEYINPUT33), .B(new_n306_), .C1(new_n295_), .C2(new_n303_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT97), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n423_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n413_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n410_), .A2(new_n412_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n262_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT101), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n434_), .A2(KEYINPUT101), .A3(new_n262_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n405_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT12), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT8), .ZN(new_n441_));
  AND2_X1   g240(.A1(G85gat), .A2(G92gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(G85gat), .A2(G92gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT66), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(G85gat), .ZN(new_n445_));
  INV_X1    g244(.A(G92gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT66), .ZN(new_n448_));
  NAND2_X1  g247(.A1(G85gat), .A2(G92gat), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n444_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G99gat), .A2(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT6), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(G99gat), .A3(G106gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT7), .ZN(new_n458_));
  INV_X1    g257(.A(G99gat), .ZN(new_n459_));
  INV_X1    g258(.A(G106gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n456_), .A2(new_n457_), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n441_), .B1(new_n451_), .B2(new_n462_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n453_), .A2(new_n455_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n457_), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT65), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n444_), .A2(new_n450_), .A3(new_n441_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT65), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n456_), .A2(new_n468_), .A3(new_n457_), .A4(new_n461_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n466_), .A2(new_n467_), .A3(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(KEYINPUT67), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT67), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n466_), .A2(new_n467_), .A3(new_n472_), .A4(new_n469_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n463_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(KEYINPUT10), .B(G99gat), .Z(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n460_), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n476_), .B(KEYINPUT64), .Z(new_n477_));
  NAND3_X1  g276(.A1(new_n447_), .A2(KEYINPUT9), .A3(new_n449_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n478_), .B(new_n456_), .C1(KEYINPUT9), .C2(new_n449_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n474_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G57gat), .B(G64gat), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n482_), .A2(KEYINPUT11), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G71gat), .B(G78gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n483_), .A2(new_n484_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n482_), .A2(KEYINPUT11), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n485_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n440_), .B1(new_n481_), .B2(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(G230gat), .A2(G233gat), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n481_), .B2(new_n488_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n463_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n444_), .A2(new_n450_), .A3(new_n441_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n493_), .B1(KEYINPUT65), .B2(new_n462_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n472_), .B1(new_n494_), .B2(new_n469_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n473_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n492_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT68), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n474_), .A2(KEYINPUT68), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n480_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  OR2_X1    g300(.A1(new_n488_), .A2(new_n440_), .ZN(new_n502_));
  OAI211_X1 g301(.A(new_n489_), .B(new_n491_), .C1(new_n501_), .C2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT69), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n481_), .A2(new_n488_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n481_), .A2(new_n488_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n490_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n474_), .A2(KEYINPUT68), .ZN(new_n510_));
  AOI211_X1 g309(.A(new_n498_), .B(new_n463_), .C1(new_n471_), .C2(new_n473_), .ZN(new_n511_));
  OAI22_X1  g310(.A1(new_n510_), .A2(new_n511_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n502_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n514_), .A2(KEYINPUT69), .A3(new_n489_), .A4(new_n491_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n505_), .A2(new_n509_), .A3(new_n515_), .ZN(new_n516_));
  XOR2_X1   g315(.A(G120gat), .B(G148gat), .Z(new_n517_));
  XNOR2_X1  g316(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G176gat), .B(G204gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n521_), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n505_), .A2(new_n515_), .A3(new_n509_), .A4(new_n523_), .ZN(new_n524_));
  AND3_X1   g323(.A1(new_n522_), .A2(KEYINPUT13), .A3(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(KEYINPUT13), .B1(new_n522_), .B2(new_n524_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(G1gat), .ZN(new_n528_));
  INV_X1    g327(.A(G8gat), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT14), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT76), .Z(new_n531_));
  XNOR2_X1  g330(.A(G15gat), .B(G22gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT75), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G1gat), .B(G8gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  XOR2_X1   g336(.A(G29gat), .B(G36gat), .Z(new_n538_));
  XOR2_X1   g337(.A(G43gat), .B(G50gat), .Z(new_n539_));
  XOR2_X1   g338(.A(new_n538_), .B(new_n539_), .Z(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n540_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n536_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n541_), .A2(new_n543_), .A3(KEYINPUT78), .ZN(new_n544_));
  OR3_X1    g343(.A1(new_n536_), .A2(KEYINPUT78), .A3(new_n542_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n544_), .A2(new_n545_), .A3(G229gat), .A4(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n540_), .B(KEYINPUT15), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n537_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n549_), .A2(new_n550_), .A3(new_n543_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n546_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G113gat), .B(G141gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G169gat), .B(G197gat), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n553_), .B(new_n554_), .Z(new_n555_));
  XOR2_X1   g354(.A(new_n552_), .B(new_n555_), .Z(new_n556_));
  NAND2_X1  g355(.A1(new_n527_), .A2(new_n556_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n439_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(G232gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT34), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(KEYINPUT71), .B(KEYINPUT35), .ZN(new_n562_));
  AOI22_X1  g361(.A1(new_n481_), .A2(new_n542_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n563_), .B1(new_n501_), .B2(new_n547_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n561_), .A2(new_n562_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n512_), .A2(new_n548_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n565_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n568_), .A3(new_n563_), .ZN(new_n569_));
  XNOR2_X1  g368(.A(G190gat), .B(G218gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G134gat), .B(G162gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n572_), .A2(KEYINPUT36), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n566_), .A2(new_n569_), .A3(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT72), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT73), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n566_), .A2(new_n569_), .A3(KEYINPUT72), .A4(new_n573_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n576_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n572_), .B(KEYINPUT36), .Z(new_n580_));
  INV_X1    g379(.A(new_n569_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n568_), .B1(new_n567_), .B2(new_n563_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n580_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n577_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT37), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n576_), .A2(new_n578_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(KEYINPUT74), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT74), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n589_), .B(new_n580_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n587_), .A2(new_n588_), .A3(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n586_), .B1(KEYINPUT37), .B2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n536_), .B(new_n488_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G127gat), .B(G155gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT16), .ZN(new_n597_));
  XOR2_X1   g396(.A(G183gat), .B(G211gat), .Z(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT17), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n599_), .A2(new_n600_), .ZN(new_n602_));
  NOR3_X1   g401(.A1(new_n595_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n603_), .B1(new_n601_), .B2(new_n595_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n592_), .A2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT77), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n558_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT102), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n406_), .A2(G1gat), .ZN(new_n610_));
  AOI21_X1  g409(.A(KEYINPUT38), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  NOR3_X1   g410(.A1(new_n262_), .A2(new_n365_), .A3(new_n404_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(new_n406_), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n434_), .A2(KEYINPUT101), .A3(new_n262_), .ZN(new_n614_));
  AOI21_X1  g413(.A(KEYINPUT101), .B1(new_n434_), .B2(new_n262_), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n613_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n591_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n604_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n617_), .A2(new_n557_), .A3(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n528_), .B1(new_n619_), .B2(new_n308_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n611_), .A2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n609_), .A2(KEYINPUT38), .A3(new_n610_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT103), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n622_), .A2(new_n623_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n621_), .B1(new_n624_), .B2(new_n625_), .ZN(G1324gat));
  NOR2_X1   g425(.A1(new_n403_), .A2(G8gat), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n609_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT39), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n619_), .A2(new_n404_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n629_), .B1(new_n630_), .B2(G8gat), .ZN(new_n631_));
  AOI211_X1 g430(.A(KEYINPUT39), .B(new_n529_), .C1(new_n619_), .C2(new_n404_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n628_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n628_), .B(new_n634_), .C1(new_n631_), .C2(new_n632_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1325gat));
  INV_X1    g437(.A(G15gat), .ZN(new_n639_));
  INV_X1    g438(.A(new_n262_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n619_), .B2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT41), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n639_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n642_), .B1(new_n607_), .B2(new_n643_), .ZN(G1326gat));
  OR3_X1    g443(.A1(new_n607_), .A2(G22gat), .A3(new_n413_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n619_), .A2(new_n365_), .ZN(new_n646_));
  XOR2_X1   g445(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n647_));
  AND3_X1   g446(.A1(new_n646_), .A2(G22gat), .A3(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n647_), .B1(new_n646_), .B2(G22gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(G1327gat));
  NOR2_X1   g449(.A1(new_n591_), .A2(new_n604_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n558_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n308_), .ZN(new_n654_));
  XOR2_X1   g453(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n656_), .B1(new_n439_), .B2(new_n592_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT37), .ZN(new_n658_));
  AND4_X1   g457(.A1(new_n658_), .A2(new_n587_), .A3(new_n588_), .A4(new_n590_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n587_), .A2(KEYINPUT73), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n660_), .A2(new_n579_), .A3(new_n583_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n659_), .B1(KEYINPUT37), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(KEYINPUT106), .A2(KEYINPUT43), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n616_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n657_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n557_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n618_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(KEYINPUT44), .B1(new_n665_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT44), .ZN(new_n670_));
  AOI211_X1 g469(.A(new_n670_), .B(new_n667_), .C1(new_n657_), .C2(new_n664_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n308_), .A2(G29gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n654_), .B1(new_n672_), .B2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(KEYINPUT46), .ZN(new_n675_));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n676_), .B1(new_n672_), .B2(new_n404_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n403_), .A2(G36gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n558_), .A2(new_n651_), .A3(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(KEYINPUT107), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT107), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n558_), .A2(new_n681_), .A3(new_n651_), .A4(new_n678_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT45), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n680_), .A2(KEYINPUT45), .A3(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n675_), .B1(new_n677_), .B2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n665_), .A2(new_n668_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(new_n670_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n665_), .A2(KEYINPUT44), .A3(new_n668_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n404_), .A3(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(G36gat), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n680_), .A2(KEYINPUT45), .A3(new_n682_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT45), .B1(new_n680_), .B2(new_n682_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n693_), .A2(KEYINPUT46), .A3(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n688_), .A2(new_n697_), .ZN(G1329gat));
  NAND4_X1  g497(.A1(new_n690_), .A2(G43gat), .A3(new_n640_), .A4(new_n691_), .ZN(new_n699_));
  INV_X1    g498(.A(G43gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n700_), .B1(new_n652_), .B2(new_n262_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT47), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n699_), .A2(new_n704_), .A3(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1330gat));
  NAND3_X1  g505(.A1(new_n653_), .A2(new_n343_), .A3(new_n365_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n690_), .A2(new_n365_), .A3(new_n691_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(new_n709_), .A3(G50gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G50gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(G1331gat));
  NOR2_X1   g511(.A1(new_n527_), .A2(new_n556_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n604_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n617_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G57gat), .B1(new_n716_), .B2(new_n406_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n616_), .A2(new_n713_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n718_), .A2(new_n606_), .ZN(new_n719_));
  INV_X1    g518(.A(G57gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n308_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n717_), .A2(new_n721_), .ZN(G1332gat));
  INV_X1    g521(.A(G64gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n715_), .B2(new_n404_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT48), .Z(new_n725_));
  NAND3_X1  g524(.A1(new_n719_), .A2(new_n723_), .A3(new_n404_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1333gat));
  INV_X1    g526(.A(G71gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n715_), .B2(new_n640_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT49), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n719_), .A2(new_n728_), .A3(new_n640_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1334gat));
  INV_X1    g531(.A(G78gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n715_), .B2(new_n365_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT50), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n719_), .A2(new_n733_), .A3(new_n365_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1335gat));
  AND2_X1   g536(.A1(new_n718_), .A2(new_n651_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n308_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n713_), .A2(new_n618_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n657_), .B2(new_n664_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n308_), .A2(G85gat), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT109), .Z(new_n743_));
  AOI21_X1  g542(.A(new_n739_), .B1(new_n741_), .B2(new_n743_), .ZN(G1336gat));
  NAND2_X1  g543(.A1(new_n718_), .A2(new_n651_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n446_), .B1(new_n745_), .B2(new_n403_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT110), .ZN(new_n747_));
  OR2_X1    g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n741_), .A2(G92gat), .A3(new_n404_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n746_), .A2(new_n747_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n748_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT111), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n748_), .A2(KEYINPUT111), .A3(new_n749_), .A4(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1337gat));
  NAND2_X1  g554(.A1(new_n741_), .A2(new_n640_), .ZN(new_n756_));
  AND2_X1   g555(.A1(new_n640_), .A2(new_n475_), .ZN(new_n757_));
  AOI22_X1  g556(.A1(new_n756_), .A2(G99gat), .B1(new_n738_), .B2(new_n757_), .ZN(new_n758_));
  XOR2_X1   g557(.A(new_n758_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g558(.A1(new_n738_), .A2(new_n460_), .A3(new_n365_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT52), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n741_), .A2(new_n365_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(G106gat), .ZN(new_n763_));
  AOI211_X1 g562(.A(KEYINPUT52), .B(new_n460_), .C1(new_n741_), .C2(new_n365_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n760_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT53), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n760_), .C1(new_n763_), .C2(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1339gat));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n546_), .A2(new_n551_), .A3(new_n555_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n544_), .A2(new_n545_), .A3(new_n550_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n550_), .B1(new_n536_), .B2(new_n542_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n555_), .B1(new_n549_), .B2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n771_), .A2(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n776_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n503_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n506_), .B(new_n489_), .C1(new_n501_), .C2(new_n502_), .ZN(new_n779_));
  AOI22_X1  g578(.A1(new_n778_), .A2(KEYINPUT55), .B1(new_n490_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n505_), .A2(new_n781_), .A3(new_n515_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(new_n521_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT56), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n523_), .A2(new_n785_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n505_), .A2(new_n781_), .A3(new_n515_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n779_), .A2(new_n490_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n789_), .B1(new_n781_), .B2(new_n503_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n787_), .B1(new_n788_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT113), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n787_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(KEYINPUT113), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n786_), .A2(new_n793_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n556_), .A2(new_n524_), .ZN(new_n798_));
  INV_X1    g597(.A(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n777_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n591_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n770_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n521_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT113), .B1(new_n783_), .B2(new_n787_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n798_), .B1(new_n805_), .B2(new_n796_), .ZN(new_n806_));
  OAI211_X1 g605(.A(KEYINPUT57), .B(new_n591_), .C1(new_n806_), .C2(new_n777_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n523_), .B1(new_n780_), .B2(new_n782_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n791_), .B1(KEYINPUT56), .B2(new_n808_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n524_), .A2(new_n771_), .A3(new_n775_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n809_), .A2(KEYINPUT114), .A3(KEYINPUT58), .A4(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n810_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT58), .B(new_n810_), .C1(new_n803_), .C2(new_n795_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n662_), .A2(new_n811_), .A3(new_n814_), .A4(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n802_), .A2(new_n807_), .A3(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(new_n618_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n525_), .A2(new_n526_), .A3(new_n556_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n592_), .A2(new_n604_), .A3(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n823_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n592_), .A2(new_n604_), .A3(new_n821_), .A4(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n820_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n828_), .A2(new_n308_), .A3(new_n612_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n833_), .A2(KEYINPUT116), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n832_), .B1(new_n829_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n556_), .ZN(new_n836_));
  OAI21_X1  g635(.A(G113gat), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n829_), .B(KEYINPUT115), .ZN(new_n838_));
  INV_X1    g637(.A(G113gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n838_), .A2(new_n839_), .A3(new_n556_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n840_), .ZN(G1340gat));
  INV_X1    g640(.A(G120gat), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(new_n527_), .B2(KEYINPUT60), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n838_), .B(new_n843_), .C1(KEYINPUT60), .C2(new_n842_), .ZN(new_n844_));
  OAI21_X1  g643(.A(G120gat), .B1(new_n835_), .B2(new_n527_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(G1341gat));
  OAI21_X1  g645(.A(G127gat), .B1(new_n835_), .B2(new_n618_), .ZN(new_n847_));
  INV_X1    g646(.A(G127gat), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n838_), .A2(new_n848_), .A3(new_n604_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(G1342gat));
  NAND2_X1  g649(.A1(new_n838_), .A2(new_n801_), .ZN(new_n851_));
  INV_X1    g650(.A(G134gat), .ZN(new_n852_));
  INV_X1    g651(.A(new_n835_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n662_), .A2(G134gat), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT117), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n851_), .A2(new_n852_), .B1(new_n853_), .B2(new_n855_), .ZN(G1343gat));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n413_), .A2(new_n404_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n262_), .A2(new_n308_), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n828_), .A2(new_n857_), .A3(new_n860_), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n819_), .A2(new_n618_), .B1(new_n826_), .B2(new_n824_), .ZN(new_n862_));
  OAI21_X1  g661(.A(KEYINPUT118), .B1(new_n862_), .B2(new_n859_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n556_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g665(.A(new_n527_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n864_), .A2(new_n867_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n864_), .B2(new_n604_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n864_), .A2(new_n870_), .A3(new_n604_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(KEYINPUT61), .B(G155gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n872_), .A2(new_n873_), .A3(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n874_), .ZN(new_n876_));
  AOI211_X1 g675(.A(KEYINPUT119), .B(new_n618_), .C1(new_n861_), .C2(new_n863_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n871_), .B2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n875_), .A2(new_n878_), .ZN(G1346gat));
  AOI21_X1  g678(.A(new_n276_), .B1(new_n864_), .B2(new_n662_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(new_n591_), .A2(G162gat), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT120), .B1(new_n880_), .B2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n864_), .A2(new_n881_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n592_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n885_), .B(new_n886_), .C1(new_n276_), .C2(new_n887_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n884_), .A2(new_n888_), .ZN(G1347gat));
  NOR2_X1   g688(.A1(new_n862_), .A2(new_n365_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n262_), .A2(new_n308_), .A3(new_n403_), .ZN(new_n891_));
  AND3_X1   g690(.A1(new_n890_), .A2(KEYINPUT122), .A3(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(KEYINPUT122), .B1(new_n890_), .B2(new_n891_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n556_), .A3(new_n225_), .ZN(new_n897_));
  INV_X1    g696(.A(G169gat), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n891_), .A2(new_n556_), .ZN(new_n899_));
  XOR2_X1   g698(.A(new_n899_), .B(KEYINPUT121), .Z(new_n900_));
  AOI21_X1  g699(.A(new_n898_), .B1(new_n890_), .B2(new_n900_), .ZN(new_n901_));
  XOR2_X1   g700(.A(new_n901_), .B(KEYINPUT62), .Z(new_n902_));
  NAND2_X1  g701(.A1(new_n897_), .A2(new_n902_), .ZN(G1348gat));
  AND2_X1   g702(.A1(new_n890_), .A2(new_n891_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n904_), .A2(G176gat), .A3(new_n867_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n867_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n905_), .B1(new_n906_), .B2(new_n224_), .ZN(G1349gat));
  AOI21_X1  g706(.A(G183gat), .B1(new_n904_), .B2(new_n604_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n618_), .A2(new_n218_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n908_), .B1(new_n896_), .B2(new_n909_), .ZN(G1350gat));
  OAI211_X1 g709(.A(new_n373_), .B(new_n801_), .C1(new_n892_), .C2(new_n894_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n592_), .B1(new_n893_), .B2(new_n895_), .ZN(new_n912_));
  INV_X1    g711(.A(G190gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(G1351gat));
  INV_X1    g713(.A(KEYINPUT123), .ZN(new_n915_));
  NOR4_X1   g714(.A1(new_n640_), .A2(new_n308_), .A3(new_n413_), .A4(new_n403_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n828_), .A2(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(new_n556_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n915_), .B1(new_n919_), .B2(new_n309_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n919_), .A2(new_n309_), .ZN(new_n921_));
  NAND4_X1  g720(.A1(new_n918_), .A2(KEYINPUT123), .A3(G197gat), .A4(new_n556_), .ZN(new_n922_));
  AND3_X1   g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(G1352gat));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n828_), .A2(new_n867_), .A3(new_n916_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n925_), .B2(G204gat), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT124), .ZN(new_n927_));
  OR2_X1    g726(.A1(new_n925_), .A2(new_n927_), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n312_), .B1(new_n925_), .B2(new_n927_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n926_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n930_));
  AND2_X1   g729(.A1(new_n928_), .A2(new_n929_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n930_), .B1(KEYINPUT125), .B2(new_n931_), .ZN(G1353gat));
  NOR2_X1   g731(.A1(new_n917_), .A2(new_n618_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n934_));
  AND2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n933_), .B1(new_n934_), .B2(new_n935_), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(new_n933_), .B2(new_n934_), .ZN(G1354gat));
  OR3_X1    g736(.A1(new_n917_), .A2(G218gat), .A3(new_n591_), .ZN(new_n938_));
  OAI21_X1  g737(.A(G218gat), .B1(new_n917_), .B2(new_n592_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n940_), .B(new_n941_), .ZN(G1355gat));
endmodule


