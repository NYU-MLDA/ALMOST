//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n839_, new_n840_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT36), .Z(new_n205_));
  NAND2_X1  g004(.A1(G232gat), .A2(G233gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n206_), .B(KEYINPUT34), .Z(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT70), .B(KEYINPUT35), .Z(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT7), .ZN(new_n211_));
  INV_X1    g010(.A(G99gat), .ZN(new_n212_));
  INV_X1    g011(.A(G106gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT66), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT6), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G99gat), .A3(G106gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222_));
  NAND4_X1  g021(.A1(new_n222_), .A2(new_n211_), .A3(new_n212_), .A4(new_n213_), .ZN(new_n223_));
  NAND4_X1  g022(.A1(new_n215_), .A2(new_n220_), .A3(new_n221_), .A4(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G85gat), .ZN(new_n225_));
  INV_X1    g024(.A(G92gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G85gat), .A2(G92gat), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n224_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT8), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n224_), .A2(KEYINPUT8), .A3(new_n229_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT10), .B(G99gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT65), .B1(new_n234_), .B2(G106gat), .ZN(new_n235_));
  OR2_X1    g034(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n237_));
  NAND2_X1  g036(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n236_), .A2(new_n237_), .A3(new_n213_), .A4(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n235_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n227_), .A2(KEYINPUT9), .A3(new_n228_), .ZN(new_n241_));
  OR2_X1    g040(.A1(new_n228_), .A2(KEYINPUT9), .ZN(new_n242_));
  AND3_X1   g041(.A1(new_n220_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n232_), .A2(new_n233_), .A3(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G29gat), .B(G36gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G43gat), .B(G50gat), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n247_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n249_), .A2(KEYINPUT15), .A3(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT15), .ZN(new_n252_));
  INV_X1    g051(.A(new_n250_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n252_), .B1(new_n253_), .B2(new_n248_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n245_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT71), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n245_), .A2(KEYINPUT71), .A3(new_n255_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n253_), .A2(new_n248_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n232_), .A2(new_n262_), .A3(new_n233_), .A4(new_n244_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n207_), .A2(new_n208_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT72), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n210_), .B1(new_n260_), .B2(new_n267_), .ZN(new_n268_));
  AOI211_X1 g067(.A(new_n209_), .B(new_n266_), .C1(new_n258_), .C2(new_n259_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n205_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n259_), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT71), .B1(new_n245_), .B2(new_n255_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n267_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n209_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n260_), .A2(new_n210_), .A3(new_n267_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n270_), .A2(KEYINPUT74), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT73), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT73), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n270_), .A2(new_n280_), .A3(new_n277_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n279_), .A2(KEYINPUT37), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT37), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n278_), .A2(KEYINPUT73), .A3(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n282_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G15gat), .B(G22gat), .ZN(new_n287_));
  INV_X1    g086(.A(G1gat), .ZN(new_n288_));
  INV_X1    g087(.A(G8gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT14), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G1gat), .B(G8gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G57gat), .B(G64gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G71gat), .B(G78gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(new_n295_), .A3(KEYINPUT11), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(KEYINPUT11), .ZN(new_n297_));
  INV_X1    g096(.A(new_n295_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n294_), .A2(KEYINPUT11), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n296_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n293_), .B(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(G231gat), .ZN(new_n303_));
  INV_X1    g102(.A(G233gat), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G127gat), .B(G155gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT16), .ZN(new_n309_));
  XOR2_X1   g108(.A(G183gat), .B(G211gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(new_n309_), .B(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT17), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n302_), .A2(new_n306_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n307_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n311_), .B(new_n312_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n317_), .B1(new_n307_), .B2(new_n314_), .ZN(new_n318_));
  OAI21_X1  g117(.A(KEYINPUT75), .B1(new_n316_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n320_));
  AND2_X1   g119(.A1(new_n307_), .A2(new_n314_), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n320_), .B(new_n315_), .C1(new_n321_), .C2(new_n317_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n319_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n286_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G120gat), .B(G148gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G176gat), .B(G204gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n232_), .A2(new_n233_), .A3(new_n244_), .A4(new_n301_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G230gat), .A2(G233gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n332_), .B(KEYINPUT64), .Z(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n230_), .A2(new_n231_), .B1(new_n240_), .B2(new_n243_), .ZN(new_n336_));
  AOI211_X1 g135(.A(KEYINPUT12), .B(new_n301_), .C1(new_n336_), .C2(new_n233_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT12), .ZN(new_n338_));
  INV_X1    g137(.A(new_n301_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n338_), .B1(new_n245_), .B2(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n335_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n245_), .A2(new_n339_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n334_), .B1(new_n343_), .B2(new_n331_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n330_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n344_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n330_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n341_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT68), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n349_), .B1(new_n350_), .B2(KEYINPUT13), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n350_), .A2(KEYINPUT13), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n350_), .A2(KEYINPUT13), .ZN(new_n353_));
  OAI211_X1 g152(.A(new_n345_), .B(new_n348_), .C1(new_n352_), .C2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n351_), .A2(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n355_), .A2(KEYINPUT69), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(KEYINPUT69), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n325_), .A2(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G127gat), .B(G134gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G113gat), .B(G120gat), .ZN(new_n361_));
  OR2_X1    g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT82), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n361_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n360_), .A2(new_n361_), .A3(KEYINPUT82), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n365_), .A2(new_n366_), .ZN(new_n367_));
  XOR2_X1   g166(.A(new_n367_), .B(KEYINPUT31), .Z(new_n368_));
  NAND2_X1  g167(.A1(G227gat), .A2(G233gat), .ZN(new_n369_));
  XOR2_X1   g168(.A(new_n369_), .B(G15gat), .Z(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(KEYINPUT30), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(KEYINPUT23), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT23), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(G183gat), .A3(G190gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(G169gat), .A2(G176gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT79), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n377_), .B1(new_n382_), .B2(KEYINPUT24), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT80), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n380_), .A2(new_n381_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n385_), .A2(new_n386_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT80), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(KEYINPUT25), .B(G183gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(KEYINPUT26), .B(G190gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(G169gat), .ZN(new_n393_));
  INV_X1    g192(.A(G176gat), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n382_), .B(KEYINPUT24), .C1(new_n393_), .C2(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n384_), .A2(new_n389_), .A3(new_n392_), .A4(new_n395_), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G183gat), .A2(G190gat), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n375_), .B2(new_n373_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(new_n375_), .B2(new_n373_), .ZN(new_n399_));
  OAI21_X1  g198(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n400_));
  OR3_X1    g199(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n399_), .A2(new_n400_), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n396_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G71gat), .B(G99gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT81), .B(G43gat), .ZN(new_n405_));
  XOR2_X1   g204(.A(new_n404_), .B(new_n405_), .Z(new_n406_));
  AND2_X1   g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n403_), .A2(new_n406_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n372_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n403_), .A2(new_n406_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n403_), .A2(new_n406_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n371_), .A3(new_n411_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n409_), .A2(new_n412_), .A3(KEYINPUT83), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT83), .B1(new_n409_), .B2(new_n412_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n368_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n409_), .A2(new_n412_), .A3(KEYINPUT83), .ZN(new_n416_));
  INV_X1    g215(.A(new_n368_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n415_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT27), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G226gat), .A2(G233gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT19), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n424_));
  XOR2_X1   g223(.A(G211gat), .B(G218gat), .Z(new_n425_));
  XOR2_X1   g224(.A(G197gat), .B(G204gat), .Z(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT21), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n425_), .B1(new_n427_), .B2(KEYINPUT87), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G197gat), .B(G204gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT21), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  OR2_X1    g230(.A1(new_n431_), .A2(KEYINPUT88), .ZN(new_n432_));
  OR3_X1    g231(.A1(new_n429_), .A2(KEYINPUT87), .A3(new_n430_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(KEYINPUT88), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n428_), .A2(new_n432_), .A3(new_n433_), .A4(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT89), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n427_), .B1(new_n436_), .B2(new_n425_), .ZN(new_n437_));
  OR2_X1    g236(.A1(new_n425_), .A2(new_n436_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n437_), .A2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n435_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n395_), .A2(new_n387_), .A3(new_n392_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(new_n402_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n424_), .B1(new_n440_), .B2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n396_), .A2(new_n439_), .A3(new_n435_), .A4(new_n402_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n423_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G8gat), .B(G36gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT18), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G64gat), .B(G92gat), .ZN(new_n449_));
  XOR2_X1   g248(.A(new_n448_), .B(new_n449_), .Z(new_n450_));
  AND2_X1   g249(.A1(new_n435_), .A2(new_n439_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n442_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n424_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n403_), .A2(new_n440_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n453_), .A2(new_n423_), .A3(new_n454_), .ZN(new_n455_));
  AND3_X1   g254(.A1(new_n446_), .A2(new_n450_), .A3(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n450_), .B1(new_n446_), .B2(new_n455_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n420_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(G155gat), .A2(G162gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(G155gat), .A2(G162gat), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n462_));
  INV_X1    g261(.A(G141gat), .ZN(new_n463_));
  INV_X1    g262(.A(G148gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  OAI22_X1  g264(.A1(KEYINPUT84), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT2), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G141gat), .A2(G148gat), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n465_), .B(new_n466_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT85), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n459_), .B(new_n461_), .C1(new_n469_), .C2(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n460_), .B1(KEYINPUT1), .B2(new_n459_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(KEYINPUT1), .B2(new_n459_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n463_), .A2(new_n464_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(new_n476_), .A3(new_n468_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n367_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n362_), .A2(new_n364_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n473_), .A2(new_n477_), .A3(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G225gat), .A2(G233gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n479_), .A2(KEYINPUT4), .A3(new_n481_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n483_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT4), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n478_), .A2(new_n487_), .A3(new_n367_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n485_), .A2(new_n486_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n484_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G29gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G57gat), .B(G85gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n490_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT95), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n484_), .A2(new_n489_), .A3(new_n495_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n497_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n490_), .A2(KEYINPUT95), .A3(new_n496_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n446_), .A2(new_n455_), .A3(new_n450_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n423_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n504_));
  AND3_X1   g303(.A1(new_n443_), .A2(new_n423_), .A3(new_n444_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(KEYINPUT27), .B(new_n503_), .C1(new_n506_), .C2(new_n450_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n458_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G78gat), .B(G106gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(G22gat), .B(G50gat), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT28), .ZN(new_n511_));
  INV_X1    g310(.A(new_n478_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT29), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n511_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NOR3_X1   g313(.A1(new_n478_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n510_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n514_), .A2(new_n515_), .A3(new_n510_), .ZN(new_n518_));
  OAI211_X1 g317(.A(KEYINPUT90), .B(new_n509_), .C1(new_n517_), .C2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n518_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n509_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(new_n516_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n440_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n524_));
  AND2_X1   g323(.A1(new_n304_), .A2(KEYINPUT86), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n304_), .A2(KEYINPUT86), .ZN(new_n526_));
  OAI21_X1  g325(.A(G228gat), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n524_), .B(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n528_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n519_), .A2(new_n530_), .A3(new_n522_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n419_), .B1(new_n508_), .B2(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n485_), .A2(new_n483_), .A3(new_n488_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT94), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n495_), .B1(new_n482_), .B2(new_n486_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n485_), .A2(new_n537_), .A3(new_n483_), .A4(new_n488_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n535_), .A2(new_n536_), .A3(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n484_), .A2(new_n489_), .A3(KEYINPUT33), .A4(new_n495_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n541_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT92), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT33), .B1(new_n499_), .B2(new_n543_), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n484_), .A2(new_n489_), .A3(KEYINPUT92), .A4(new_n495_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT93), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT93), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n544_), .A2(new_n548_), .A3(new_n545_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n542_), .A2(new_n547_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n531_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n530_), .B1(new_n519_), .B2(new_n522_), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n450_), .A2(KEYINPUT32), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n506_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n446_), .A2(new_n455_), .A3(new_n554_), .ZN(new_n556_));
  NAND4_X1  g355(.A1(new_n555_), .A2(new_n501_), .A3(new_n500_), .A4(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n550_), .A2(new_n553_), .A3(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n415_), .A2(new_n418_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n502_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n458_), .A2(new_n507_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n532_), .A2(new_n562_), .ZN(new_n563_));
  AOI22_X1  g362(.A1(new_n533_), .A2(new_n558_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n293_), .B(new_n261_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n255_), .A2(new_n293_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n293_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n567_), .B1(new_n570_), .B2(new_n262_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n568_), .A2(new_n572_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G113gat), .B(G141gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT77), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G169gat), .B(G197gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(KEYINPUT78), .B1(new_n573_), .B2(new_n578_), .ZN(new_n579_));
  AOI22_X1  g378(.A1(new_n565_), .A2(new_n567_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT78), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n580_), .A2(new_n581_), .A3(new_n577_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n573_), .A2(KEYINPUT76), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT76), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n584_), .A2(new_n586_), .A3(new_n578_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n564_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n359_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n592_), .A2(KEYINPUT96), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(KEYINPUT96), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n502_), .A2(G1gat), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n593_), .A2(KEYINPUT38), .A3(new_n594_), .A4(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT97), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n358_), .A2(new_n589_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n316_), .A2(new_n318_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(KEYINPUT98), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n274_), .A2(new_n275_), .A3(new_n276_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n205_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n603_), .A2(new_n605_), .A3(KEYINPUT99), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT99), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n270_), .B2(new_n277_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n564_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT98), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n599_), .A2(new_n611_), .A3(new_n600_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n602_), .A2(new_n610_), .A3(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G1gat), .B1(new_n613_), .B2(new_n502_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT100), .Z(new_n615_));
  NAND3_X1  g414(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT38), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT101), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n616_), .A2(KEYINPUT101), .A3(new_n617_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n598_), .B(new_n615_), .C1(new_n618_), .C2(new_n619_), .ZN(G1324gat));
  NAND4_X1  g419(.A1(new_n593_), .A2(new_n289_), .A3(new_n562_), .A4(new_n594_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n622_));
  INV_X1    g421(.A(new_n562_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G8gat), .B1(new_n613_), .B2(new_n623_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n624_), .A2(KEYINPUT39), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n624_), .A2(KEYINPUT39), .ZN(new_n626_));
  OAI211_X1 g425(.A(new_n621_), .B(new_n622_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n624_), .B(KEYINPUT39), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n622_), .B1(new_n629_), .B2(new_n621_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n628_), .A2(new_n630_), .ZN(G1325gat));
  OR2_X1    g430(.A1(new_n613_), .A2(new_n559_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(G15gat), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT41), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT41), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n632_), .A2(new_n635_), .A3(G15gat), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(KEYINPUT103), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n634_), .A2(new_n639_), .A3(new_n636_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n591_), .A2(G15gat), .A3(new_n559_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT104), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n638_), .A2(new_n640_), .A3(new_n642_), .ZN(G1326gat));
  OAI21_X1  g442(.A(G22gat), .B1(new_n613_), .B2(new_n553_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT42), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n553_), .A2(G22gat), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n645_), .B1(new_n591_), .B2(new_n646_), .ZN(G1327gat));
  INV_X1    g446(.A(new_n358_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n590_), .A2(new_n648_), .A3(new_n323_), .A4(new_n609_), .ZN(new_n649_));
  OR3_X1    g448(.A1(new_n649_), .A2(G29gat), .A3(new_n502_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n558_), .A2(new_n533_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n561_), .A2(new_n563_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(new_n285_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n324_), .B1(new_n654_), .B2(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n653_), .A2(KEYINPUT43), .A3(new_n285_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n656_), .A2(KEYINPUT44), .A3(new_n599_), .A4(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n655_), .B1(new_n564_), .B2(new_n286_), .ZN(new_n659_));
  NAND4_X1  g458(.A1(new_n659_), .A2(new_n657_), .A3(new_n323_), .A4(new_n599_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT44), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n658_), .A2(new_n662_), .A3(new_n560_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT105), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(G29gat), .B1(new_n663_), .B2(new_n664_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n650_), .B1(new_n665_), .B2(new_n666_), .ZN(G1328gat));
  OR2_X1    g466(.A1(new_n623_), .A2(KEYINPUT107), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n623_), .A2(KEYINPUT107), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n649_), .A2(G36gat), .A3(new_n671_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT45), .Z(new_n673_));
  NAND3_X1  g472(.A1(new_n658_), .A2(new_n662_), .A3(new_n562_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n674_), .A2(KEYINPUT106), .A3(G36gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT106), .B1(new_n674_), .B2(G36gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n673_), .B1(new_n675_), .B2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n673_), .B(KEYINPUT46), .C1(new_n675_), .C2(new_n676_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1329gat));
  NAND2_X1  g480(.A1(new_n658_), .A2(new_n662_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G43gat), .B1(new_n682_), .B2(new_n559_), .ZN(new_n683_));
  OR3_X1    g482(.A1(new_n649_), .A2(G43gat), .A3(new_n559_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  XOR2_X1   g484(.A(new_n685_), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g485(.A(G50gat), .B1(new_n682_), .B2(new_n553_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n553_), .A2(G50gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT108), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n687_), .B1(new_n649_), .B2(new_n689_), .ZN(G1331gat));
  NAND4_X1  g489(.A1(new_n610_), .A2(new_n589_), .A3(new_n358_), .A4(new_n324_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n691_), .A2(KEYINPUT109), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(KEYINPUT109), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n692_), .A2(new_n560_), .A3(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(G57gat), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n564_), .A2(new_n588_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n325_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n696_), .A2(new_n358_), .A3(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n560_), .A2(new_n695_), .ZN(new_n699_));
  OAI22_X1  g498(.A1(new_n694_), .A2(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(G1332gat));
  OR3_X1    g499(.A1(new_n698_), .A2(G64gat), .A3(new_n671_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n692_), .A2(new_n670_), .A3(new_n693_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT48), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n702_), .A2(new_n703_), .A3(G64gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n702_), .B2(G64gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(G1333gat));
  OR3_X1    g505(.A1(new_n698_), .A2(G71gat), .A3(new_n559_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n692_), .A2(new_n419_), .A3(new_n693_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT110), .B(KEYINPUT49), .ZN(new_n709_));
  AND3_X1   g508(.A1(new_n708_), .A2(G71gat), .A3(new_n709_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n708_), .B2(G71gat), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n707_), .B1(new_n710_), .B2(new_n711_), .ZN(G1334gat));
  OR3_X1    g511(.A1(new_n698_), .A2(G78gat), .A3(new_n553_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n692_), .A2(new_n532_), .A3(new_n693_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT50), .ZN(new_n715_));
  AND3_X1   g514(.A1(new_n714_), .A2(new_n715_), .A3(G78gat), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n714_), .B2(G78gat), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n713_), .B1(new_n716_), .B2(new_n717_), .ZN(G1335gat));
  NAND4_X1  g517(.A1(new_n656_), .A2(new_n589_), .A3(new_n358_), .A4(new_n657_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G85gat), .B1(new_n719_), .B2(new_n502_), .ZN(new_n720_));
  NAND4_X1  g519(.A1(new_n696_), .A2(new_n358_), .A3(new_n323_), .A4(new_n609_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n722_), .A2(new_n225_), .A3(new_n560_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n720_), .A2(new_n723_), .ZN(G1336gat));
  OAI21_X1  g523(.A(G92gat), .B1(new_n719_), .B2(new_n671_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n722_), .A2(new_n226_), .A3(new_n562_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1337gat));
  OAI21_X1  g526(.A(G99gat), .B1(new_n719_), .B2(new_n559_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n559_), .A2(new_n234_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT111), .B1(new_n722_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g531(.A(G106gat), .B1(new_n719_), .B2(new_n553_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT112), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n735_), .B(G106gat), .C1(new_n719_), .C2(new_n553_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n734_), .A2(KEYINPUT52), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT52), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n733_), .A2(KEYINPUT112), .A3(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n722_), .A2(new_n213_), .A3(new_n532_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(KEYINPUT53), .B1(new_n737_), .B2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n734_), .A2(KEYINPUT52), .A3(new_n736_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT53), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(new_n739_), .A4(new_n740_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n742_), .A2(new_n745_), .ZN(G1339gat));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n569_), .B(new_n567_), .C1(new_n261_), .C2(new_n293_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n577_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n573_), .A2(KEYINPUT78), .A3(new_n578_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n581_), .B1(new_n580_), .B2(new_n577_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n750_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n345_), .B2(new_n348_), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n331_), .B1(new_n337_), .B2(new_n340_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n333_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n341_), .A2(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(KEYINPUT55), .B(new_n335_), .C1(new_n337_), .C2(new_n340_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n756_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT56), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n347_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  AOI22_X1  g562(.A1(new_n333_), .A2(new_n755_), .B1(new_n341_), .B2(new_n757_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n347_), .B1(new_n764_), .B2(new_n759_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n763_), .B1(new_n765_), .B2(KEYINPUT56), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n588_), .A2(new_n348_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n754_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n747_), .B1(new_n768_), .B2(new_n609_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT57), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT99), .B1(new_n603_), .B2(new_n605_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n270_), .A2(new_n607_), .A3(new_n277_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n588_), .A2(new_n348_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n760_), .A2(new_n330_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n761_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n774_), .B1(new_n776_), .B2(new_n763_), .ZN(new_n777_));
  OAI211_X1 g576(.A(KEYINPUT114), .B(new_n773_), .C1(new_n777_), .C2(new_n754_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n769_), .A2(new_n770_), .A3(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT57), .B1(new_n606_), .B2(new_n608_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT116), .B1(new_n768_), .B2(new_n780_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n782_), .B(new_n783_), .C1(new_n777_), .C2(new_n754_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT58), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n760_), .A2(KEYINPUT115), .A3(new_n762_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT56), .B1(new_n760_), .B2(new_n330_), .ZN(new_n789_));
  AOI21_X1  g588(.A(KEYINPUT115), .B1(new_n760_), .B2(new_n762_), .ZN(new_n790_));
  NOR3_X1   g589(.A1(new_n788_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n753_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n348_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n786_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT115), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n763_), .A2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n776_), .A2(new_n796_), .A3(new_n787_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n793_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n797_), .A2(KEYINPUT58), .A3(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n794_), .A2(new_n285_), .A3(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n779_), .A2(new_n785_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n323_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT117), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n319_), .A2(new_n322_), .A3(new_n583_), .A4(new_n587_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n351_), .B2(new_n354_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n282_), .A2(new_n805_), .A3(new_n284_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT54), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n806_), .B(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n801_), .A2(new_n810_), .A3(new_n323_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n803_), .A2(new_n809_), .A3(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  NOR4_X1   g612(.A1(new_n559_), .A2(new_n532_), .A3(new_n562_), .A4(new_n502_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT59), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n600_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n801_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n809_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n819_), .A2(new_n814_), .ZN(new_n820_));
  OAI22_X1  g619(.A1(new_n813_), .A2(new_n816_), .B1(new_n820_), .B2(new_n815_), .ZN(new_n821_));
  OAI21_X1  g620(.A(G113gat), .B1(new_n821_), .B2(new_n589_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n819_), .A2(new_n814_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n823_), .A2(G113gat), .A3(new_n589_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n822_), .A2(KEYINPUT118), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827_));
  INV_X1    g626(.A(G113gat), .ZN(new_n828_));
  INV_X1    g627(.A(new_n816_), .ZN(new_n829_));
  AOI22_X1  g628(.A1(new_n812_), .A2(new_n829_), .B1(new_n823_), .B2(KEYINPUT59), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n828_), .B1(new_n830_), .B2(new_n588_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n827_), .B1(new_n831_), .B2(new_n824_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n826_), .A2(new_n832_), .ZN(G1340gat));
  XNOR2_X1  g632(.A(KEYINPUT119), .B(G120gat), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n358_), .A2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n820_), .B1(KEYINPUT60), .B2(new_n835_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n830_), .A2(new_n836_), .A3(new_n358_), .ZN(new_n837_));
  OAI22_X1  g636(.A1(new_n837_), .A2(new_n834_), .B1(KEYINPUT60), .B2(new_n836_), .ZN(G1341gat));
  OAI21_X1  g637(.A(G127gat), .B1(new_n821_), .B2(new_n817_), .ZN(new_n839_));
  OR3_X1    g638(.A1(new_n823_), .A2(G127gat), .A3(new_n323_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1342gat));
  OAI21_X1  g640(.A(G134gat), .B1(new_n821_), .B2(new_n286_), .ZN(new_n842_));
  OR3_X1    g641(.A1(new_n823_), .A2(G134gat), .A3(new_n773_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1343gat));
  NOR2_X1   g643(.A1(new_n553_), .A2(new_n419_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n670_), .A2(new_n502_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n797_), .A2(new_n798_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n847_), .A2(new_n786_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n848_));
  AOI22_X1  g647(.A1(new_n848_), .A2(new_n799_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n600_), .B1(new_n849_), .B2(new_n779_), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n845_), .B(new_n846_), .C1(new_n850_), .C2(new_n808_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(KEYINPUT120), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT120), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n819_), .A2(new_n853_), .A3(new_n845_), .A4(new_n846_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(new_n588_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n358_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n855_), .B2(new_n324_), .ZN(new_n861_));
  AOI211_X1 g660(.A(KEYINPUT121), .B(new_n323_), .C1(new_n852_), .C2(new_n854_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT61), .B(G155gat), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n861_), .A2(new_n862_), .A3(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n845_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n866_), .B1(new_n818_), .B2(new_n809_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n853_), .B1(new_n867_), .B2(new_n846_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n808_), .B1(new_n801_), .B2(new_n817_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n846_), .ZN(new_n870_));
  NOR4_X1   g669(.A1(new_n869_), .A2(KEYINPUT120), .A3(new_n866_), .A4(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n324_), .B1(new_n868_), .B2(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(KEYINPUT121), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n855_), .A2(new_n860_), .A3(new_n324_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n863_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n865_), .A2(new_n875_), .ZN(G1346gat));
  AOI21_X1  g675(.A(G162gat), .B1(new_n855_), .B2(new_n609_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n285_), .A2(G162gat), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n878_), .B(KEYINPUT122), .Z(new_n879_));
  AOI21_X1  g678(.A(new_n877_), .B1(new_n855_), .B2(new_n879_), .ZN(G1347gat));
  NOR2_X1   g679(.A1(new_n671_), .A2(new_n560_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n419_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n553_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n884_), .A2(new_n589_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n393_), .B1(new_n885_), .B2(new_n812_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887_));
  OR3_X1    g686(.A1(new_n886_), .A2(new_n887_), .A3(KEYINPUT62), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT22), .B(G169gat), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n885_), .A2(new_n812_), .A3(new_n889_), .ZN(new_n890_));
  AND2_X1   g689(.A1(new_n886_), .A2(new_n887_), .ZN(new_n891_));
  OAI21_X1  g690(.A(KEYINPUT62), .B1(new_n886_), .B2(new_n887_), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n888_), .B(new_n890_), .C1(new_n891_), .C2(new_n892_), .ZN(G1348gat));
  NAND3_X1  g692(.A1(new_n812_), .A2(new_n553_), .A3(new_n883_), .ZN(new_n894_));
  INV_X1    g693(.A(new_n894_), .ZN(new_n895_));
  AOI21_X1  g694(.A(G176gat), .B1(new_n895_), .B2(new_n358_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n869_), .A2(new_n532_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(KEYINPUT124), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n882_), .A2(new_n394_), .A3(new_n648_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n896_), .B1(new_n898_), .B2(new_n899_), .ZN(G1349gat));
  NOR3_X1   g699(.A1(new_n894_), .A2(new_n390_), .A3(new_n817_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n898_), .A2(new_n324_), .A3(new_n883_), .ZN(new_n902_));
  INV_X1    g701(.A(G183gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(G1350gat));
  OAI21_X1  g703(.A(G190gat), .B1(new_n894_), .B2(new_n286_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n609_), .A2(new_n391_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n905_), .B1(new_n894_), .B2(new_n906_), .ZN(G1351gat));
  INV_X1    g706(.A(G197gat), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n867_), .A2(new_n881_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n909_), .B2(new_n589_), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n911_));
  NAND4_X1  g710(.A1(new_n867_), .A2(G197gat), .A3(new_n588_), .A4(new_n881_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n913_), .B1(new_n911_), .B2(new_n912_), .ZN(G1352gat));
  INV_X1    g713(.A(G204gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n358_), .B1(KEYINPUT126), .B2(new_n915_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n909_), .A2(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(KEYINPUT126), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n917_), .B(new_n918_), .Z(G1353gat));
  NAND2_X1  g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n600_), .A2(new_n920_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(KEYINPUT127), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n909_), .A2(new_n922_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1354gat));
  OAI21_X1  g724(.A(G218gat), .B1(new_n909_), .B2(new_n286_), .ZN(new_n926_));
  OR2_X1    g725(.A1(new_n773_), .A2(G218gat), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n909_), .B2(new_n927_), .ZN(G1355gat));
endmodule


