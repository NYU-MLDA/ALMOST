//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n618_, new_n619_, new_n620_, new_n622_, new_n623_, new_n624_,
    new_n625_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n705_, new_n706_, new_n707_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n830_, new_n831_, new_n832_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT6), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT6), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G99gat), .A3(G106gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n203_), .A2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT10), .B(G99gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(new_n207_), .B2(G106gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT65), .ZN(new_n210_));
  OR2_X1    g009(.A1(G85gat), .A2(G92gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT64), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G85gat), .A2(G92gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT9), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  AND2_X1   g015(.A1(G85gat), .A2(G92gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n219_), .A2(new_n212_), .A3(KEYINPUT9), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n210_), .B1(new_n221_), .B2(new_n211_), .ZN(new_n222_));
  AOI211_X1 g021(.A(KEYINPUT65), .B(new_n218_), .C1(new_n216_), .C2(new_n220_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n209_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT7), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  OAI211_X1 g029(.A(KEYINPUT66), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n206_), .A2(new_n227_), .A3(new_n230_), .A4(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT67), .B(KEYINPUT8), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n232_), .A2(new_n219_), .A3(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT68), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n219_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT8), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n232_), .A2(new_n238_), .A3(new_n219_), .A4(new_n233_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n235_), .A2(new_n237_), .A3(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n224_), .A2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT69), .B(G71gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G78gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G57gat), .B(G64gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT11), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n244_), .A2(KEYINPUT11), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n243_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(G78gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n242_), .B(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(new_n245_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n241_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT12), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(KEYINPUT71), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT71), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n252_), .B1(new_n224_), .B2(new_n240_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(KEYINPUT12), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n256_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n224_), .A2(new_n252_), .A3(new_n240_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n219_), .ZN(new_n263_));
  AND2_X1   g062(.A1(new_n230_), .A2(new_n231_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n203_), .A2(new_n205_), .B1(new_n226_), .B2(new_n225_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT8), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n239_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n238_), .B1(new_n266_), .B2(new_n233_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT70), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT70), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n235_), .A2(new_n237_), .A3(new_n271_), .A4(new_n239_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n224_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n252_), .A2(new_n255_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n262_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(G230gat), .A2(G233gat), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n260_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n277_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(new_n262_), .B2(new_n258_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  XOR2_X1   g080(.A(G120gat), .B(G148gat), .Z(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT5), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G176gat), .B(G204gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n281_), .A2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n281_), .A2(new_n285_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT13), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n286_), .A2(KEYINPUT13), .A3(new_n287_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G29gat), .B(G36gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G43gat), .B(G50gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n294_), .B(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT74), .B(KEYINPUT15), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G15gat), .B(G22gat), .ZN(new_n299_));
  INV_X1    g098(.A(G1gat), .ZN(new_n300_));
  INV_X1    g099(.A(G8gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT14), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G1gat), .B(G8gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n298_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n305_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n296_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G229gat), .A2(G233gat), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n309_), .B(KEYINPUT81), .Z(new_n310_));
  NAND3_X1  g109(.A1(new_n306_), .A2(new_n308_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n296_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n305_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n308_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n311_), .B1(new_n315_), .B2(new_n309_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G113gat), .B(G141gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G169gat), .B(G197gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n317_), .B(new_n318_), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n316_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT82), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n293_), .A2(KEYINPUT106), .A3(new_n322_), .ZN(new_n323_));
  XOR2_X1   g122(.A(G127gat), .B(G155gat), .Z(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT16), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G183gat), .B(G211gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT17), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G231gat), .A2(G233gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n305_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(new_n252_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT80), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n329_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n334_), .B1(new_n333_), .B2(new_n332_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n332_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT79), .B1(new_n327_), .B2(new_n328_), .ZN(new_n337_));
  OR3_X1    g136(.A1(new_n327_), .A2(KEYINPUT79), .A3(new_n328_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n336_), .A2(new_n337_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT106), .ZN(new_n342_));
  INV_X1    g141(.A(new_n322_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n342_), .B1(new_n292_), .B2(new_n343_), .ZN(new_n344_));
  AND3_X1   g143(.A1(new_n323_), .A2(new_n341_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n221_), .A2(new_n211_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT65), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n221_), .A2(new_n210_), .A3(new_n211_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n208_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n298_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G232gat), .A2(G233gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n353_), .B(KEYINPUT34), .Z(new_n354_));
  XOR2_X1   g153(.A(KEYINPUT73), .B(KEYINPUT35), .Z(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  OAI211_X1 g155(.A(KEYINPUT76), .B(new_n356_), .C1(new_n241_), .C2(new_n312_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n352_), .A2(new_n357_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n354_), .A2(new_n355_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(new_n358_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G190gat), .B(G218gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT75), .ZN(new_n363_));
  XOR2_X1   g162(.A(G134gat), .B(G162gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT36), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n361_), .A2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n358_), .B(new_n359_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT36), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n371_), .A3(new_n365_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n361_), .A2(KEYINPUT77), .A3(new_n366_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n369_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(G169gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT83), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT83), .B1(G183gat), .B2(G190gat), .ZN(new_n381_));
  OAI21_X1  g180(.A(KEYINPUT23), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT23), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n378_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n377_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NOR3_X1   g186(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n383_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n378_), .A2(KEYINPUT23), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n388_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  AND2_X1   g190(.A1(new_n391_), .A2(KEYINPUT84), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT25), .B(G183gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT26), .B(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(G169gat), .ZN(new_n398_));
  INV_X1    g197(.A(G176gat), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n397_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  AND2_X1   g199(.A1(new_n395_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n401_), .B1(new_n391_), .B2(KEYINPUT84), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n387_), .B1(new_n392_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT87), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n387_), .B(new_n404_), .C1(new_n392_), .C2(new_n402_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G227gat), .A2(G233gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(G15gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(KEYINPUT86), .B(G43gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  XOR2_X1   g212(.A(G71gat), .B(G99gat), .Z(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n409_), .A2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(G127gat), .B(G134gat), .ZN(new_n417_));
  AND2_X1   g216(.A1(new_n417_), .A2(KEYINPUT88), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n417_), .A2(KEYINPUT88), .ZN(new_n419_));
  XOR2_X1   g218(.A(G113gat), .B(G120gat), .Z(new_n420_));
  OR3_X1    g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n420_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT31), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n409_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n407_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n416_), .B(new_n425_), .C1(new_n428_), .C2(new_n415_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n406_), .A2(new_n408_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT87), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n415_), .B1(new_n431_), .B2(new_n409_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n416_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n424_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n429_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G228gat), .ZN(new_n436_));
  INV_X1    g235(.A(G233gat), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT93), .ZN(new_n439_));
  INV_X1    g238(.A(G204gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n439_), .B1(new_n440_), .B2(G197gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(G197gat), .ZN(new_n442_));
  INV_X1    g241(.A(G197gat), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n443_), .A2(KEYINPUT93), .A3(G204gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n442_), .A3(new_n444_), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n445_), .A2(KEYINPUT96), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(KEYINPUT96), .ZN(new_n447_));
  XOR2_X1   g246(.A(G211gat), .B(G218gat), .Z(new_n448_));
  NAND4_X1  g247(.A1(new_n446_), .A2(new_n447_), .A3(KEYINPUT21), .A4(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT21), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n441_), .A2(new_n444_), .A3(new_n451_), .A4(new_n442_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT94), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n443_), .A2(G204gat), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n451_), .B1(new_n455_), .B2(new_n442_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n456_), .A2(new_n448_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(KEYINPUT95), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT95), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n454_), .A2(new_n460_), .A3(new_n457_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n450_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT92), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(G141gat), .A2(G148gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT3), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G141gat), .A2(G148gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT89), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n465_), .B(new_n467_), .C1(KEYINPUT2), .C2(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G155gat), .B(G162gat), .Z(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G155gat), .A2(G162gat), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT1), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n474_), .B1(G155gat), .B2(G162gat), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(G155gat), .A3(G162gat), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT91), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n473_), .A2(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n477_), .B2(new_n476_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n469_), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n466_), .B(KEYINPUT90), .Z(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n472_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT29), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n438_), .B1(new_n462_), .B2(new_n485_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n454_), .A2(new_n460_), .A3(new_n457_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n460_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n449_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n489_), .B(new_n484_), .C1(new_n436_), .C2(new_n437_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G78gat), .B(G106gat), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n486_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT97), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n483_), .A2(KEYINPUT29), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G22gat), .B(G50gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT28), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n496_), .B(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n486_), .A2(new_n490_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n491_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n493_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n500_), .A2(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n502_), .A2(KEYINPUT97), .A3(new_n493_), .A4(new_n499_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT100), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G226gat), .A2(G233gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(KEYINPUT19), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT98), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT20), .B1(new_n489_), .B2(new_n403_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n389_), .A2(new_n390_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(G183gat), .B2(G190gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n377_), .B(KEYINPUT99), .Z(new_n514_));
  INV_X1    g313(.A(new_n388_), .ZN(new_n515_));
  AND2_X1   g314(.A1(new_n401_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n385_), .ZN(new_n517_));
  AOI22_X1  g316(.A1(new_n513_), .A2(new_n514_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n462_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n510_), .B1(new_n511_), .B2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G8gat), .B(G36gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT18), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G64gat), .B(G92gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  OAI211_X1 g323(.A(new_n518_), .B(new_n449_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n489_), .A2(new_n403_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n509_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(KEYINPUT20), .A4(new_n527_), .ZN(new_n528_));
  AND3_X1   g327(.A1(new_n520_), .A2(new_n524_), .A3(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n524_), .B1(new_n520_), .B2(new_n528_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n507_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n520_), .A2(new_n528_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n524_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n520_), .A2(new_n524_), .A3(new_n528_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(KEYINPUT100), .A3(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G1gat), .B(G29gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(KEYINPUT102), .ZN(new_n538_));
  XOR2_X1   g337(.A(G57gat), .B(G85gat), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n483_), .A2(new_n423_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(G225gat), .A2(G233gat), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n472_), .A2(new_n482_), .A3(new_n421_), .A4(new_n422_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n544_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n543_), .A2(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n544_), .A2(KEYINPUT4), .A3(new_n547_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT4), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n483_), .A2(new_n423_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(new_n546_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n546_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n546_), .B1(new_n544_), .B2(new_n547_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n543_), .B1(new_n556_), .B2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT33), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n545_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n542_), .B1(new_n562_), .B2(new_n557_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(KEYINPUT33), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n555_), .B1(new_n561_), .B2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n531_), .A2(new_n536_), .A3(new_n565_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n562_), .A2(new_n542_), .A3(new_n557_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n559_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n524_), .A2(KEYINPUT32), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n520_), .A2(new_n570_), .A3(new_n528_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n511_), .A2(new_n519_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n510_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n525_), .A2(new_n526_), .A3(KEYINPUT20), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n572_), .A2(new_n573_), .B1(new_n574_), .B2(new_n509_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n569_), .B(new_n571_), .C1(new_n570_), .C2(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n506_), .B1(new_n566_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT27), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n578_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n579_));
  OAI211_X1 g378(.A(KEYINPUT27), .B(new_n535_), .C1(new_n575_), .C2(new_n524_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n504_), .A2(new_n505_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n581_), .A2(new_n582_), .A3(new_n569_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n435_), .B1(new_n577_), .B2(new_n583_), .ZN(new_n584_));
  AND3_X1   g383(.A1(new_n568_), .A2(new_n429_), .A3(new_n434_), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n582_), .A2(new_n585_), .A3(new_n579_), .A4(new_n580_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT103), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n579_), .A2(new_n580_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT103), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(new_n582_), .A4(new_n585_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n375_), .B1(new_n584_), .B2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n345_), .A2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(G1gat), .B1(new_n593_), .B2(new_n568_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n292_), .B(KEYINPUT72), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n343_), .B1(new_n584_), .B2(new_n591_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT78), .B(KEYINPUT37), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n369_), .A2(new_n372_), .A3(new_n373_), .A4(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n372_), .A2(new_n367_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(KEYINPUT37), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  NAND4_X1  g401(.A1(new_n596_), .A2(new_n597_), .A3(new_n602_), .A4(new_n341_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT104), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n604_), .A2(new_n300_), .A3(new_n569_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n604_), .A2(KEYINPUT38), .A3(new_n300_), .A4(new_n569_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT105), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n606_), .A2(new_n607_), .ZN(new_n609_));
  OAI221_X1 g408(.A(new_n594_), .B1(KEYINPUT38), .B2(new_n605_), .C1(new_n608_), .C2(new_n609_), .ZN(G1324gat));
  NAND3_X1  g409(.A1(new_n604_), .A2(new_n301_), .A3(new_n581_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n345_), .A2(new_n581_), .A3(new_n592_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT107), .B(KEYINPUT39), .ZN(new_n613_));
  AND3_X1   g412(.A1(new_n612_), .A2(G8gat), .A3(new_n613_), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n613_), .B1(new_n612_), .B2(G8gat), .ZN(new_n615_));
  OAI21_X1  g414(.A(new_n611_), .B1(new_n614_), .B2(new_n615_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g416(.A(G15gat), .B1(new_n593_), .B2(new_n435_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT41), .ZN(new_n619_));
  NOR3_X1   g418(.A1(new_n603_), .A2(G15gat), .A3(new_n435_), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1326gat));
  OAI21_X1  g420(.A(G22gat), .B1(new_n593_), .B2(new_n582_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  OR2_X1    g423(.A1(new_n582_), .A2(G22gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n624_), .B1(new_n603_), .B2(new_n625_), .ZN(G1327gat));
  NAND2_X1  g425(.A1(new_n375_), .A2(new_n340_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n292_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n597_), .A2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(G29gat), .B1(new_n629_), .B2(new_n569_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n584_), .A2(new_n591_), .ZN(new_n631_));
  AND2_X1   g430(.A1(new_n599_), .A2(new_n601_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT110), .ZN(new_n634_));
  XOR2_X1   g433(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n635_));
  NAND3_X1  g434(.A1(new_n633_), .A2(new_n634_), .A3(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n602_), .B1(new_n584_), .B2(new_n591_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT43), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n635_), .ZN(new_n640_));
  OAI21_X1  g439(.A(KEYINPUT110), .B1(new_n637_), .B2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n636_), .A2(new_n639_), .A3(new_n641_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n323_), .A2(new_n340_), .A3(new_n344_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(KEYINPUT44), .A3(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n642_), .A2(new_n643_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(KEYINPUT111), .B(KEYINPUT44), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n644_), .B1(new_n645_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n569_), .A2(G29gat), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n630_), .B1(new_n648_), .B2(new_n649_), .ZN(G1328gat));
  INV_X1    g449(.A(G36gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n629_), .A2(new_n651_), .A3(new_n581_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT45), .Z(new_n653_));
  OAI211_X1 g452(.A(new_n581_), .B(new_n644_), .C1(new_n645_), .C2(new_n646_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n653_), .B1(new_n654_), .B2(G36gat), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT112), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT46), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n656_), .A2(new_n657_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n655_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n658_), .A2(new_n661_), .ZN(G1329gat));
  INV_X1    g461(.A(new_n435_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G43gat), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n629_), .A2(new_n663_), .ZN(new_n665_));
  OAI22_X1  g464(.A1(new_n647_), .A2(new_n664_), .B1(G43gat), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g466(.A(G50gat), .B1(new_n629_), .B2(new_n506_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n506_), .A2(G50gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n648_), .B2(new_n669_), .ZN(G1331gat));
  NOR2_X1   g469(.A1(new_n322_), .A2(new_n340_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n595_), .A2(new_n592_), .A3(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G57gat), .B1(new_n672_), .B2(new_n568_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n631_), .A2(new_n343_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT113), .Z(new_n675_));
  NAND4_X1  g474(.A1(new_n675_), .A2(new_n292_), .A3(new_n602_), .A4(new_n341_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n568_), .A2(G57gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(G1332gat));
  OAI21_X1  g477(.A(G64gat), .B1(new_n672_), .B2(new_n588_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT48), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n588_), .A2(G64gat), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n676_), .B2(new_n681_), .ZN(G1333gat));
  OAI21_X1  g481(.A(G71gat), .B1(new_n672_), .B2(new_n435_), .ZN(new_n683_));
  XOR2_X1   g482(.A(KEYINPUT114), .B(KEYINPUT49), .Z(new_n684_));
  XNOR2_X1  g483(.A(new_n683_), .B(new_n684_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n435_), .A2(G71gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n676_), .B2(new_n686_), .ZN(G1334gat));
  OAI21_X1  g486(.A(G78gat), .B1(new_n672_), .B2(new_n582_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT50), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n506_), .A2(new_n249_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n676_), .B2(new_n690_), .ZN(G1335gat));
  NOR3_X1   g490(.A1(new_n293_), .A2(new_n322_), .A3(new_n341_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n642_), .A2(new_n692_), .ZN(new_n693_));
  OAI21_X1  g492(.A(G85gat), .B1(new_n693_), .B2(new_n568_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n596_), .A2(new_n627_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n675_), .A2(new_n695_), .ZN(new_n696_));
  OR2_X1    g495(.A1(new_n568_), .A2(G85gat), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n694_), .B1(new_n696_), .B2(new_n697_), .ZN(G1336gat));
  INV_X1    g497(.A(new_n696_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G92gat), .B1(new_n699_), .B2(new_n581_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n693_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n581_), .A2(G92gat), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT115), .Z(new_n703_));
  AOI21_X1  g502(.A(new_n700_), .B1(new_n701_), .B2(new_n703_), .ZN(G1337gat));
  OAI21_X1  g503(.A(G99gat), .B1(new_n693_), .B2(new_n435_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n435_), .A2(new_n207_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n696_), .B2(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g507(.A1(new_n696_), .A2(G106gat), .A3(new_n582_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n642_), .A2(new_n506_), .A3(new_n692_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(G106gat), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n711_), .A2(KEYINPUT52), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n711_), .A2(KEYINPUT52), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n709_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n714_), .B(new_n716_), .ZN(G1339gat));
  AND3_X1   g516(.A1(new_n290_), .A2(new_n291_), .A3(new_n671_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT54), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n718_), .A2(KEYINPUT117), .A3(new_n719_), .A4(new_n602_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n290_), .A2(new_n291_), .A3(new_n671_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n632_), .A2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n722_), .B2(new_n719_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT117), .B1(new_n722_), .B2(new_n719_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT118), .ZN(new_n726_));
  INV_X1    g525(.A(new_n275_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n261_), .B1(new_n350_), .B2(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n259_), .B2(new_n256_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n726_), .B1(new_n729_), .B2(new_n277_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT55), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n278_), .A2(new_n731_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n260_), .A2(new_n276_), .A3(KEYINPUT55), .A4(new_n277_), .ZN(new_n733_));
  AOI21_X1  g532(.A(KEYINPUT71), .B1(new_n254_), .B2(new_n255_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n258_), .A2(new_n257_), .A3(KEYINPUT12), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n734_), .A2(new_n735_), .ZN(new_n736_));
  OAI211_X1 g535(.A(KEYINPUT118), .B(new_n279_), .C1(new_n736_), .C2(new_n728_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n730_), .A2(new_n732_), .A3(new_n733_), .A4(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n285_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT56), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n739_), .A2(KEYINPUT121), .A3(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n319_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n316_), .A2(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n319_), .B1(new_n314_), .B2(new_n310_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n744_), .A2(KEYINPUT120), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n310_), .B1(new_n307_), .B2(new_n296_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n306_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n744_), .A2(KEYINPUT120), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n743_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n286_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n738_), .A2(KEYINPUT56), .A3(new_n285_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT121), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  AOI21_X1  g552(.A(KEYINPUT56), .B1(new_n738_), .B2(new_n285_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n741_), .B(new_n750_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT58), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n739_), .A2(new_n740_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n758_), .A2(new_n752_), .A3(new_n751_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n759_), .A2(KEYINPUT58), .A3(new_n741_), .A4(new_n750_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n757_), .A2(new_n632_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n288_), .A2(new_n749_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT119), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n751_), .A2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n764_), .A2(new_n754_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n739_), .A2(KEYINPUT119), .A3(new_n740_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n322_), .A2(new_n286_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n762_), .B1(new_n765_), .B2(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(KEYINPUT57), .A3(new_n374_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT57), .ZN(new_n772_));
  INV_X1    g571(.A(new_n762_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n758_), .A2(new_n763_), .A3(new_n751_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n767_), .B1(new_n754_), .B2(KEYINPUT119), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n773_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n776_), .B2(new_n375_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n761_), .A2(new_n771_), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n725_), .B1(new_n778_), .B2(new_n340_), .ZN(new_n779_));
  NOR4_X1   g578(.A1(new_n506_), .A2(new_n581_), .A3(new_n435_), .A4(new_n568_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT59), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n779_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT123), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n771_), .A2(new_n777_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n602_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT122), .B1(new_n786_), .B2(new_n760_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n786_), .A2(KEYINPUT122), .A3(new_n760_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n341_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n784_), .B1(new_n790_), .B2(new_n725_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT122), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n761_), .A2(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n793_), .A2(new_n789_), .A3(new_n777_), .A4(new_n771_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n340_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n725_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n795_), .A2(KEYINPUT123), .A3(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n791_), .A2(new_n797_), .A3(new_n780_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n783_), .B1(new_n798_), .B2(KEYINPUT59), .ZN(new_n799_));
  INV_X1    g598(.A(G113gat), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n343_), .A2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT123), .B1(new_n795_), .B2(new_n796_), .ZN(new_n802_));
  AOI211_X1 g601(.A(new_n784_), .B(new_n725_), .C1(new_n794_), .C2(new_n340_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n804_), .A2(new_n322_), .A3(new_n780_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n799_), .A2(new_n801_), .B1(new_n805_), .B2(new_n800_), .ZN(G1340gat));
  OAI21_X1  g605(.A(new_n595_), .B1(new_n779_), .B2(new_n782_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n798_), .B2(KEYINPUT59), .ZN(new_n808_));
  INV_X1    g607(.A(G120gat), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n809_), .B1(new_n293_), .B2(KEYINPUT60), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(KEYINPUT60), .B2(new_n809_), .ZN(new_n811_));
  OAI22_X1  g610(.A1(new_n808_), .A2(new_n809_), .B1(new_n798_), .B2(new_n811_), .ZN(G1341gat));
  INV_X1    g611(.A(KEYINPUT124), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n341_), .A2(new_n813_), .A3(G127gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n813_), .B2(G127gat), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n804_), .A2(new_n341_), .A3(new_n780_), .ZN(new_n816_));
  INV_X1    g615(.A(G127gat), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n799_), .A2(new_n815_), .B1(new_n816_), .B2(new_n817_), .ZN(G1342gat));
  INV_X1    g617(.A(G134gat), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n602_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n804_), .A2(new_n375_), .A3(new_n780_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n799_), .A2(new_n820_), .B1(new_n821_), .B2(new_n819_), .ZN(G1343gat));
  NOR3_X1   g621(.A1(new_n802_), .A2(new_n803_), .A3(new_n663_), .ZN(new_n823_));
  INV_X1    g622(.A(G141gat), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n581_), .A2(new_n582_), .A3(new_n568_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n823_), .A2(new_n824_), .A3(new_n322_), .A4(new_n825_), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n791_), .A2(new_n435_), .A3(new_n797_), .A4(new_n825_), .ZN(new_n827_));
  OAI21_X1  g626(.A(G141gat), .B1(new_n827_), .B2(new_n343_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1344gat));
  INV_X1    g628(.A(G148gat), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n823_), .A2(new_n830_), .A3(new_n595_), .A4(new_n825_), .ZN(new_n831_));
  OAI21_X1  g630(.A(G148gat), .B1(new_n827_), .B2(new_n596_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(G1345gat));
  XNOR2_X1  g632(.A(KEYINPUT61), .B(G155gat), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n823_), .A2(new_n341_), .A3(new_n825_), .A4(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n827_), .B2(new_n340_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1346gat));
  OAI21_X1  g637(.A(G162gat), .B1(new_n827_), .B2(new_n602_), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n374_), .A2(G162gat), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n839_), .B1(new_n827_), .B2(new_n840_), .ZN(G1347gat));
  INV_X1    g640(.A(KEYINPUT62), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n581_), .A2(new_n585_), .ZN(new_n843_));
  NOR4_X1   g642(.A1(new_n779_), .A2(new_n343_), .A3(new_n506_), .A4(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT22), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n842_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(G169gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n398_), .B1(new_n844_), .B2(new_n842_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n847_), .B1(new_n846_), .B2(new_n848_), .ZN(G1348gat));
  NOR3_X1   g648(.A1(new_n596_), .A2(new_n399_), .A3(new_n843_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n791_), .A2(new_n582_), .A3(new_n797_), .A4(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n804_), .A2(KEYINPUT125), .A3(new_n582_), .A4(new_n850_), .ZN(new_n854_));
  OR3_X1    g653(.A1(new_n779_), .A2(new_n506_), .A3(new_n843_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n855_), .A2(new_n293_), .ZN(new_n856_));
  AOI22_X1  g655(.A1(new_n853_), .A2(new_n854_), .B1(new_n856_), .B2(new_n399_), .ZN(G1349gat));
  NOR2_X1   g656(.A1(new_n843_), .A2(new_n340_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n804_), .A2(new_n582_), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(G183gat), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n779_), .A2(new_n506_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n843_), .A2(new_n393_), .A3(new_n340_), .ZN(new_n862_));
  AOI22_X1  g661(.A1(new_n859_), .A2(new_n860_), .B1(new_n861_), .B2(new_n862_), .ZN(G1350gat));
  OAI21_X1  g662(.A(G190gat), .B1(new_n855_), .B2(new_n602_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n375_), .A2(new_n394_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n855_), .B2(new_n865_), .ZN(G1351gat));
  NOR3_X1   g665(.A1(new_n588_), .A2(new_n582_), .A3(new_n569_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n791_), .A2(new_n435_), .A3(new_n797_), .A4(new_n867_), .ZN(new_n868_));
  OAI211_X1 g667(.A(KEYINPUT126), .B(G197gat), .C1(new_n868_), .C2(new_n343_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT126), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n343_), .B1(new_n870_), .B2(new_n443_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n823_), .A2(new_n867_), .A3(new_n871_), .A4(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n869_), .A2(new_n873_), .ZN(G1352gat));
  NAND4_X1  g673(.A1(new_n823_), .A2(new_n440_), .A3(new_n595_), .A4(new_n867_), .ZN(new_n875_));
  OAI21_X1  g674(.A(G204gat), .B1(new_n868_), .B2(new_n596_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n875_), .A2(new_n876_), .ZN(G1353gat));
  NOR2_X1   g676(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n341_), .A2(new_n880_), .ZN(new_n881_));
  XOR2_X1   g680(.A(new_n881_), .B(KEYINPUT127), .Z(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n823_), .A2(new_n867_), .A3(new_n879_), .A4(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n878_), .B1(new_n868_), .B2(new_n882_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1354gat));
  OAI21_X1  g685(.A(G218gat), .B1(new_n868_), .B2(new_n602_), .ZN(new_n887_));
  OR2_X1    g686(.A1(new_n374_), .A2(G218gat), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n868_), .B2(new_n888_), .ZN(G1355gat));
endmodule


