//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n734_, new_n735_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n857_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n879_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n886_, new_n887_, new_n889_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G211gat), .B(G218gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT96), .ZN(new_n204_));
  XOR2_X1   g003(.A(G197gat), .B(G204gat), .Z(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT21), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT95), .ZN(new_n208_));
  OR3_X1    g007(.A1(new_n205_), .A2(new_n208_), .A3(KEYINPUT21), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n208_), .B1(new_n205_), .B2(KEYINPUT21), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n209_), .A2(new_n204_), .A3(new_n206_), .A4(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n207_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n215_), .B(new_n216_), .C1(G183gat), .C2(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  XOR2_X1   g017(.A(KEYINPUT22), .B(G169gat), .Z(new_n219_));
  OAI211_X1 g018(.A(new_n217_), .B(new_n218_), .C1(G176gat), .C2(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n221_), .B(KEYINPUT100), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT25), .B(G183gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n222_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n213_), .B(KEYINPUT23), .ZN(new_n226_));
  OR3_X1    g025(.A1(KEYINPUT90), .A2(G169gat), .A3(G176gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT90), .B1(G169gat), .B2(G176gat), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n227_), .A2(KEYINPUT24), .A3(new_n228_), .ZN(new_n229_));
  AOI22_X1  g028(.A1(new_n227_), .A2(new_n228_), .B1(KEYINPUT24), .B2(new_n218_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n226_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n220_), .B1(new_n225_), .B2(new_n231_), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n212_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G226gat), .A2(G233gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(KEYINPUT19), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT20), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT91), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n219_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G176gat), .ZN(new_n240_));
  INV_X1    g039(.A(G169gat), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n241_), .A2(KEYINPUT22), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n240_), .B1(new_n242_), .B2(new_n238_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n217_), .B(new_n218_), .C1(new_n239_), .C2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT89), .B1(new_n245_), .B2(G183gat), .ZN(new_n246_));
  OAI211_X1 g045(.A(new_n221_), .B(new_n246_), .C1(new_n223_), .C2(KEYINPUT89), .ZN(new_n247_));
  OAI211_X1 g046(.A(new_n247_), .B(new_n226_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n244_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n237_), .B1(new_n212_), .B2(new_n249_), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n233_), .A2(new_n236_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n212_), .A2(new_n232_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT20), .B1(new_n212_), .B2(new_n249_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n235_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT101), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(KEYINPUT101), .B(new_n235_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n251_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G8gat), .B(G36gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(G64gat), .B(G92gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT102), .B(KEYINPUT18), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n259_), .A2(new_n265_), .ZN(new_n266_));
  AOI211_X1 g065(.A(new_n264_), .B(new_n251_), .C1(new_n257_), .C2(new_n258_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n202_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n202_), .B1(new_n259_), .B2(new_n265_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n264_), .B(KEYINPUT107), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT105), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n232_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT97), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n207_), .A2(new_n211_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n212_), .A2(KEYINPUT97), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n232_), .A2(new_n271_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n272_), .A2(new_n274_), .A3(new_n275_), .A4(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n236_), .B1(new_n277_), .B2(new_n250_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n252_), .B(KEYINPUT20), .C1(new_n212_), .C2(new_n249_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n279_), .A2(new_n235_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n270_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n269_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n268_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n274_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n273_), .B1(new_n207_), .B2(new_n211_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT29), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G155gat), .B(G162gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n287_), .A2(KEYINPUT1), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n288_), .A2(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n289_), .B(KEYINPUT3), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT92), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT2), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT2), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n292_), .A2(new_n296_), .A3(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n295_), .A2(new_n298_), .A3(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT93), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n287_), .B1(new_n301_), .B2(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n295_), .A2(KEYINPUT93), .A3(new_n298_), .A4(new_n300_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n294_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  OAI22_X1  g104(.A1(new_n284_), .A2(new_n285_), .B1(new_n286_), .B2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(G228gat), .ZN(new_n307_));
  INV_X1    g106(.A(G233gat), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(KEYINPUT98), .A3(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n310_), .ZN(new_n311_));
  AOI21_X1  g110(.A(KEYINPUT98), .B1(new_n306_), .B2(new_n309_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n305_), .A2(new_n286_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n309_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n212_), .A2(new_n314_), .ZN(new_n315_));
  OAI22_X1  g114(.A1(new_n311_), .A2(new_n312_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G78gat), .B(G106gat), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n319_));
  XOR2_X1   g118(.A(G22gat), .B(G50gat), .Z(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n305_), .A2(new_n286_), .A3(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n321_), .B1(new_n305_), .B2(new_n286_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n319_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n324_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n319_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n322_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n318_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n317_), .A2(KEYINPUT99), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n325_), .A2(new_n328_), .A3(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n316_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n313_), .A2(new_n315_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT98), .ZN(new_n335_));
  INV_X1    g134(.A(new_n305_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n274_), .A2(new_n275_), .B1(new_n336_), .B2(KEYINPUT29), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n335_), .B1(new_n337_), .B2(new_n314_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n334_), .B1(new_n338_), .B2(new_n310_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n332_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(new_n329_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n333_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n283_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G71gat), .B(G99gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(G43gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n249_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G127gat), .B(G134gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(G113gat), .B(G120gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n347_), .B(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G227gat), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(G15gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n352_), .B(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT30), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT31), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n351_), .B(new_n356_), .Z(new_n357_));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n305_), .A2(new_n350_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n305_), .A2(new_n350_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363_));
  NOR3_X1   g162(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n363_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n359_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  XNOR2_X1  g166(.A(G1gat), .B(G29gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(G85gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT0), .B(G57gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n369_), .B(new_n370_), .Z(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n358_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n367_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n305_), .A2(new_n350_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(KEYINPUT4), .A3(new_n360_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n358_), .B1(new_n376_), .B2(new_n365_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n373_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n371_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n357_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n344_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n251_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n258_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT101), .B1(new_n279_), .B2(new_n235_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n384_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n264_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n259_), .A2(new_n265_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n390_), .A2(new_n202_), .B1(new_n281_), .B2(new_n269_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n380_), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n391_), .A2(KEYINPUT108), .A3(new_n343_), .A4(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT108), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n341_), .A3(new_n333_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n394_), .B1(new_n283_), .B2(new_n395_), .ZN(new_n396_));
  OAI211_X1 g195(.A(KEYINPUT33), .B(new_n371_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT104), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n375_), .A2(KEYINPUT104), .A3(new_n360_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n359_), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n376_), .A2(new_n358_), .A3(new_n365_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n401_), .A2(new_n372_), .A3(new_n402_), .ZN(new_n403_));
  AND4_X1   g202(.A1(new_n389_), .A2(new_n388_), .A3(new_n397_), .A4(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT33), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n379_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT103), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n379_), .A2(KEYINPUT103), .A3(new_n405_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n265_), .A2(KEYINPUT32), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT106), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n413_), .B(new_n414_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n374_), .A2(new_n379_), .B1(new_n259_), .B2(new_n411_), .ZN(new_n416_));
  AOI22_X1  g215(.A1(new_n404_), .A2(new_n410_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n393_), .B(new_n396_), .C1(new_n417_), .C2(new_n343_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n383_), .B1(new_n418_), .B2(new_n357_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G15gat), .B(G22gat), .ZN(new_n420_));
  INV_X1    g219(.A(G1gat), .ZN(new_n421_));
  INV_X1    g220(.A(G8gat), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT14), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n420_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G1gat), .B(G8gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G29gat), .B(G36gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G43gat), .B(G50gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  XOR2_X1   g228(.A(new_n426_), .B(new_n429_), .Z(new_n430_));
  NAND2_X1  g229(.A1(G229gat), .A2(G233gat), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n429_), .B(KEYINPUT15), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(new_n426_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n426_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n432_), .B1(new_n435_), .B2(new_n429_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n430_), .A2(new_n432_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G113gat), .B(G141gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G169gat), .B(G197gat), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n438_), .B(new_n439_), .Z(new_n440_));
  XOR2_X1   g239(.A(new_n440_), .B(KEYINPUT86), .Z(new_n441_));
  OR2_X1    g240(.A1(new_n437_), .A2(new_n441_), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n437_), .A2(KEYINPUT87), .A3(new_n440_), .ZN(new_n443_));
  AOI21_X1  g242(.A(KEYINPUT87), .B1(new_n437_), .B2(new_n440_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n442_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  OAI211_X1 g246(.A(KEYINPUT88), .B(new_n442_), .C1(new_n443_), .C2(new_n444_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n419_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT13), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G57gat), .B(G64gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT11), .ZN(new_n454_));
  XNOR2_X1  g253(.A(KEYINPUT69), .B(G71gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(G78gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(G78gat), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n455_), .B(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n453_), .A2(KEYINPUT11), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n457_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT66), .ZN(new_n463_));
  INV_X1    g262(.A(G99gat), .ZN(new_n464_));
  INV_X1    g263(.A(G106gat), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .A4(KEYINPUT7), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT7), .ZN(new_n467_));
  OAI22_X1  g266(.A1(new_n467_), .A2(KEYINPUT66), .B1(G99gat), .B2(G106gat), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n463_), .A2(KEYINPUT7), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n466_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT6), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT64), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT64), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT6), .ZN(new_n474_));
  AND2_X1   g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n472_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n475_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n470_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  AND2_X1   g277(.A1(G85gat), .A2(G92gat), .ZN(new_n479_));
  NOR2_X1   g278(.A1(G85gat), .A2(G92gat), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(KEYINPUT67), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT8), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT65), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n476_), .A2(new_n477_), .ZN(new_n486_));
  OR2_X1    g285(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n487_), .A2(new_n465_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(G85gat), .ZN(new_n490_));
  INV_X1    g289(.A(G92gat), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G85gat), .A2(G92gat), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n492_), .A2(KEYINPUT9), .A3(new_n493_), .ZN(new_n494_));
  NOR2_X1   g293(.A1(new_n493_), .A2(KEYINPUT9), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n489_), .A2(new_n494_), .A3(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n485_), .B1(new_n486_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n475_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n473_), .A2(KEYINPUT6), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n471_), .A2(KEYINPUT64), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n499_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n472_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n495_), .B1(new_n481_), .B2(KEYINPUT9), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n504_), .A2(KEYINPUT65), .A3(new_n489_), .A4(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n498_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n484_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n481_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n509_), .B1(new_n504_), .B2(new_n470_), .ZN(new_n510_));
  AND2_X1   g309(.A1(KEYINPUT68), .A2(KEYINPUT8), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI22_X1  g311(.A1(new_n482_), .A2(KEYINPUT68), .B1(new_n510_), .B2(new_n512_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n462_), .B1(new_n508_), .B2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT71), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n482_), .A2(KEYINPUT68), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n510_), .A2(new_n512_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  AOI22_X1  g318(.A1(new_n483_), .A2(new_n482_), .B1(new_n498_), .B2(new_n506_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n462_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT70), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n519_), .A2(new_n520_), .A3(KEYINPUT70), .A4(new_n521_), .ZN(new_n525_));
  OAI211_X1 g324(.A(KEYINPUT71), .B(new_n462_), .C1(new_n508_), .C2(new_n513_), .ZN(new_n526_));
  NAND4_X1  g325(.A1(new_n516_), .A2(new_n524_), .A3(new_n525_), .A4(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(G230gat), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n528_), .A2(new_n308_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n508_), .A2(new_n513_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n529_), .B1(new_n531_), .B2(new_n521_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(KEYINPUT72), .B(KEYINPUT12), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n514_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n519_), .A2(new_n520_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT72), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n537_), .A2(KEYINPUT12), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n536_), .A2(new_n462_), .A3(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n532_), .A2(new_n535_), .A3(new_n540_), .ZN(new_n541_));
  XOR2_X1   g340(.A(G120gat), .B(G148gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT74), .B(KEYINPUT5), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G176gat), .B(G204gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n530_), .A2(new_n541_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT75), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n530_), .A2(KEYINPUT75), .A3(new_n541_), .A4(new_n547_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n530_), .A2(new_n541_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT73), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT73), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n530_), .A2(new_n555_), .A3(new_n541_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(new_n546_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT76), .ZN(new_n558_));
  AND3_X1   g357(.A1(new_n552_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n558_), .B1(new_n552_), .B2(new_n557_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n452_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n514_), .A2(new_n538_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n533_), .B1(new_n536_), .B2(new_n462_), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n529_), .A2(new_n527_), .B1(new_n564_), .B2(new_n532_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT75), .B1(new_n565_), .B2(new_n547_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n551_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n530_), .A2(new_n555_), .A3(new_n541_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n555_), .B1(new_n530_), .B2(new_n541_), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n569_), .A2(new_n570_), .A3(new_n547_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT76), .B1(new_n568_), .B2(new_n571_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n552_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(KEYINPUT13), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n561_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n426_), .B(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(new_n521_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(G127gat), .B(G155gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G183gat), .B(G211gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT17), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n584_), .A2(KEYINPUT17), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n579_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT85), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n579_), .A2(new_n585_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT84), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(KEYINPUT81), .A2(KEYINPUT37), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT35), .ZN(new_n593_));
  XNOR2_X1  g392(.A(KEYINPUT77), .B(KEYINPUT34), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G232gat), .A2(G233gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n594_), .B(new_n595_), .ZN(new_n596_));
  AOI22_X1  g395(.A1(new_n531_), .A2(new_n429_), .B1(new_n593_), .B2(new_n596_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n536_), .A2(KEYINPUT78), .A3(new_n433_), .ZN(new_n598_));
  AOI21_X1  g397(.A(KEYINPUT78), .B1(new_n536_), .B2(new_n433_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n597_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n596_), .A2(new_n593_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  OAI221_X1 g401(.A(new_n597_), .B1(new_n593_), .B2(new_n596_), .C1(new_n598_), .C2(new_n599_), .ZN(new_n603_));
  XOR2_X1   g402(.A(G190gat), .B(G218gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT79), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(KEYINPUT80), .B(KEYINPUT36), .Z(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  AND3_X1   g408(.A1(new_n602_), .A2(new_n603_), .A3(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n607_), .B(KEYINPUT36), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n611_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n592_), .B1(new_n610_), .B2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(KEYINPUT81), .A2(KEYINPUT37), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT82), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n592_), .B(new_n615_), .C1(new_n610_), .C2(new_n612_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n591_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  AND3_X1   g418(.A1(new_n451_), .A2(new_n576_), .A3(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(new_n421_), .A3(new_n380_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT38), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n610_), .A2(new_n612_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n419_), .A2(new_n591_), .A3(new_n624_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n575_), .A2(new_n450_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n421_), .B1(new_n627_), .B2(new_n380_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n623_), .A2(new_n628_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n629_), .B1(new_n622_), .B2(new_n621_), .ZN(G1324gat));
  NAND3_X1  g429(.A1(new_n620_), .A2(new_n422_), .A3(new_n283_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT39), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n627_), .A2(new_n283_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n633_), .B2(G8gat), .ZN(new_n634_));
  AOI211_X1 g433(.A(KEYINPUT39), .B(new_n422_), .C1(new_n627_), .C2(new_n283_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n631_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT40), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(G1325gat));
  INV_X1    g437(.A(new_n357_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n353_), .B1(new_n627_), .B2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT41), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n620_), .A2(new_n353_), .A3(new_n639_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1326gat));
  INV_X1    g442(.A(G22gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n620_), .A2(new_n644_), .A3(new_n343_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n627_), .A2(new_n343_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n646_), .B1(new_n647_), .B2(G22gat), .ZN(new_n648_));
  AOI211_X1 g447(.A(KEYINPUT42), .B(new_n644_), .C1(new_n627_), .C2(new_n343_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT109), .ZN(G1327gat));
  NAND2_X1  g450(.A1(new_n624_), .A2(new_n591_), .ZN(new_n652_));
  NOR4_X1   g451(.A1(new_n419_), .A2(new_n450_), .A3(new_n575_), .A4(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(G29gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n653_), .A2(new_n654_), .A3(new_n380_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT112), .B1(KEYINPUT111), .B2(KEYINPUT44), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n626_), .A2(new_n591_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT110), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n658_), .B(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n418_), .A2(new_n357_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(new_n382_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n617_), .A2(new_n618_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n661_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n419_), .A2(KEYINPUT43), .A3(new_n664_), .ZN(new_n667_));
  OAI22_X1  g466(.A1(new_n666_), .A2(new_n667_), .B1(KEYINPUT112), .B2(KEYINPUT44), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n657_), .B1(new_n660_), .B2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n658_), .B(KEYINPUT110), .ZN(new_n670_));
  NOR2_X1   g469(.A1(KEYINPUT112), .A2(KEYINPUT44), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n663_), .A2(new_n661_), .A3(new_n665_), .ZN(new_n672_));
  OAI21_X1  g471(.A(KEYINPUT43), .B1(new_n419_), .B2(new_n664_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n671_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n670_), .A2(new_n674_), .A3(new_n656_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n392_), .B1(new_n669_), .B2(new_n675_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n655_), .B1(new_n676_), .B2(new_n654_), .ZN(G1328gat));
  INV_X1    g476(.A(G36gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n653_), .A2(new_n678_), .A3(new_n283_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT45), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n391_), .B1(new_n669_), .B2(new_n675_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n680_), .B1(new_n681_), .B2(new_n678_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT46), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n680_), .B(KEYINPUT46), .C1(new_n681_), .C2(new_n678_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(G1329gat));
  INV_X1    g485(.A(G43gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n653_), .A2(new_n687_), .A3(new_n639_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n357_), .B1(new_n669_), .B2(new_n675_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(new_n687_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT47), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI211_X1 g491(.A(KEYINPUT47), .B(new_n688_), .C1(new_n689_), .C2(new_n687_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1330gat));
  AOI21_X1  g493(.A(G50gat), .B1(new_n653_), .B2(new_n343_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n669_), .A2(new_n675_), .ZN(new_n696_));
  AND2_X1   g495(.A1(new_n343_), .A2(G50gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n695_), .B1(new_n696_), .B2(new_n697_), .ZN(G1331gat));
  NOR2_X1   g497(.A1(new_n576_), .A2(new_n449_), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n625_), .A2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G57gat), .B1(new_n701_), .B2(new_n392_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n419_), .A2(new_n449_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n703_), .A2(new_n575_), .A3(new_n619_), .ZN(new_n704_));
  INV_X1    g503(.A(G57gat), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(new_n380_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n702_), .A2(new_n706_), .ZN(G1332gat));
  INV_X1    g506(.A(G64gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n708_), .B1(new_n700_), .B2(new_n283_), .ZN(new_n709_));
  XOR2_X1   g508(.A(new_n709_), .B(KEYINPUT48), .Z(new_n710_));
  NAND3_X1  g509(.A1(new_n704_), .A2(new_n708_), .A3(new_n283_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1333gat));
  INV_X1    g511(.A(G71gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n713_), .B1(new_n700_), .B2(new_n639_), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT113), .B(KEYINPUT49), .Z(new_n715_));
  XNOR2_X1  g514(.A(new_n714_), .B(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n704_), .A2(new_n713_), .A3(new_n639_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1334gat));
  AOI21_X1  g517(.A(new_n458_), .B1(new_n700_), .B2(new_n343_), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n704_), .A2(new_n458_), .A3(new_n343_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1335gat));
  INV_X1    g522(.A(new_n591_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n576_), .A2(new_n449_), .A3(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n725_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n726_), .A2(new_n490_), .A3(new_n392_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n703_), .A2(new_n575_), .A3(new_n591_), .A4(new_n624_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT115), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n490_), .B1(new_n729_), .B2(new_n392_), .ZN(new_n730_));
  OR2_X1    g529(.A1(new_n730_), .A2(KEYINPUT116), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(KEYINPUT116), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n727_), .B1(new_n731_), .B2(new_n732_), .ZN(G1336gat));
  OAI21_X1  g532(.A(G92gat), .B1(new_n726_), .B2(new_n391_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n283_), .A2(new_n491_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n729_), .B2(new_n735_), .ZN(G1337gat));
  XOR2_X1   g535(.A(new_n728_), .B(KEYINPUT115), .Z(new_n737_));
  NAND4_X1  g536(.A1(new_n737_), .A2(new_n639_), .A3(new_n487_), .A4(new_n488_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G99gat), .B1(new_n726_), .B2(new_n357_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT51), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n738_), .A2(new_n742_), .A3(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1338gat));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745_));
  OAI211_X1 g544(.A(new_n343_), .B(new_n725_), .C1(new_n666_), .C2(new_n667_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT117), .ZN(new_n747_));
  AND3_X1   g546(.A1(new_n746_), .A2(new_n747_), .A3(G106gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n746_), .B2(G106gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n746_), .A2(G106gat), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT117), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n746_), .A2(new_n747_), .A3(G106gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n752_), .A2(KEYINPUT52), .A3(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n342_), .A2(G106gat), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n737_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n750_), .A2(new_n754_), .A3(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n757_), .A2(new_n759_), .ZN(new_n760_));
  NAND4_X1  g559(.A1(new_n750_), .A2(new_n754_), .A3(new_n756_), .A4(new_n758_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1339gat));
  NOR2_X1   g561(.A1(new_n443_), .A2(new_n444_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n431_), .B1(new_n435_), .B2(new_n429_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n434_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n440_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n763_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n767_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT55), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n541_), .A2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n532_), .A2(new_n535_), .A3(KEYINPUT55), .A4(new_n540_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n564_), .A2(KEYINPUT119), .A3(new_n524_), .A4(new_n525_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n529_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n535_), .A2(new_n524_), .A3(new_n540_), .A4(new_n525_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT119), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n774_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n772_), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT56), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n778_), .A2(new_n779_), .A3(new_n547_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n773_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n781_), .A2(new_n770_), .A3(new_n771_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT56), .B1(new_n782_), .B2(new_n546_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n449_), .B(new_n552_), .C1(new_n780_), .C2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n624_), .B1(new_n768_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT57), .B1(new_n785_), .B2(KEYINPUT120), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT120), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT57), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n552_), .A2(new_n449_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n779_), .B1(new_n778_), .B2(new_n547_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n782_), .A2(KEYINPUT56), .A3(new_n546_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n789_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n572_), .A2(new_n573_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n792_), .B1(new_n793_), .B2(new_n767_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n787_), .B(new_n788_), .C1(new_n794_), .C2(new_n624_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n552_), .A2(new_n767_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n796_), .B1(new_n780_), .B2(new_n783_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT58), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n796_), .B(KEYINPUT58), .C1(new_n783_), .C2(new_n780_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n665_), .A3(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n786_), .A2(new_n795_), .A3(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n591_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n561_), .A2(new_n574_), .A3(new_n450_), .A4(new_n619_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT54), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n804_), .B(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n803_), .A2(new_n807_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n344_), .A2(new_n380_), .A3(new_n639_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT59), .B1(new_n808_), .B2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n806_), .B1(new_n802_), .B2(new_n591_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT59), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n812_), .A2(new_n813_), .A3(new_n809_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n811_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(G113gat), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n450_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n809_), .B1(new_n803_), .B2(new_n807_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n816_), .B1(new_n819_), .B2(new_n450_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n820_), .A2(new_n821_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n817_), .B1(new_n822_), .B2(new_n823_), .ZN(G1340gat));
  OAI21_X1  g623(.A(G120gat), .B1(new_n815_), .B2(new_n576_), .ZN(new_n825_));
  INV_X1    g624(.A(G120gat), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n826_), .B1(new_n576_), .B2(KEYINPUT60), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(KEYINPUT60), .B2(new_n826_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n825_), .B1(new_n819_), .B2(new_n828_), .ZN(G1341gat));
  INV_X1    g628(.A(G127gat), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n815_), .A2(new_n830_), .A3(new_n591_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n830_), .B1(new_n819_), .B2(new_n591_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT122), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  OR2_X1    g633(.A1(new_n832_), .A2(new_n833_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(G1342gat));
  INV_X1    g635(.A(G134gat), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n664_), .A2(new_n837_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n811_), .B2(new_n814_), .ZN(new_n839_));
  AOI211_X1 g638(.A(KEYINPUT123), .B(G134gat), .C1(new_n818_), .C2(new_n624_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT123), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n799_), .A2(new_n665_), .A3(new_n800_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n787_), .B1(new_n794_), .B2(new_n624_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(KEYINPUT57), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n724_), .B1(new_n844_), .B2(new_n795_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n624_), .B(new_n810_), .C1(new_n845_), .C2(new_n806_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n841_), .B1(new_n846_), .B2(new_n837_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n839_), .B1(new_n840_), .B2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(KEYINPUT124), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT124), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n839_), .B(new_n850_), .C1(new_n840_), .C2(new_n847_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n849_), .A2(new_n851_), .ZN(G1343gat));
  NOR3_X1   g651(.A1(new_n283_), .A2(new_n392_), .A3(new_n639_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n808_), .A2(new_n343_), .A3(new_n853_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n854_), .A2(new_n450_), .ZN(new_n855_));
  XOR2_X1   g654(.A(new_n855_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g655(.A1(new_n854_), .A2(new_n576_), .ZN(new_n857_));
  XOR2_X1   g656(.A(new_n857_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g657(.A1(new_n854_), .A2(new_n591_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT61), .B(G155gat), .Z(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1346gat));
  OAI21_X1  g660(.A(G162gat), .B1(new_n854_), .B2(new_n664_), .ZN(new_n862_));
  INV_X1    g661(.A(G162gat), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n624_), .A2(new_n863_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n862_), .B1(new_n854_), .B2(new_n864_), .ZN(G1347gat));
  AND2_X1   g664(.A1(new_n283_), .A2(new_n381_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n866_), .A2(KEYINPUT125), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n342_), .B1(new_n866_), .B2(KEYINPUT125), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n812_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n449_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G169gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n872_), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n870_), .A2(G169gat), .A3(new_n874_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n873_), .B(new_n875_), .C1(new_n219_), .C2(new_n870_), .ZN(G1348gat));
  NAND2_X1  g675(.A1(new_n869_), .A2(new_n575_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g677(.A1(new_n869_), .A2(new_n724_), .ZN(new_n879_));
  MUX2_X1   g678(.A(new_n223_), .B(G183gat), .S(new_n879_), .Z(G1350gat));
  INV_X1    g679(.A(new_n222_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n869_), .A2(new_n881_), .A3(new_n624_), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n869_), .A2(new_n665_), .ZN(new_n883_));
  INV_X1    g682(.A(G190gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(G1351gat));
  NOR4_X1   g684(.A1(new_n812_), .A2(new_n391_), .A3(new_n639_), .A4(new_n395_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n449_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n575_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g689(.A(KEYINPUT63), .ZN(new_n891_));
  INV_X1    g690(.A(G211gat), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n724_), .B1(new_n891_), .B2(new_n892_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n893_), .B(KEYINPUT127), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n886_), .A2(new_n894_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n891_), .A2(new_n892_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1354gat));
  INV_X1    g696(.A(G218gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n886_), .A2(new_n898_), .A3(new_n624_), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n886_), .A2(new_n665_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n898_), .ZN(G1355gat));
endmodule


