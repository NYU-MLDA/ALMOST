//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n784_,
    new_n785_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT27), .ZN(new_n203_));
  XNOR2_X1  g002(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G226gat), .A2(G233gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  OR2_X1    g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G197gat), .A2(G204gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT21), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(KEYINPUT21), .A3(new_n208_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G211gat), .B(G218gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n212_), .A3(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n212_), .A2(new_n213_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT25), .B(G183gat), .ZN(new_n218_));
  XNOR2_X1  g017(.A(KEYINPUT26), .B(G190gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT76), .ZN(new_n221_));
  INV_X1    g020(.A(G169gat), .ZN(new_n222_));
  INV_X1    g021(.A(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n221_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT76), .B1(G169gat), .B2(G176gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n224_), .A2(KEYINPUT24), .A3(new_n225_), .A4(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n220_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT23), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT78), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT78), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(KEYINPUT23), .ZN(new_n233_));
  AND2_X1   g032(.A1(G183gat), .A2(G190gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT81), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G183gat), .A2(G190gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT23), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT80), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n238_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT78), .B(KEYINPUT23), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(KEYINPUT81), .A3(new_n234_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n237_), .A2(new_n243_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT89), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n224_), .A2(new_n226_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT24), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n246_), .A2(new_n247_), .A3(new_n250_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n247_), .B1(new_n246_), .B2(new_n250_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n229_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n234_), .A2(new_n230_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n254_), .B1(new_n244_), .B2(new_n234_), .ZN(new_n255_));
  OR2_X1    g054(.A1(G183gat), .A2(G190gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT90), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT77), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n225_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(KEYINPUT77), .A2(G169gat), .A3(G176gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT79), .B(G176gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT22), .B(G169gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n262_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n257_), .A2(new_n258_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n258_), .B1(new_n257_), .B2(new_n265_), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n217_), .B1(new_n253_), .B2(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n224_), .A2(KEYINPUT24), .A3(new_n226_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(new_n262_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n273_), .A2(new_n255_), .A3(new_n220_), .A4(new_n250_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n246_), .A2(new_n256_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n263_), .A2(new_n264_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n262_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n274_), .B1(new_n275_), .B2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT20), .B1(new_n279_), .B2(new_n216_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n206_), .B1(new_n270_), .B2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n278_), .B1(new_n246_), .B2(new_n256_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n255_), .A2(new_n250_), .A3(new_n220_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(new_n272_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n216_), .B1(new_n282_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n206_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(KEYINPUT20), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n253_), .A2(new_n269_), .A3(new_n217_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G8gat), .B(G36gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT18), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G64gat), .B(G92gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n281_), .A2(new_n290_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n294_), .B1(new_n281_), .B2(new_n290_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n203_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n294_), .ZN(new_n299_));
  NOR3_X1   g098(.A1(new_n270_), .A2(new_n280_), .A3(new_n206_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n257_), .A2(new_n265_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n253_), .A2(new_n217_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT20), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n303_), .B1(new_n279_), .B2(new_n216_), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n286_), .B1(new_n302_), .B2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n299_), .B1(new_n300_), .B2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n306_), .A2(KEYINPUT27), .A3(new_n295_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n298_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G127gat), .B(G134gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G113gat), .B(G120gat), .ZN(new_n310_));
  AND2_X1   g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n309_), .A2(new_n310_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT83), .ZN(new_n314_));
  INV_X1    g113(.A(G155gat), .ZN(new_n315_));
  INV_X1    g114(.A(G162gat), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(KEYINPUT83), .B1(G155gat), .B2(G162gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT3), .ZN(new_n321_));
  INV_X1    g120(.A(G141gat), .ZN(new_n322_));
  INV_X1    g121(.A(G148gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G141gat), .A2(G148gat), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT2), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n324_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(KEYINPUT84), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT84), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n332_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n320_), .B1(new_n329_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n322_), .A2(new_n323_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n325_), .ZN(new_n337_));
  AND2_X1   g136(.A1(new_n317_), .A2(new_n318_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n319_), .A2(KEYINPUT1), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT1), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n340_), .A2(G155gat), .A3(G162gat), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n337_), .B1(new_n338_), .B2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n313_), .B1(new_n335_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n320_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n331_), .A2(new_n333_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n324_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(G127gat), .B(G134gat), .Z(new_n349_));
  XOR2_X1   g148(.A(G113gat), .B(G120gat), .Z(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n309_), .A2(new_n310_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n317_), .A2(new_n339_), .A3(new_n341_), .A4(new_n318_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(new_n336_), .A3(new_n325_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n348_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(G225gat), .A2(G233gat), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n344_), .A2(new_n356_), .A3(new_n357_), .ZN(new_n358_));
  AND3_X1   g157(.A1(new_n344_), .A2(KEYINPUT4), .A3(new_n356_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n357_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(new_n344_), .B2(KEYINPUT4), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n358_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G1gat), .B(G29gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G57gat), .B(G85gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n363_), .B(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n367_), .ZN(new_n369_));
  OAI211_X1 g168(.A(new_n358_), .B(new_n369_), .C1(new_n359_), .C2(new_n361_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT87), .B(G106gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT29), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n373_), .B1(new_n348_), .B2(new_n355_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G78gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n375_), .A2(new_n376_), .A3(new_n216_), .ZN(new_n377_));
  OAI21_X1  g176(.A(G78gat), .B1(new_n374_), .B2(new_n217_), .ZN(new_n378_));
  AND2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n216_), .A2(KEYINPUT86), .ZN(new_n380_));
  INV_X1    g179(.A(G228gat), .ZN(new_n381_));
  INV_X1    g180(.A(G233gat), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G22gat), .B(G50gat), .Z(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n380_), .A2(new_n384_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT86), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n214_), .B2(new_n215_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n385_), .B1(new_n389_), .B2(new_n383_), .ZN(new_n390_));
  XOR2_X1   g189(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n391_));
  NAND2_X1  g190(.A1(new_n348_), .A2(new_n355_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n391_), .B1(new_n392_), .B2(KEYINPUT29), .ZN(new_n393_));
  INV_X1    g192(.A(new_n391_), .ZN(new_n394_));
  NAND4_X1  g193(.A1(new_n348_), .A2(new_n373_), .A3(new_n355_), .A4(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n387_), .A2(new_n390_), .A3(new_n393_), .A4(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n387_), .A2(new_n390_), .B1(new_n393_), .B2(new_n395_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n379_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n387_), .A2(new_n390_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n393_), .A2(new_n395_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n377_), .A2(new_n378_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n396_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n372_), .B1(new_n399_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n399_), .A2(new_n372_), .A3(new_n404_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n371_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n294_), .A2(KEYINPUT32), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n246_), .A2(new_n250_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(KEYINPUT89), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n246_), .A2(new_n247_), .A3(new_n250_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n228_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n268_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n266_), .ZN(new_n415_));
  NOR3_X1   g214(.A1(new_n413_), .A2(new_n415_), .A3(new_n216_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n409_), .B1(new_n416_), .B2(new_n287_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n216_), .B1(new_n413_), .B2(new_n415_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n282_), .A2(new_n284_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n303_), .B1(new_n419_), .B2(new_n217_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n286_), .B1(new_n418_), .B2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n371_), .B1(new_n417_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n418_), .A2(new_n420_), .A3(new_n286_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n217_), .A2(new_n301_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n413_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n285_), .A2(KEYINPUT20), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n206_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n409_), .B1(new_n423_), .B2(new_n427_), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT94), .B1(new_n422_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n409_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n431_), .A2(new_n281_), .B1(new_n370_), .B2(new_n368_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n430_), .B1(new_n300_), .B2(new_n305_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT94), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT92), .B1(new_n344_), .B2(new_n356_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n436_), .A2(new_n357_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n344_), .A2(KEYINPUT92), .A3(new_n356_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n369_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n353_), .B1(new_n348_), .B2(new_n355_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT4), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n360_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT93), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n344_), .A2(KEYINPUT4), .A3(new_n356_), .ZN(new_n444_));
  AND3_X1   g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n443_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n370_), .A2(KEYINPUT33), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n444_), .B(new_n360_), .C1(KEYINPUT4), .C2(new_n344_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT33), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n449_), .A2(new_n450_), .A3(new_n358_), .A4(new_n369_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n439_), .A2(new_n447_), .B1(new_n448_), .B2(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n413_), .A2(new_n415_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n287_), .B1(new_n453_), .B2(new_n217_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n299_), .B1(new_n421_), .B2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n455_), .A3(new_n295_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n429_), .A2(new_n435_), .A3(new_n456_), .ZN(new_n457_));
  AND3_X1   g256(.A1(new_n399_), .A2(new_n372_), .A3(new_n404_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n458_), .A2(new_n405_), .ZN(new_n459_));
  AOI22_X1  g258(.A1(new_n308_), .A2(new_n408_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G71gat), .B(G99gat), .ZN(new_n461_));
  INV_X1    g260(.A(G43gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n419_), .B(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(G227gat), .A2(G233gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n465_), .B(G15gat), .Z(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT30), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT31), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n464_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n464_), .A2(new_n468_), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT82), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n471_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT82), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n473_), .A2(new_n474_), .A3(new_n469_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n472_), .A2(new_n475_), .A3(new_n313_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n313_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT95), .B1(new_n460_), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n298_), .A2(new_n459_), .A3(new_n307_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT96), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT96), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n298_), .A2(new_n459_), .A3(new_n482_), .A4(new_n307_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NOR3_X1   g283(.A1(new_n476_), .A2(new_n477_), .A3(new_n371_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n457_), .A2(new_n459_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n408_), .A2(new_n298_), .A3(new_n307_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT95), .ZN(new_n490_));
  INV_X1    g289(.A(new_n478_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n479_), .A2(new_n486_), .A3(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(G232gat), .A2(G233gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT34), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT35), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT72), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n495_), .A2(KEYINPUT35), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G85gat), .B(G92gat), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n500_), .A2(KEYINPUT65), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G99gat), .A2(G106gat), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT6), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n502_), .B(new_n503_), .ZN(new_n504_));
  OR3_X1    g303(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n505_));
  OAI21_X1  g304(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n505_), .A2(new_n506_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n501_), .B1(new_n504_), .B2(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n508_), .A2(KEYINPUT8), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n508_), .A2(KEYINPUT8), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT10), .B(G99gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n511_), .B(KEYINPUT64), .ZN(new_n512_));
  INV_X1    g311(.A(G106gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT9), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n500_), .A2(new_n515_), .ZN(new_n516_));
  AND3_X1   g315(.A1(new_n515_), .A2(G85gat), .A3(G92gat), .ZN(new_n517_));
  NOR3_X1   g316(.A1(new_n516_), .A2(new_n504_), .A3(new_n517_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n509_), .A2(new_n510_), .B1(new_n514_), .B2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G29gat), .B(G36gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G43gat), .B(G50gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n520_), .B(new_n521_), .ZN(new_n522_));
  AOI211_X1 g321(.A(new_n498_), .B(new_n499_), .C1(new_n519_), .C2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n514_), .A2(new_n518_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n510_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n508_), .A2(KEYINPUT8), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n524_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n522_), .B(KEYINPUT15), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n529_), .A2(KEYINPUT70), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(KEYINPUT70), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n523_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n496_), .A2(new_n497_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n529_), .B(KEYINPUT70), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(new_n533_), .A3(new_n523_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G190gat), .B(G218gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT71), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G134gat), .B(G162gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT36), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n535_), .A2(new_n537_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n541_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n544_), .A2(KEYINPUT36), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n546_), .B1(new_n535_), .B2(new_n537_), .ZN(new_n547_));
  OAI21_X1  g346(.A(KEYINPUT100), .B1(new_n543_), .B2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n535_), .A2(new_n537_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n545_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT100), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n535_), .A2(new_n537_), .A3(new_n542_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n548_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(new_n493_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT12), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n524_), .B(new_n557_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n559_), .A2(KEYINPUT11), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(KEYINPUT11), .ZN(new_n561_));
  XOR2_X1   g360(.A(G71gat), .B(G78gat), .Z(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n561_), .A2(new_n562_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT66), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT12), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n558_), .B(new_n566_), .C1(new_n519_), .C2(new_n568_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n527_), .A2(new_n567_), .A3(KEYINPUT12), .A4(new_n565_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G230gat), .A2(G233gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n572_), .B1(new_n527_), .B2(new_n565_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n574_), .B1(new_n565_), .B2(new_n527_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  XOR2_X1   g375(.A(KEYINPUT67), .B(KEYINPUT5), .Z(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT68), .ZN(new_n578_));
  XNOR2_X1  g377(.A(G120gat), .B(G148gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G176gat), .B(G204gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n576_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n573_), .A2(new_n575_), .A3(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n586_), .B1(KEYINPUT69), .B2(KEYINPUT13), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT69), .B(KEYINPUT13), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n583_), .A2(new_n585_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G15gat), .B(G22gat), .ZN(new_n592_));
  INV_X1    g391(.A(G8gat), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G1gat), .B(G8gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(new_n522_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G229gat), .A2(G233gat), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n528_), .A2(new_n601_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n600_), .B1(new_n597_), .B2(new_n522_), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n598_), .A2(new_n600_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(G113gat), .B(G141gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(G169gat), .B(G197gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n604_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n604_), .A2(new_n607_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G127gat), .B(G155gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT16), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G183gat), .B(G211gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT17), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT73), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n597_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(new_n566_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n615_), .A2(KEYINPUT17), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n617_), .B(new_n620_), .C1(new_n567_), .C2(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(KEYINPUT66), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n620_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n622_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n591_), .A2(new_n611_), .A3(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n556_), .A2(new_n627_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n202_), .B1(new_n628_), .B2(new_n371_), .ZN(new_n629_));
  OR2_X1    g428(.A1(new_n629_), .A2(KEYINPUT101), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(KEYINPUT101), .ZN(new_n631_));
  INV_X1    g430(.A(new_n611_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n493_), .A2(new_n632_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n625_), .B(KEYINPUT74), .ZN(new_n634_));
  OAI21_X1  g433(.A(KEYINPUT37), .B1(new_n543_), .B2(new_n547_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT37), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n550_), .A2(new_n636_), .A3(new_n552_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n634_), .A2(new_n638_), .A3(new_n590_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT75), .Z(new_n640_));
  NAND2_X1  g439(.A1(new_n633_), .A2(new_n640_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n641_), .A2(KEYINPUT97), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(KEYINPUT97), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n642_), .A2(new_n202_), .A3(new_n371_), .A4(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n645_));
  AOI22_X1  g444(.A1(new_n630_), .A2(new_n631_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n644_), .A2(new_n645_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n647_), .A2(KEYINPUT99), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT99), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n644_), .A2(new_n649_), .A3(new_n645_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n646_), .B1(new_n648_), .B2(new_n650_), .ZN(G1324gat));
  INV_X1    g450(.A(KEYINPUT39), .ZN(new_n652_));
  INV_X1    g451(.A(new_n308_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n628_), .A2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n654_), .B2(G8gat), .ZN(new_n655_));
  AOI211_X1 g454(.A(KEYINPUT39), .B(new_n593_), .C1(new_n628_), .C2(new_n653_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n642_), .A2(new_n643_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n653_), .A2(new_n593_), .ZN(new_n658_));
  OAI22_X1  g457(.A1(new_n655_), .A2(new_n656_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(G1325gat));
  NAND2_X1  g460(.A1(new_n628_), .A2(new_n478_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(G15gat), .ZN(new_n663_));
  XOR2_X1   g462(.A(new_n663_), .B(KEYINPUT41), .Z(new_n664_));
  OR2_X1    g463(.A1(new_n491_), .A2(G15gat), .ZN(new_n665_));
  OR3_X1    g464(.A1(new_n657_), .A2(KEYINPUT102), .A3(new_n665_), .ZN(new_n666_));
  OAI21_X1  g465(.A(KEYINPUT102), .B1(new_n657_), .B2(new_n665_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n664_), .A2(new_n666_), .A3(new_n667_), .ZN(G1326gat));
  INV_X1    g467(.A(G22gat), .ZN(new_n669_));
  INV_X1    g468(.A(new_n459_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n669_), .B1(new_n628_), .B2(new_n670_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT42), .Z(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n669_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n657_), .B2(new_n673_), .ZN(G1327gat));
  OAI21_X1  g473(.A(KEYINPUT106), .B1(new_n555_), .B2(new_n634_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT74), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n625_), .B(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT106), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n677_), .A2(new_n554_), .A3(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n591_), .B1(new_n675_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n633_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(G29gat), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n371_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n677_), .A2(new_n590_), .A3(new_n632_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n638_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(KEYINPUT103), .A2(KEYINPUT43), .ZN(new_n688_));
  AND3_X1   g487(.A1(new_n493_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n689_));
  XOR2_X1   g488(.A(KEYINPUT103), .B(KEYINPUT43), .Z(new_n690_));
  AOI21_X1  g489(.A(new_n690_), .B1(new_n493_), .B2(new_n687_), .ZN(new_n691_));
  OAI211_X1 g490(.A(KEYINPUT44), .B(new_n686_), .C1(new_n689_), .C2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n492_), .A2(new_n486_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n490_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n687_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n690_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n695_), .A2(new_n696_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n493_), .A2(new_n687_), .A3(new_n688_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n685_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n699_), .A2(KEYINPUT104), .A3(KEYINPUT44), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT104), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n686_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n371_), .B(new_n692_), .C1(new_n700_), .C2(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(KEYINPUT105), .B1(new_n705_), .B2(G29gat), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n692_), .A2(new_n371_), .ZN(new_n707_));
  OAI21_X1  g506(.A(KEYINPUT104), .B1(new_n699_), .B2(KEYINPUT44), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n702_), .A2(new_n701_), .A3(new_n703_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n710_), .A2(new_n711_), .A3(new_n683_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n684_), .B1(new_n706_), .B2(new_n712_), .ZN(G1328gat));
  OR2_X1    g512(.A1(new_n653_), .A2(KEYINPUT107), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n653_), .A2(KEYINPUT107), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n717_), .A2(G36gat), .ZN(new_n718_));
  INV_X1    g517(.A(new_n718_), .ZN(new_n719_));
  OR3_X1    g518(.A1(new_n681_), .A2(KEYINPUT45), .A3(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(KEYINPUT45), .B1(new_n681_), .B2(new_n719_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n692_), .A2(new_n653_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n724_));
  INV_X1    g523(.A(G36gat), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n722_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT46), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT46), .B(new_n722_), .C1(new_n724_), .C2(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(G1329gat));
  NOR2_X1   g529(.A1(new_n491_), .A2(new_n462_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n692_), .B(new_n731_), .C1(new_n700_), .C2(new_n704_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n462_), .B1(new_n681_), .B2(new_n491_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1330gat));
  AOI21_X1  g536(.A(G50gat), .B1(new_n682_), .B2(new_n670_), .ZN(new_n738_));
  AOI22_X1  g537(.A1(new_n708_), .A2(new_n709_), .B1(KEYINPUT44), .B2(new_n699_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n670_), .A2(G50gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n739_), .B2(new_n740_), .ZN(G1331gat));
  INV_X1    g540(.A(G57gat), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n591_), .A2(new_n611_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n556_), .A2(new_n634_), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n742_), .B1(new_n747_), .B2(new_n371_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n493_), .A2(new_n611_), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n687_), .A2(new_n677_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(new_n591_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n371_), .ZN(new_n752_));
  NOR3_X1   g551(.A1(new_n751_), .A2(G57gat), .A3(new_n752_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n748_), .A2(new_n753_), .ZN(G1332gat));
  OR3_X1    g553(.A1(new_n751_), .A2(G64gat), .A3(new_n717_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n747_), .A2(new_n716_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(KEYINPUT110), .B(KEYINPUT48), .ZN(new_n757_));
  AND3_X1   g556(.A1(new_n756_), .A2(G64gat), .A3(new_n757_), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n757_), .B1(new_n756_), .B2(G64gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(G1333gat));
  OR3_X1    g559(.A1(new_n751_), .A2(G71gat), .A3(new_n491_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n747_), .A2(new_n478_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT49), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n762_), .A2(new_n763_), .A3(G71gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n762_), .B2(G71gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(G1334gat));
  INV_X1    g565(.A(KEYINPUT50), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n747_), .A2(new_n670_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(G78gat), .ZN(new_n769_));
  AOI211_X1 g568(.A(KEYINPUT50), .B(new_n376_), .C1(new_n747_), .C2(new_n670_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n670_), .A2(new_n376_), .ZN(new_n771_));
  OAI22_X1  g570(.A1(new_n769_), .A2(new_n770_), .B1(new_n751_), .B2(new_n771_), .ZN(G1335gat));
  NOR2_X1   g571(.A1(new_n689_), .A2(new_n691_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT111), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n743_), .A2(new_n634_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n776_), .B1(new_n689_), .B2(new_n691_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n774_), .A2(new_n775_), .A3(new_n777_), .ZN(new_n778_));
  OAI21_X1  g577(.A(G85gat), .B1(new_n778_), .B2(new_n752_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n675_), .A2(new_n679_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n749_), .A2(new_n591_), .A3(new_n780_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n752_), .A2(G85gat), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n779_), .B1(new_n781_), .B2(new_n782_), .ZN(G1336gat));
  OAI21_X1  g582(.A(G92gat), .B1(new_n778_), .B2(new_n717_), .ZN(new_n784_));
  OR2_X1    g583(.A1(new_n308_), .A2(G92gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n784_), .B1(new_n781_), .B2(new_n785_), .ZN(G1337gat));
  OAI21_X1  g585(.A(G99gat), .B1(new_n778_), .B2(new_n491_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n781_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n788_), .A2(new_n478_), .A3(new_n512_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n791_), .A2(KEYINPUT112), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n787_), .B(new_n789_), .C1(KEYINPUT112), .C2(new_n791_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(G1338gat));
  XNOR2_X1  g594(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n513_), .B1(KEYINPUT113), .B2(KEYINPUT52), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n775_), .A2(new_n670_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n773_), .B2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(KEYINPUT113), .A2(KEYINPUT52), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n788_), .A2(new_n513_), .A3(new_n670_), .ZN(new_n802_));
  AND2_X1   g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  OR2_X1    g602(.A1(new_n799_), .A2(new_n800_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n796_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  AND4_X1   g604(.A1(new_n804_), .A2(new_n801_), .A3(new_n802_), .A4(new_n796_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(new_n806_), .ZN(G1339gat));
  XNOR2_X1  g606(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n750_), .A2(new_n611_), .A3(new_n590_), .A4(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n808_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n639_), .B2(new_n632_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(KEYINPUT58), .ZN(new_n814_));
  INV_X1    g613(.A(new_n572_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n569_), .A2(new_n815_), .A3(new_n570_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT116), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT116), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n569_), .A2(new_n818_), .A3(new_n815_), .A4(new_n570_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n817_), .A2(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(KEYINPUT55), .B1(new_n571_), .B2(new_n572_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822_));
  AOI211_X1 g621(.A(new_n822_), .B(new_n815_), .C1(new_n569_), .C2(new_n570_), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n584_), .B1(new_n820_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT56), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n599_), .B1(new_n597_), .B2(new_n522_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n602_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n607_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n609_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n827_), .A2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n585_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n814_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n585_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n573_), .A2(new_n822_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n571_), .A2(KEYINPUT55), .A3(new_n572_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(new_n817_), .A4(new_n819_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n582_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n835_), .B1(new_n839_), .B2(KEYINPUT56), .ZN(new_n840_));
  INV_X1    g639(.A(new_n814_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n840_), .A2(new_n831_), .A3(new_n827_), .A4(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n834_), .A2(new_n687_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT117), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n611_), .B1(new_n839_), .B2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n825_), .A2(KEYINPUT117), .A3(new_n826_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n840_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n586_), .A2(new_n831_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n844_), .B1(new_n850_), .B2(new_n555_), .ZN(new_n851_));
  AOI211_X1 g650(.A(KEYINPUT57), .B(new_n554_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n843_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n812_), .B1(new_n853_), .B2(new_n626_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n491_), .A2(new_n752_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n855_), .A2(new_n484_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n854_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(G113gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n858_), .A2(new_n859_), .A3(new_n632_), .ZN(new_n860_));
  OAI21_X1  g659(.A(KEYINPUT59), .B1(new_n854_), .B2(new_n857_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n812_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n843_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n849_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n632_), .B1(new_n825_), .B2(KEYINPUT117), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n833_), .A2(new_n865_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n866_), .B2(new_n847_), .ZN(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT57), .B1(new_n867_), .B2(new_n554_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n850_), .A2(new_n844_), .A3(new_n555_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n863_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n862_), .B1(new_n870_), .B2(new_n634_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT59), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n856_), .B2(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n874_), .B1(new_n873_), .B2(new_n856_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT120), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n861_), .A2(new_n876_), .A3(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n877_), .B1(new_n861_), .B2(new_n876_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n878_), .A2(new_n879_), .A3(new_n611_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n860_), .B1(new_n880_), .B2(new_n859_), .ZN(G1340gat));
  INV_X1    g680(.A(G120gat), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(new_n590_), .B2(KEYINPUT60), .ZN(new_n883_));
  OAI211_X1 g682(.A(new_n858_), .B(new_n883_), .C1(KEYINPUT60), .C2(new_n882_), .ZN(new_n884_));
  AND3_X1   g683(.A1(new_n861_), .A2(new_n876_), .A3(new_n591_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n882_), .ZN(G1341gat));
  INV_X1    g685(.A(G127gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n858_), .A2(new_n887_), .A3(new_n634_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n878_), .A2(new_n879_), .A3(new_n626_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n889_), .B2(new_n887_), .ZN(G1342gat));
  AOI21_X1  g689(.A(G134gat), .B1(new_n858_), .B2(new_n554_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n878_), .A2(new_n879_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n687_), .A2(G134gat), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(KEYINPUT121), .Z(new_n894_));
  AOI21_X1  g693(.A(new_n891_), .B1(new_n892_), .B2(new_n894_), .ZN(G1343gat));
  NAND4_X1  g694(.A1(new_n717_), .A2(new_n491_), .A3(new_n371_), .A4(new_n670_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT122), .Z(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n854_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n632_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n591_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g701(.A1(new_n898_), .A2(new_n634_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G155gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  AOI21_X1  g704(.A(G162gat), .B1(new_n898_), .B2(new_n554_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n638_), .A2(new_n316_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT123), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n906_), .B1(new_n898_), .B2(new_n908_), .ZN(G1347gat));
  AOI21_X1  g708(.A(new_n812_), .B1(new_n853_), .B2(new_n677_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n485_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n717_), .A2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n459_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n910_), .A2(new_n611_), .A3(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT124), .ZN(new_n915_));
  OAI21_X1  g714(.A(G169gat), .B1(new_n914_), .B2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n914_), .A2(new_n915_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n917_), .A2(KEYINPUT62), .A3(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT62), .ZN(new_n920_));
  INV_X1    g719(.A(new_n918_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n921_), .B2(new_n916_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n914_), .A2(new_n264_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n919_), .A2(new_n922_), .A3(new_n923_), .ZN(G1348gat));
  NOR2_X1   g723(.A1(new_n910_), .A2(new_n913_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n591_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n854_), .A2(new_n670_), .ZN(new_n927_));
  NOR4_X1   g726(.A1(new_n717_), .A2(new_n223_), .A3(new_n911_), .A4(new_n590_), .ZN(new_n928_));
  AOI22_X1  g727(.A1(new_n926_), .A2(new_n263_), .B1(new_n927_), .B2(new_n928_), .ZN(G1349gat));
  INV_X1    g728(.A(new_n218_), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n925_), .A2(new_n930_), .A3(new_n625_), .ZN(new_n931_));
  AND3_X1   g730(.A1(new_n927_), .A2(new_n634_), .A3(new_n912_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n932_), .B2(G183gat), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  OAI211_X1 g734(.A(KEYINPUT125), .B(new_n931_), .C1(new_n932_), .C2(G183gat), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(G1350gat));
  NAND2_X1  g736(.A1(new_n554_), .A2(new_n219_), .ZN(new_n938_));
  XOR2_X1   g737(.A(new_n938_), .B(KEYINPUT126), .Z(new_n939_));
  NAND2_X1  g738(.A1(new_n925_), .A2(new_n939_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n910_), .A2(new_n638_), .A3(new_n913_), .ZN(new_n941_));
  INV_X1    g740(.A(G190gat), .ZN(new_n942_));
  OAI21_X1  g741(.A(new_n940_), .B1(new_n941_), .B2(new_n942_), .ZN(G1351gat));
  INV_X1    g742(.A(new_n854_), .ZN(new_n944_));
  AND3_X1   g743(.A1(new_n716_), .A2(new_n491_), .A3(new_n408_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n944_), .A2(new_n945_), .ZN(new_n946_));
  INV_X1    g745(.A(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n632_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n948_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g748(.A1(new_n946_), .A2(new_n590_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT127), .ZN(new_n951_));
  AND2_X1   g750(.A1(new_n951_), .A2(G204gat), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n951_), .A2(G204gat), .ZN(new_n953_));
  OAI21_X1  g752(.A(new_n950_), .B1(new_n952_), .B2(new_n953_), .ZN(new_n954_));
  OAI21_X1  g753(.A(new_n954_), .B1(new_n950_), .B2(new_n953_), .ZN(G1353gat));
  AOI211_X1 g754(.A(KEYINPUT63), .B(G211gat), .C1(new_n947_), .C2(new_n625_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(KEYINPUT63), .B(G211gat), .ZN(new_n957_));
  NOR3_X1   g756(.A1(new_n946_), .A2(new_n626_), .A3(new_n957_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n956_), .A2(new_n958_), .ZN(G1354gat));
  OR3_X1    g758(.A1(new_n946_), .A2(G218gat), .A3(new_n555_), .ZN(new_n960_));
  OAI21_X1  g759(.A(G218gat), .B1(new_n946_), .B2(new_n638_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1355gat));
endmodule


