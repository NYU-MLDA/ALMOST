//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 1 0 1 0 1 1 1 0 1 1 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:07 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n624_,
    new_n625_, new_n626_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n830_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n885_, new_n886_,
    new_n887_;
  XOR2_X1   g000(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n205_), .B(KEYINPUT81), .Z(new_n206_));
  NOR2_X1   g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(KEYINPUT80), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT80), .ZN(new_n209_));
  NOR3_X1   g008(.A1(new_n209_), .A2(G155gat), .A3(G162gat), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n204_), .A2(KEYINPUT1), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n206_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  INV_X1    g014(.A(G141gat), .ZN(new_n216_));
  INV_X1    g015(.A(G148gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT84), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n216_), .A2(new_n217_), .A3(KEYINPUT3), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(G141gat), .B2(G148gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n215_), .A2(KEYINPUT82), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT2), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n215_), .A2(KEYINPUT82), .A3(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n224_), .A2(new_n226_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT83), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND4_X1  g030(.A1(new_n224_), .A2(new_n226_), .A3(KEYINPUT83), .A4(new_n228_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n204_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n220_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  AOI211_X1 g035(.A(KEYINPUT84), .B(new_n234_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n219_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT85), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT85), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n240_), .B(new_n219_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT29), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n203_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  AOI211_X1 g043(.A(KEYINPUT29), .B(new_n202_), .C1(new_n239_), .C2(new_n241_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n239_), .A2(KEYINPUT29), .A3(new_n241_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT21), .ZN(new_n248_));
  INV_X1    g047(.A(G204gat), .ZN(new_n249_));
  OR2_X1    g048(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(KEYINPUT87), .A2(G197gat), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(G197gat), .A2(G204gat), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n248_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G211gat), .B(G218gat), .Z(new_n255_));
  NAND3_X1  g054(.A1(new_n250_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n248_), .B1(G197gat), .B2(G204gat), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n255_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n255_), .A2(KEYINPUT21), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n252_), .A2(new_n253_), .ZN(new_n260_));
  AOI22_X1  g059(.A1(new_n254_), .A2(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n261_), .B1(G228gat), .B2(G233gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n247_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n258_), .A2(new_n254_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n259_), .A2(new_n260_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  AND3_X1   g065(.A1(new_n214_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n233_), .A2(new_n235_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT84), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n233_), .A2(new_n220_), .A3(new_n235_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n267_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n266_), .B1(new_n271_), .B2(new_n243_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n272_), .A2(G228gat), .A3(G233gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G78gat), .B(G106gat), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n263_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n274_), .B1(new_n263_), .B2(new_n273_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n246_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n263_), .A2(new_n273_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n274_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n263_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n242_), .A2(new_n243_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(new_n202_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n242_), .A2(new_n243_), .A3(new_n203_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n280_), .A2(new_n281_), .A3(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G22gat), .B(G50gat), .ZN(new_n287_));
  XOR2_X1   g086(.A(new_n287_), .B(KEYINPUT88), .Z(new_n288_));
  AND3_X1   g087(.A1(new_n277_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n288_), .B1(new_n277_), .B2(new_n286_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G1gat), .B(G29gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT94), .B(G85gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT0), .B(G57gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n294_), .B(new_n295_), .Z(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G225gat), .A2(G233gat), .ZN(new_n298_));
  XOR2_X1   g097(.A(new_n298_), .B(KEYINPUT93), .Z(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G127gat), .B(G134gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G113gat), .B(G120gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT79), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n301_), .B(new_n302_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n305_), .B1(new_n306_), .B2(new_n304_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n239_), .A2(new_n241_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n271_), .A2(new_n306_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT4), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT4), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n308_), .A2(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n300_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n308_), .A2(new_n298_), .A3(new_n309_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT95), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND4_X1  g116(.A1(new_n308_), .A2(KEYINPUT95), .A3(new_n298_), .A4(new_n309_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n297_), .B1(new_n314_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n313_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n312_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n299_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n323_), .A2(new_n296_), .A3(new_n317_), .A4(new_n318_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n320_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G64gat), .B(G92gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT92), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G8gat), .B(G36gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT32), .ZN(new_n332_));
  OAI21_X1  g131(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n333_));
  NOR3_X1   g132(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G183gat), .ZN(new_n336_));
  INV_X1    g135(.A(G190gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT23), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(G183gat), .A3(G190gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(KEYINPUT78), .A3(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n342_), .B(KEYINPUT23), .C1(new_n336_), .C2(new_n337_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n333_), .B(new_n335_), .C1(new_n344_), .C2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT26), .B(G190gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT25), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n347_), .B1(new_n348_), .B2(G183gat), .ZN(new_n349_));
  AND2_X1   g148(.A1(new_n348_), .A2(KEYINPUT76), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n348_), .A2(KEYINPUT76), .ZN(new_n351_));
  OAI21_X1  g150(.A(G183gat), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT77), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT77), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n354_), .B(G183gat), .C1(new_n350_), .C2(new_n351_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n349_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  AND2_X1   g155(.A1(new_n338_), .A2(new_n340_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NOR3_X1   g157(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n359_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n358_), .A2(new_n363_), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n261_), .B(new_n346_), .C1(new_n356_), .C2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT20), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n335_), .A2(KEYINPUT89), .A3(new_n333_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT89), .ZN(new_n368_));
  INV_X1    g167(.A(new_n333_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(new_n334_), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n367_), .B(new_n370_), .C1(new_n357_), .C2(new_n345_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT25), .B(G183gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n347_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n363_), .A2(new_n373_), .A3(new_n341_), .A4(new_n343_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n366_), .B1(new_n266_), .B2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G226gat), .A2(G233gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT19), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n365_), .A2(new_n376_), .A3(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n346_), .B1(new_n356_), .B2(new_n364_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n266_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT96), .B(KEYINPUT20), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n385_), .B1(new_n266_), .B2(new_n375_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n378_), .B1(new_n383_), .B2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n332_), .B1(new_n380_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT90), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(new_n266_), .B2(new_n375_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n378_), .A2(new_n366_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n261_), .A2(KEYINPUT90), .A3(new_n371_), .A4(new_n374_), .ZN(new_n392_));
  AND4_X1   g191(.A1(new_n382_), .A2(new_n390_), .A3(new_n391_), .A4(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n379_), .B1(new_n365_), .B2(new_n376_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n388_), .B1(new_n395_), .B2(new_n332_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n325_), .A2(new_n396_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n314_), .A2(new_n319_), .ZN(new_n398_));
  AOI21_X1  g197(.A(KEYINPUT33), .B1(new_n398_), .B2(new_n296_), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n329_), .B(new_n330_), .Z(new_n400_));
  OAI21_X1  g199(.A(new_n400_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n394_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n382_), .A2(new_n390_), .A3(new_n391_), .A4(new_n392_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n402_), .A2(new_n331_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n298_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n310_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n296_), .B1(new_n407_), .B2(new_n299_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n405_), .B1(new_n406_), .B2(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n296_), .A2(KEYINPUT33), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n323_), .A2(new_n317_), .A3(new_n318_), .A4(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n291_), .B(new_n397_), .C1(new_n399_), .C2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G227gat), .A2(G233gat), .ZN(new_n414_));
  INV_X1    g213(.A(G15gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n416_), .B(KEYINPUT30), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n381_), .B(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(new_n418_), .B(new_n307_), .Z(new_n419_));
  XNOR2_X1  g218(.A(G71gat), .B(G99gat), .ZN(new_n420_));
  INV_X1    g219(.A(G43gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT31), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n419_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n288_), .ZN(new_n426_));
  NOR3_X1   g225(.A1(new_n275_), .A2(new_n276_), .A3(new_n246_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n285_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n426_), .B1(new_n427_), .B2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n277_), .A2(new_n286_), .A3(new_n288_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT27), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT98), .B1(new_n405_), .B2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT98), .ZN(new_n434_));
  AOI211_X1 g233(.A(new_n434_), .B(KEYINPUT27), .C1(new_n401_), .C2(new_n404_), .ZN(new_n435_));
  OR2_X1    g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  OR2_X1    g235(.A1(new_n404_), .A2(KEYINPUT97), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n404_), .A2(KEYINPUT97), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n387_), .A2(new_n380_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n432_), .B1(new_n439_), .B2(new_n400_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n437_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n320_), .A2(new_n436_), .A3(new_n324_), .A4(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n425_), .B1(new_n431_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n441_), .B1(new_n433_), .B2(new_n435_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT99), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT99), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n441_), .B(new_n446_), .C1(new_n433_), .C2(new_n435_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n448_), .A2(new_n430_), .A3(new_n429_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n325_), .A2(new_n424_), .ZN(new_n450_));
  AOI22_X1  g249(.A1(new_n413_), .A2(new_n443_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(KEYINPUT10), .B(G99gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(KEYINPUT64), .ZN(new_n453_));
  INV_X1    g252(.A(G106gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G99gat), .A2(G106gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT6), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT6), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n458_), .A2(G99gat), .A3(G106gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G85gat), .A2(G92gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n460_), .B1(KEYINPUT9), .B2(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G85gat), .B(G92gat), .Z(new_n463_));
  AOI21_X1  g262(.A(new_n462_), .B1(KEYINPUT9), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n455_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT68), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT8), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT65), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n460_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n457_), .A2(new_n459_), .A3(KEYINPUT65), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT66), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT66), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(new_n474_), .A3(new_n471_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G99gat), .A2(G106gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT7), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n473_), .A2(new_n475_), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n468_), .B1(new_n478_), .B2(new_n463_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n463_), .A2(new_n468_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n480_), .B1(new_n460_), .B2(new_n477_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n467_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G29gat), .B(G36gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G43gat), .B(G50gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT15), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n482_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT71), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n482_), .A2(KEYINPUT71), .A3(new_n486_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT72), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G232gat), .A2(G233gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT34), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n494_), .B2(KEYINPUT35), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n465_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT67), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OAI211_X1 g297(.A(KEYINPUT67), .B(new_n465_), .C1(new_n479_), .C2(new_n481_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n495_), .B1(new_n500_), .B2(new_n485_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n491_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n494_), .A2(KEYINPUT35), .ZN(new_n503_));
  XOR2_X1   g302(.A(new_n503_), .B(KEYINPUT70), .Z(new_n504_));
  NAND2_X1  g303(.A1(new_n502_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n504_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n491_), .A2(new_n506_), .A3(new_n501_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G190gat), .B(G218gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G134gat), .B(G162gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(new_n510_), .B(KEYINPUT36), .Z(new_n511_));
  AND3_X1   g310(.A1(new_n505_), .A2(new_n507_), .A3(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(new_n510_), .A2(KEYINPUT36), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n513_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n451_), .A2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G57gat), .B(G64gat), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n517_), .A2(KEYINPUT11), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(KEYINPUT11), .ZN(new_n519_));
  XOR2_X1   g318(.A(G71gat), .B(G78gat), .Z(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n519_), .A2(new_n520_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G15gat), .B(G22gat), .ZN(new_n524_));
  INV_X1    g323(.A(G1gat), .ZN(new_n525_));
  INV_X1    g324(.A(G8gat), .ZN(new_n526_));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n524_), .A2(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G1gat), .B(G8gat), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n528_), .B(new_n529_), .Z(new_n530_));
  XNOR2_X1  g329(.A(new_n523_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G231gat), .A2(G233gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535_));
  XOR2_X1   g334(.A(G127gat), .B(G155gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT16), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n537_), .B(new_n538_), .ZN(new_n539_));
  OR3_X1    g338(.A1(new_n534_), .A2(new_n535_), .A3(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(KEYINPUT17), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n534_), .A2(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n530_), .A2(new_n485_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT73), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n545_), .B1(new_n485_), .B2(new_n530_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G229gat), .A2(G233gat), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n530_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n486_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n545_), .A2(new_n547_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT74), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n545_), .A2(KEYINPUT74), .A3(new_n547_), .A4(new_n551_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n549_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  XOR2_X1   g355(.A(G113gat), .B(G141gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT75), .ZN(new_n558_));
  XOR2_X1   g357(.A(G169gat), .B(G197gat), .Z(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n556_), .B(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n523_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n523_), .A2(KEYINPUT12), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n500_), .A2(new_n562_), .B1(new_n482_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(new_n500_), .B2(new_n562_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G230gat), .A2(G233gat), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n565_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n500_), .A2(new_n562_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n523_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  XOR2_X1   g372(.A(G120gat), .B(G148gat), .Z(new_n574_));
  XNOR2_X1  g373(.A(G176gat), .B(G204gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  NAND3_X1  g377(.A1(new_n569_), .A2(new_n573_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n578_), .B1(new_n569_), .B2(new_n573_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT13), .Z(new_n583_));
  NAND4_X1  g382(.A1(new_n516_), .A2(new_n543_), .A3(new_n561_), .A4(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT100), .Z(new_n585_));
  INV_X1    g384(.A(new_n325_), .ZN(new_n586_));
  OAI21_X1  g385(.A(G1gat), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n583_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT37), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n505_), .A2(new_n507_), .A3(new_n511_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n505_), .A2(new_n507_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n589_), .B(new_n590_), .C1(new_n591_), .C2(new_n513_), .ZN(new_n592_));
  OAI21_X1  g391(.A(KEYINPUT37), .B1(new_n512_), .B2(new_n514_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n543_), .ZN(new_n596_));
  NOR3_X1   g395(.A1(new_n588_), .A2(new_n595_), .A3(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(new_n561_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n451_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n525_), .A3(new_n325_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT38), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n587_), .A2(new_n603_), .ZN(G1324gat));
  INV_X1    g403(.A(new_n448_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(new_n526_), .A3(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n584_), .A2(new_n448_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n526_), .B1(new_n607_), .B2(KEYINPUT101), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT101), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n610_), .B1(new_n584_), .B2(new_n448_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n608_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n609_), .B1(new_n608_), .B2(new_n611_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n606_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT40), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OAI211_X1 g415(.A(KEYINPUT40), .B(new_n606_), .C1(new_n612_), .C2(new_n613_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n616_), .A2(new_n617_), .ZN(G1325gat));
  OAI21_X1  g417(.A(G15gat), .B1(new_n585_), .B2(new_n424_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT41), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n619_), .B(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n601_), .A2(new_n415_), .A3(new_n425_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1326gat));
  OAI21_X1  g422(.A(G22gat), .B1(new_n585_), .B2(new_n291_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT42), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n291_), .A2(G22gat), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n625_), .B1(new_n600_), .B2(new_n626_), .ZN(G1327gat));
  NAND2_X1  g426(.A1(new_n515_), .A2(new_n596_), .ZN(new_n628_));
  NOR4_X1   g427(.A1(new_n451_), .A2(new_n588_), .A3(new_n598_), .A4(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(G29gat), .B1(new_n629_), .B2(new_n325_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n442_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n631_));
  OAI211_X1 g430(.A(new_n430_), .B(new_n429_), .C1(new_n399_), .C2(new_n412_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n325_), .A2(new_n396_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n424_), .B(new_n631_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n449_), .A2(new_n450_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n594_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n637_));
  OAI21_X1  g436(.A(KEYINPUT103), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639_));
  INV_X1    g438(.A(new_n637_), .ZN(new_n640_));
  OAI211_X1 g439(.A(new_n639_), .B(new_n640_), .C1(new_n451_), .C2(new_n594_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT43), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n636_), .A2(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n638_), .A2(new_n641_), .A3(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n588_), .A2(new_n543_), .A3(new_n598_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(KEYINPUT44), .A3(new_n645_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n325_), .A2(G29gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n630_), .B1(new_n650_), .B2(new_n651_), .ZN(G1328gat));
  NAND3_X1  g451(.A1(new_n648_), .A2(new_n605_), .A3(new_n649_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(G36gat), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n448_), .A2(G36gat), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n629_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n655_), .B1(new_n629_), .B2(new_n656_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT105), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n659_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n654_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n660_), .A2(new_n661_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n663_), .B(new_n665_), .ZN(G1329gat));
  AOI21_X1  g465(.A(G43gat), .B1(new_n629_), .B2(new_n425_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n424_), .A2(new_n421_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n650_), .B2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT47), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(G1330gat));
  AOI21_X1  g470(.A(G50gat), .B1(new_n629_), .B2(new_n431_), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n431_), .A2(G50gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n672_), .B1(new_n650_), .B2(new_n673_), .ZN(G1331gat));
  NAND4_X1  g473(.A1(new_n516_), .A2(new_n543_), .A3(new_n598_), .A4(new_n588_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G57gat), .B1(new_n675_), .B2(new_n586_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n588_), .A2(new_n598_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n677_), .A2(new_n451_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n595_), .A2(new_n596_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT106), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n586_), .A2(G57gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n676_), .B1(new_n681_), .B2(new_n682_), .ZN(G1332gat));
  OAI21_X1  g482(.A(G64gat), .B1(new_n675_), .B2(new_n448_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT48), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n448_), .A2(G64gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n685_), .B1(new_n681_), .B2(new_n686_), .ZN(G1333gat));
  OAI21_X1  g486(.A(G71gat), .B1(new_n675_), .B2(new_n424_), .ZN(new_n688_));
  XOR2_X1   g487(.A(KEYINPUT107), .B(KEYINPUT49), .Z(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n424_), .A2(G71gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n681_), .B2(new_n691_), .ZN(G1334gat));
  OAI21_X1  g491(.A(G78gat), .B1(new_n675_), .B2(new_n291_), .ZN(new_n693_));
  XOR2_X1   g492(.A(KEYINPUT108), .B(KEYINPUT50), .Z(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n291_), .A2(G78gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n681_), .B2(new_n696_), .ZN(G1335gat));
  NOR3_X1   g496(.A1(new_n677_), .A2(new_n451_), .A3(new_n628_), .ZN(new_n698_));
  INV_X1    g497(.A(G85gat), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(new_n699_), .A3(new_n325_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n677_), .A2(new_n543_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n644_), .A2(new_n701_), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n702_), .A2(new_n325_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n700_), .B1(new_n703_), .B2(new_n699_), .ZN(G1336gat));
  NAND2_X1  g503(.A1(new_n702_), .A2(new_n605_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n448_), .A2(G92gat), .ZN(new_n706_));
  AOI22_X1  g505(.A1(new_n705_), .A2(G92gat), .B1(new_n698_), .B2(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT109), .Z(G1337gat));
  AND3_X1   g507(.A1(new_n698_), .A2(new_n425_), .A3(new_n453_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n702_), .A2(new_n425_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(G99gat), .ZN(new_n711_));
  XOR2_X1   g510(.A(new_n711_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g511(.A1(new_n698_), .A2(new_n454_), .A3(new_n431_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT52), .ZN(new_n714_));
  NAND4_X1  g513(.A1(new_n644_), .A2(KEYINPUT110), .A3(new_n431_), .A4(new_n701_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(G106gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n644_), .A2(new_n431_), .A3(new_n701_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT110), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n714_), .B1(new_n716_), .B2(new_n719_), .ZN(new_n720_));
  AND4_X1   g519(.A1(new_n714_), .A2(new_n719_), .A3(G106gat), .A4(new_n715_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n713_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT53), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT53), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n724_), .B(new_n713_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1339gat));
  INV_X1    g525(.A(KEYINPUT119), .ZN(new_n727_));
  INV_X1    g526(.A(G113gat), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n729_));
  NAND4_X1  g528(.A1(new_n679_), .A2(new_n598_), .A3(new_n583_), .A4(new_n729_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n583_), .A2(new_n543_), .A3(new_n598_), .A4(new_n594_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n729_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n730_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT118), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n546_), .A2(new_n547_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n545_), .A2(new_n548_), .A3(new_n551_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(new_n560_), .A3(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT113), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n556_), .A2(new_n560_), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n579_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n565_), .A2(new_n567_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT55), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n570_), .B2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n578_), .B1(new_n743_), .B2(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n744_), .B2(new_n570_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n565_), .A2(new_n567_), .A3(new_n748_), .ZN(new_n749_));
  AND3_X1   g548(.A1(new_n747_), .A2(KEYINPUT56), .A3(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(KEYINPUT56), .B1(new_n747_), .B2(new_n749_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n750_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n751_), .A2(KEYINPUT114), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n742_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT58), .B1(new_n756_), .B2(KEYINPUT115), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n743_), .A2(new_n746_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n578_), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(new_n749_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n753_), .B1(new_n760_), .B2(KEYINPUT56), .ZN(new_n761_));
  INV_X1    g560(.A(new_n750_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n761_), .A2(new_n755_), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n742_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT115), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT58), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n757_), .A2(new_n767_), .A3(new_n595_), .ZN(new_n768_));
  AND2_X1   g567(.A1(new_n561_), .A2(new_n579_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n769_), .B1(new_n750_), .B2(new_n751_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n741_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n515_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(KEYINPUT57), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT57), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n774_), .B(new_n515_), .C1(new_n770_), .C2(new_n771_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n773_), .A2(new_n775_), .ZN(new_n776_));
  AOI211_X1 g575(.A(new_n735_), .B(new_n543_), .C1(new_n768_), .C2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n595_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n778_));
  NOR3_X1   g577(.A1(new_n756_), .A2(KEYINPUT115), .A3(KEYINPUT58), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n776_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT118), .B1(new_n780_), .B2(new_n596_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n734_), .B1(new_n777_), .B2(new_n781_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n449_), .A2(new_n325_), .A3(new_n425_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT117), .ZN(new_n784_));
  XOR2_X1   g583(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n785_));
  NOR2_X1   g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n783_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n543_), .B1(new_n768_), .B2(new_n776_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n730_), .A2(new_n733_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n787_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  AOI22_X1  g589(.A1(new_n782_), .A2(new_n786_), .B1(KEYINPUT59), .B2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n728_), .B1(new_n791_), .B2(new_n561_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n790_), .A2(G113gat), .A3(new_n598_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n727_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n790_), .A2(KEYINPUT59), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n780_), .A2(new_n596_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n735_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n788_), .A2(KEYINPUT118), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n789_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n786_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n795_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  OAI21_X1  g600(.A(G113gat), .B1(new_n801_), .B2(new_n598_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n793_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(KEYINPUT119), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n794_), .A2(new_n804_), .ZN(G1340gat));
  OAI21_X1  g604(.A(G120gat), .B1(new_n801_), .B2(new_n583_), .ZN(new_n806_));
  INV_X1    g605(.A(G120gat), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n583_), .B2(KEYINPUT60), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(KEYINPUT60), .B2(new_n807_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n806_), .B1(new_n790_), .B2(new_n809_), .ZN(G1341gat));
  INV_X1    g609(.A(G127gat), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n811_), .B1(new_n791_), .B2(new_n543_), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n790_), .A2(G127gat), .A3(new_n596_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT120), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(G127gat), .B1(new_n801_), .B2(new_n596_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n816_));
  INV_X1    g615(.A(new_n813_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n814_), .A2(new_n818_), .ZN(G1342gat));
  INV_X1    g618(.A(new_n790_), .ZN(new_n820_));
  AOI21_X1  g619(.A(G134gat), .B1(new_n820_), .B2(new_n515_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n595_), .A2(G134gat), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT121), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(new_n791_), .B2(new_n823_), .ZN(G1343gat));
  AOI211_X1 g623(.A(new_n291_), .B(new_n425_), .C1(new_n796_), .C2(new_n734_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n605_), .A2(new_n586_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(new_n598_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(new_n216_), .ZN(G1344gat));
  NOR2_X1   g628(.A1(new_n827_), .A2(new_n583_), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(new_n217_), .ZN(G1345gat));
  NOR2_X1   g630(.A1(new_n827_), .A2(new_n596_), .ZN(new_n832_));
  XOR2_X1   g631(.A(KEYINPUT61), .B(G155gat), .Z(new_n833_));
  XNOR2_X1  g632(.A(new_n832_), .B(new_n833_), .ZN(G1346gat));
  INV_X1    g633(.A(new_n827_), .ZN(new_n835_));
  AOI21_X1  g634(.A(G162gat), .B1(new_n835_), .B2(new_n515_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n595_), .A2(G162gat), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT122), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n836_), .B1(new_n835_), .B2(new_n838_), .ZN(G1347gat));
  INV_X1    g638(.A(G169gat), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n448_), .A2(new_n325_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n425_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n431_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n844_), .A2(new_n598_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n840_), .B1(new_n782_), .B2(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  OR3_X1    g647(.A1(new_n846_), .A2(KEYINPUT124), .A3(new_n848_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(KEYINPUT22), .B(G169gat), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n782_), .A2(new_n845_), .A3(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n846_), .A2(KEYINPUT124), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n848_), .B1(new_n846_), .B2(KEYINPUT124), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n849_), .B(new_n851_), .C1(new_n852_), .C2(new_n853_), .ZN(G1348gat));
  NOR2_X1   g653(.A1(new_n799_), .A2(new_n844_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G176gat), .B1(new_n855_), .B2(new_n588_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n431_), .B1(new_n796_), .B2(new_n734_), .ZN(new_n857_));
  INV_X1    g656(.A(G176gat), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n583_), .A2(new_n858_), .A3(new_n842_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n856_), .B1(new_n857_), .B2(new_n859_), .ZN(G1349gat));
  NOR2_X1   g659(.A1(new_n842_), .A2(new_n596_), .ZN(new_n861_));
  AOI21_X1  g660(.A(G183gat), .B1(new_n857_), .B2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n596_), .A2(new_n372_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n855_), .B2(new_n863_), .ZN(G1350gat));
  NAND3_X1  g663(.A1(new_n855_), .A2(new_n347_), .A3(new_n515_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n855_), .A2(new_n595_), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT125), .B1(new_n866_), .B2(G190gat), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT125), .ZN(new_n868_));
  AOI211_X1 g667(.A(new_n868_), .B(new_n337_), .C1(new_n855_), .C2(new_n595_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n865_), .B1(new_n867_), .B2(new_n869_), .ZN(G1351gat));
  NAND2_X1  g669(.A1(new_n825_), .A2(new_n841_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n561_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G197gat), .ZN(G1352gat));
  NOR2_X1   g673(.A1(new_n871_), .A2(new_n583_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(new_n249_), .ZN(G1353gat));
  NOR2_X1   g675(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT127), .ZN(new_n878_));
  NOR3_X1   g677(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n879_));
  NAND2_X1  g678(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n543_), .A2(new_n880_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(KEYINPUT126), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n871_), .A2(new_n882_), .ZN(new_n883_));
  MUX2_X1   g682(.A(new_n878_), .B(new_n879_), .S(new_n883_), .Z(G1354gat));
  OAI21_X1  g683(.A(G218gat), .B1(new_n871_), .B2(new_n594_), .ZN(new_n885_));
  INV_X1    g684(.A(G218gat), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n515_), .A2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n885_), .B1(new_n871_), .B2(new_n887_), .ZN(G1355gat));
endmodule


