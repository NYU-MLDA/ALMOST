//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n754_,
    new_n755_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n916_, new_n917_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n937_, new_n938_, new_n939_, new_n940_, new_n941_,
    new_n942_, new_n943_, new_n945_, new_n946_, new_n948_, new_n949_,
    new_n950_, new_n952_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n959_, new_n960_, new_n961_;
  XOR2_X1   g000(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G190gat), .B(G218gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G134gat), .B(G162gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT36), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G232gat), .A2(G233gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(KEYINPUT34), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(KEYINPUT35), .ZN(new_n210_));
  OR2_X1    g009(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(KEYINPUT64), .A3(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n214_));
  AND2_X1   g013(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n214_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(G106gat), .B1(new_n213_), .B2(new_n217_), .ZN(new_n218_));
  OR2_X1    g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n219_), .A2(KEYINPUT9), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G99gat), .A2(G106gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT6), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(G99gat), .A3(G106gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n223_), .A2(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n220_), .A2(KEYINPUT9), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n221_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n218_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n219_), .A2(new_n220_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n223_), .A2(new_n225_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT7), .ZN(new_n233_));
  INV_X1    g032(.A(G99gat), .ZN(new_n234_));
  INV_X1    g033(.A(G106gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n231_), .B1(new_n232_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT8), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n224_), .B1(G99gat), .B2(G106gat), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n237_), .B(new_n236_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT8), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(new_n231_), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n229_), .B1(new_n240_), .B2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G29gat), .B(G36gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G43gat), .B(G50gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n210_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n251_));
  INV_X1    g050(.A(new_n237_), .ZN(new_n252_));
  NOR3_X1   g051(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  AOI211_X1 g053(.A(KEYINPUT8), .B(new_n230_), .C1(new_n254_), .C2(new_n226_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n244_), .B1(new_n243_), .B2(new_n231_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n251_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n240_), .A2(KEYINPUT67), .A3(new_n245_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n229_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT15), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n249_), .B(new_n260_), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n250_), .B(KEYINPUT72), .C1(new_n259_), .C2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT71), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n209_), .A2(KEYINPUT35), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n265_), .B(KEYINPUT70), .Z(new_n266_));
  OAI211_X1 g065(.A(new_n250_), .B(KEYINPUT71), .C1(new_n259_), .C2(new_n261_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n264_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n266_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n262_), .A2(new_n263_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n206_), .A2(KEYINPUT36), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n207_), .B1(new_n268_), .B2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n264_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n207_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n274_), .A2(new_n275_), .A3(new_n271_), .A4(new_n270_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n273_), .A2(KEYINPUT37), .A3(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(KEYINPUT37), .B1(new_n273_), .B2(new_n276_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G230gat), .A2(G233gat), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  NOR3_X1   g080(.A1(new_n215_), .A2(new_n216_), .A3(new_n214_), .ZN(new_n282_));
  AOI21_X1  g081(.A(KEYINPUT64), .B1(new_n211_), .B2(new_n212_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n235_), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n221_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n287_));
  XOR2_X1   g086(.A(G71gat), .B(G78gat), .Z(new_n288_));
  XNOR2_X1  g087(.A(G57gat), .B(G64gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n288_), .B1(KEYINPUT11), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT65), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n289_), .B2(KEYINPUT11), .ZN(new_n292_));
  INV_X1    g091(.A(G64gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(G57gat), .ZN(new_n294_));
  INV_X1    g093(.A(G57gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(G64gat), .ZN(new_n296_));
  AND4_X1   g095(.A1(new_n291_), .A2(new_n294_), .A3(new_n296_), .A4(KEYINPUT11), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n290_), .B1(new_n292_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n294_), .A2(new_n296_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT11), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT65), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n289_), .A2(new_n291_), .A3(KEYINPUT11), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n300_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n303_), .A4(new_n288_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n298_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n287_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n240_), .A2(new_n245_), .ZN(new_n307_));
  AOI22_X1  g106(.A1(new_n307_), .A2(new_n286_), .B1(new_n304_), .B2(new_n298_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n281_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT66), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(KEYINPUT66), .B(new_n281_), .C1(new_n306_), .C2(new_n308_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n280_), .B1(new_n287_), .B2(new_n305_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT68), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  OAI211_X1 g115(.A(KEYINPUT68), .B(new_n280_), .C1(new_n287_), .C2(new_n305_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT12), .B1(new_n287_), .B2(new_n305_), .ZN(new_n319_));
  NOR3_X1   g118(.A1(new_n255_), .A2(new_n256_), .A3(new_n251_), .ZN(new_n320_));
  AOI21_X1  g119(.A(KEYINPUT67), .B1(new_n240_), .B2(new_n245_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n286_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n305_), .A2(KEYINPUT12), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n319_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n318_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n313_), .A2(new_n326_), .ZN(new_n327_));
  XOR2_X1   g126(.A(G120gat), .B(G148gat), .Z(new_n328_));
  XNOR2_X1  g127(.A(G176gat), .B(G204gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n327_), .A2(new_n333_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n311_), .A2(new_n312_), .B1(new_n318_), .B2(new_n325_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(new_n332_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n334_), .A2(KEYINPUT13), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT13), .B1(new_n334_), .B2(new_n336_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G127gat), .B(G155gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT16), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G183gat), .B(G211gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n341_), .B(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT17), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n343_), .A2(new_n344_), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n298_), .A2(new_n304_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT73), .B(G15gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(G22gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(G1gat), .B(G8gat), .Z(new_n350_));
  INV_X1    g149(.A(G1gat), .ZN(new_n351_));
  INV_X1    g150(.A(G8gat), .ZN(new_n352_));
  OAI21_X1  g151(.A(KEYINPUT14), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(new_n350_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n350_), .B1(new_n349_), .B2(new_n353_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n347_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  AND2_X1   g156(.A1(new_n348_), .A2(G22gat), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n348_), .A2(G22gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n353_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n350_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n305_), .A2(new_n362_), .A3(new_n354_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(G231gat), .ZN(new_n365_));
  INV_X1    g164(.A(G233gat), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n364_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n365_), .A2(new_n366_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n357_), .A2(new_n368_), .A3(new_n363_), .ZN(new_n369_));
  AOI211_X1 g168(.A(new_n345_), .B(new_n346_), .C1(new_n367_), .C2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n367_), .A2(KEYINPUT74), .A3(new_n345_), .A4(new_n369_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n367_), .A2(new_n345_), .A3(new_n369_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT74), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n370_), .B1(new_n371_), .B2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT75), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n279_), .A2(new_n339_), .A3(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G127gat), .B(G134gat), .Z(new_n379_));
  XOR2_X1   g178(.A(G113gat), .B(G120gat), .Z(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G227gat), .A2(G233gat), .ZN(new_n382_));
  INV_X1    g181(.A(G71gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G99gat), .ZN(new_n385_));
  XOR2_X1   g184(.A(G15gat), .B(G43gat), .Z(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT79), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n385_), .B(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G183gat), .A2(G190gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT23), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  OR2_X1    g190(.A1(G183gat), .A2(G190gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT22), .ZN(new_n396_));
  INV_X1    g195(.A(G169gat), .ZN(new_n397_));
  INV_X1    g196(.A(G176gat), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n394_), .A2(new_n395_), .A3(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n397_), .A2(new_n398_), .A3(KEYINPUT78), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT78), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n402_), .B1(G169gat), .B2(G176gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT24), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(G169gat), .B2(G176gat), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n407_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n391_), .A2(new_n393_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n408_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT76), .ZN(new_n412_));
  INV_X1    g211(.A(G183gat), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n412_), .B1(new_n413_), .B2(KEYINPUT25), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(KEYINPUT25), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT25), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n416_), .A2(KEYINPUT76), .A3(G183gat), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n414_), .A2(new_n415_), .A3(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT26), .ZN(new_n419_));
  INV_X1    g218(.A(G190gat), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n419_), .B1(new_n420_), .B2(KEYINPUT77), .ZN(new_n421_));
  OR3_X1    g220(.A1(new_n419_), .A2(new_n420_), .A3(KEYINPUT77), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n418_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n400_), .B1(new_n411_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT30), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n409_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n422_), .A2(new_n421_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n427_), .B(new_n408_), .C1(new_n428_), .C2(new_n418_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n429_), .A2(KEYINPUT30), .A3(new_n400_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT80), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n426_), .A2(new_n430_), .A3(KEYINPUT80), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n388_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n388_), .ZN(new_n436_));
  AOI21_X1  g235(.A(KEYINPUT80), .B1(new_n426_), .B2(new_n430_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT31), .B1(new_n435_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n434_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n436_), .B1(new_n440_), .B2(new_n437_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT31), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n433_), .A2(new_n388_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT81), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n439_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n445_), .B1(new_n439_), .B2(new_n444_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n381_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n439_), .A2(new_n444_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT81), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n379_), .B(new_n380_), .Z(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n452_), .A3(new_n446_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n449_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G1gat), .B(G29gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G57gat), .B(G85gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G225gat), .A2(G233gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G155gat), .ZN(new_n463_));
  INV_X1    g262(.A(G162gat), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT1), .B1(new_n463_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT1), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(G155gat), .A3(G162gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n463_), .A2(new_n464_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n465_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G141gat), .A2(G148gat), .ZN(new_n470_));
  INV_X1    g269(.A(G141gat), .ZN(new_n471_));
  INV_X1    g270(.A(G148gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n469_), .A2(new_n470_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT3), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n475_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT2), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n470_), .A2(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n476_), .A2(new_n478_), .A3(new_n479_), .A4(new_n480_), .ZN(new_n481_));
  XOR2_X1   g280(.A(G155gat), .B(G162gat), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n474_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT82), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT82), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n474_), .A2(new_n483_), .A3(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n485_), .A2(new_n487_), .A3(new_n452_), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n462_), .B1(new_n488_), .B2(KEYINPUT4), .ZN(new_n489_));
  INV_X1    g288(.A(new_n484_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n381_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n488_), .A2(KEYINPUT4), .A3(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT94), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n488_), .A2(KEYINPUT94), .A3(KEYINPUT4), .A4(new_n491_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n489_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n488_), .A2(new_n491_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n497_), .A2(new_n461_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n460_), .B1(new_n496_), .B2(new_n498_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n496_), .A2(new_n498_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(new_n459_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G78gat), .B(G106gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT87), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT29), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n474_), .A2(new_n483_), .A3(new_n486_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n486_), .B1(new_n474_), .B2(new_n483_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT28), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n485_), .A2(new_n487_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT28), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(new_n505_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G22gat), .B(G50gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n509_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n514_), .B1(new_n509_), .B2(new_n512_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n504_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n509_), .A2(new_n512_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n513_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n502_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n509_), .A2(new_n512_), .A3(new_n514_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  NOR2_X1   g321(.A1(G197gat), .A2(G204gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT85), .B(G197gat), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n523_), .B1(new_n524_), .B2(G204gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G211gat), .B(G218gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(KEYINPUT21), .A3(new_n527_), .ZN(new_n528_));
  NOR2_X1   g327(.A1(new_n524_), .A2(G204gat), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT21), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n530_), .B1(G197gat), .B2(G204gat), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n526_), .B1(new_n529_), .B2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n525_), .A2(KEYINPUT21), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n528_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(KEYINPUT83), .A2(G233gat), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  NOR2_X1   g336(.A1(KEYINPUT83), .A2(G233gat), .ZN(new_n538_));
  OAI21_X1  g337(.A(G228gat), .B1(new_n537_), .B2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT84), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n535_), .B(new_n540_), .C1(new_n510_), .C2(new_n505_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT86), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n535_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(KEYINPUT86), .B(new_n528_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n490_), .A2(new_n505_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n541_), .B1(new_n547_), .B2(new_n539_), .ZN(new_n548_));
  AND3_X1   g347(.A1(new_n517_), .A2(new_n522_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n517_), .B2(new_n522_), .ZN(new_n550_));
  OAI211_X1 g349(.A(new_n499_), .B(new_n501_), .C1(new_n549_), .C2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT27), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n553_));
  NAND2_X1  g352(.A1(G226gat), .A2(G233gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT20), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n535_), .B2(new_n424_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n399_), .A2(new_n395_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT90), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT90), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n399_), .A2(new_n561_), .A3(new_n395_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT92), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n391_), .A2(new_n392_), .A3(new_n565_), .A4(new_n393_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n394_), .A2(KEYINPUT91), .ZN(new_n567_));
  NAND4_X1  g366(.A1(new_n563_), .A2(new_n564_), .A3(new_n566_), .A4(new_n567_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n567_), .A2(new_n560_), .A3(new_n566_), .A4(new_n562_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT92), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n416_), .A2(G183gat), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n415_), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n573_), .B(KEYINPUT89), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT26), .B(G190gat), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n411_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n577_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n556_), .B(new_n558_), .C1(new_n578_), .C2(new_n535_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT20), .B1(new_n535_), .B2(new_n424_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n580_), .B1(new_n578_), .B2(new_n535_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n579_), .B1(new_n581_), .B2(new_n556_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G8gat), .B(G36gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G64gat), .B(G92gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n582_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n587_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n535_), .A2(new_n424_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n576_), .B1(new_n570_), .B2(new_n568_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n535_), .ZN(new_n592_));
  OAI211_X1 g391(.A(KEYINPUT20), .B(new_n590_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(new_n555_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n589_), .B1(new_n594_), .B2(new_n579_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n552_), .B1(new_n588_), .B2(new_n595_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n543_), .A2(new_n577_), .A3(new_n569_), .A4(new_n544_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n556_), .B1(new_n597_), .B2(new_n558_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n581_), .A2(new_n556_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n601_), .A2(new_n587_), .ZN(new_n602_));
  AND2_X1   g401(.A1(new_n558_), .A2(new_n556_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n591_), .A2(new_n592_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n593_), .A2(new_n555_), .B1(new_n603_), .B2(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n552_), .B1(new_n605_), .B2(new_n589_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n602_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n596_), .A2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT97), .B1(new_n551_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n582_), .A2(new_n587_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n594_), .A2(new_n589_), .A3(new_n579_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  AOI22_X1  g411(.A1(new_n612_), .A2(new_n552_), .B1(new_n602_), .B2(new_n606_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n550_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n517_), .A2(new_n522_), .A3(new_n548_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n501_), .A2(new_n499_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n613_), .A2(new_n616_), .A3(new_n618_), .A4(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n609_), .A2(new_n620_), .ZN(new_n621_));
  AOI21_X1  g420(.A(KEYINPUT33), .B1(new_n500_), .B2(new_n459_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n612_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n500_), .A2(KEYINPUT33), .A3(new_n459_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n459_), .B1(new_n497_), .B2(new_n462_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n494_), .A2(new_n495_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n461_), .B1(new_n488_), .B2(KEYINPUT4), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n626_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .A4(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n589_), .A2(KEYINPUT32), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n631_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n501_), .B2(new_n499_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n605_), .A2(new_n631_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT96), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT96), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n605_), .A2(new_n636_), .A3(new_n631_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n633_), .A2(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n616_), .B1(new_n630_), .B2(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n454_), .B1(new_n621_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n616_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(new_n613_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n449_), .A2(new_n453_), .A3(new_n618_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n643_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n641_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT98), .ZN(new_n648_));
  NAND2_X1  g447(.A1(G229gat), .A2(G233gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n362_), .A2(new_n354_), .A3(new_n249_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n249_), .B1(new_n362_), .B2(new_n354_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n650_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n355_), .A2(new_n356_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n651_), .B(new_n649_), .C1(new_n655_), .C2(new_n261_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(G113gat), .B(G141gat), .ZN(new_n657_));
  XNOR2_X1  g456(.A(G169gat), .B(G197gat), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n657_), .B(new_n658_), .Z(new_n659_));
  AND3_X1   g458(.A1(new_n654_), .A2(new_n656_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n659_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n647_), .A2(new_n648_), .A3(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n629_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(new_n622_), .ZN(new_n666_));
  AOI22_X1  g465(.A1(new_n666_), .A2(new_n625_), .B1(new_n633_), .B2(new_n638_), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n609_), .B(new_n620_), .C1(new_n667_), .C2(new_n616_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n645_), .B1(new_n668_), .B2(new_n454_), .ZN(new_n669_));
  OAI21_X1  g468(.A(KEYINPUT98), .B1(new_n669_), .B2(new_n662_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n378_), .B1(new_n664_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n617_), .A2(new_n351_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n203_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n273_), .A2(KEYINPUT101), .A3(new_n276_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT101), .B1(new_n273_), .B2(new_n276_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n669_), .A2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n377_), .A2(new_n663_), .A3(new_n339_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT100), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n679_), .A2(new_n681_), .ZN(new_n682_));
  OAI21_X1  g481(.A(G1gat), .B1(new_n682_), .B2(new_n618_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n671_), .A2(new_n351_), .A3(new_n617_), .A4(new_n202_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n674_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT102), .ZN(G1324gat));
  OAI21_X1  g485(.A(G8gat), .B1(new_n682_), .B2(new_n613_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT39), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n671_), .A2(new_n352_), .A3(new_n608_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n688_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n690_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1325gat));
  INV_X1    g493(.A(G15gat), .ZN(new_n695_));
  INV_X1    g494(.A(new_n454_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n671_), .A2(new_n695_), .A3(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT105), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n679_), .A2(new_n696_), .A3(new_n681_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G15gat), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT41), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(KEYINPUT41), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(KEYINPUT104), .A3(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n698_), .A2(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(KEYINPUT104), .B1(new_n701_), .B2(new_n702_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n704_), .A2(new_n705_), .ZN(G1326gat));
  OAI21_X1  g505(.A(G22gat), .B1(new_n682_), .B2(new_n642_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT42), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n642_), .A2(G22gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n672_), .B2(new_n709_), .ZN(G1327gat));
  NOR2_X1   g509(.A1(new_n677_), .A2(new_n377_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n339_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n664_), .B2(new_n670_), .ZN(new_n713_));
  AOI21_X1  g512(.A(G29gat), .B1(new_n713_), .B2(new_n617_), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n337_), .A2(new_n338_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n715_), .A2(new_n377_), .A3(new_n662_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n717_));
  INV_X1    g516(.A(new_n279_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n647_), .B2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(KEYINPUT106), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n669_), .A2(new_n279_), .A3(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n716_), .B1(new_n719_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  OAI211_X1 g524(.A(KEYINPUT44), .B(new_n716_), .C1(new_n719_), .C2(new_n722_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n617_), .A2(G29gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n714_), .B1(new_n727_), .B2(new_n728_), .ZN(G1328gat));
  NAND3_X1  g528(.A1(new_n725_), .A2(new_n608_), .A3(new_n726_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G36gat), .ZN(new_n731_));
  NOR2_X1   g530(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n664_), .A2(new_n670_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n712_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n613_), .A2(G36gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n733_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  XOR2_X1   g535(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n737_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n713_), .A2(new_n735_), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n732_), .B1(new_n738_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT109), .Z(new_n743_));
  AND3_X1   g542(.A1(new_n731_), .A2(new_n741_), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n731_), .B2(new_n741_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1329gat));
  NAND4_X1  g545(.A1(new_n725_), .A2(G43gat), .A3(new_n696_), .A4(new_n726_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n713_), .A2(new_n696_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(G43gat), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT47), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n747_), .B(new_n751_), .C1(G43gat), .C2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1330gat));
  AOI21_X1  g552(.A(G50gat), .B1(new_n713_), .B2(new_n616_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n616_), .A2(G50gat), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n727_), .B2(new_n755_), .ZN(G1331gat));
  XNOR2_X1  g555(.A(new_n375_), .B(KEYINPUT75), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n757_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n715_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT110), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n669_), .A2(new_n663_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(G57gat), .B1(new_n763_), .B2(new_n617_), .ZN(new_n764_));
  NOR3_X1   g563(.A1(new_n757_), .A2(new_n339_), .A3(new_n663_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n679_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n618_), .A2(KEYINPUT111), .ZN(new_n768_));
  MUX2_X1   g567(.A(KEYINPUT111), .B(new_n768_), .S(G57gat), .Z(new_n769_));
  AOI21_X1  g568(.A(new_n764_), .B1(new_n767_), .B2(new_n769_), .ZN(G1332gat));
  OAI21_X1  g569(.A(G64gat), .B1(new_n766_), .B2(new_n613_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT48), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n763_), .A2(new_n293_), .A3(new_n608_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(G1333gat));
  OAI21_X1  g573(.A(G71gat), .B1(new_n766_), .B2(new_n454_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT49), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n763_), .A2(new_n383_), .A3(new_n696_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(G1334gat));
  OAI21_X1  g577(.A(G78gat), .B1(new_n766_), .B2(new_n642_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT50), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n642_), .A2(G78gat), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n780_), .B1(new_n762_), .B2(new_n781_), .ZN(G1335gat));
  AND3_X1   g581(.A1(new_n761_), .A2(new_n715_), .A3(new_n711_), .ZN(new_n783_));
  AOI21_X1  g582(.A(G85gat), .B1(new_n783_), .B2(new_n617_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n719_), .A2(new_n722_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n377_), .A2(new_n339_), .A3(new_n663_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n617_), .A2(G85gat), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT112), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n784_), .B1(new_n788_), .B2(new_n790_), .ZN(G1336gat));
  INV_X1    g590(.A(G92gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n783_), .A2(new_n792_), .A3(new_n608_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n785_), .A2(new_n613_), .A3(new_n787_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(new_n792_), .ZN(G1337gat));
  OAI211_X1 g594(.A(new_n783_), .B(new_n696_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n796_));
  NOR3_X1   g595(.A1(new_n785_), .A2(new_n454_), .A3(new_n787_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n796_), .B1(new_n797_), .B2(new_n234_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g598(.A1(new_n783_), .A2(new_n235_), .A3(new_n616_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n616_), .B(new_n786_), .C1(new_n719_), .C2(new_n722_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n801_), .A2(new_n802_), .A3(G106gat), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n801_), .B2(G106gat), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n800_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g605(.A1(new_n643_), .A2(new_n454_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n651_), .B(new_n650_), .C1(new_n655_), .C2(new_n261_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n659_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n660_), .B1(new_n808_), .B2(new_n811_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n313_), .A2(new_n326_), .A3(new_n332_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n332_), .B1(new_n313_), .B2(new_n326_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OAI211_X1 g616(.A(KEYINPUT114), .B(new_n812_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n662_), .B1(new_n335_), .B2(new_n332_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820_));
  INV_X1    g619(.A(new_n319_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n246_), .A2(new_n347_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n821_), .B(new_n822_), .C1(new_n259_), .C2(new_n323_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n326_), .A2(new_n820_), .B1(new_n281_), .B2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n318_), .A2(new_n325_), .A3(KEYINPUT55), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n332_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(KEYINPUT113), .A2(KEYINPUT56), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n819_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT68), .B1(new_n822_), .B2(new_n280_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n317_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n821_), .B1(new_n259_), .B2(new_n323_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n820_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n823_), .A2(new_n281_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n834_), .A2(new_n825_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837_));
  AND4_X1   g636(.A1(new_n829_), .A2(new_n836_), .A3(new_n837_), .A4(new_n333_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n817_), .B(new_n818_), .C1(new_n828_), .C2(new_n838_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n839_), .A2(KEYINPUT57), .A3(new_n677_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT57), .B1(new_n839_), .B2(new_n677_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n836_), .A2(new_n837_), .A3(new_n333_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n844_), .A2(new_n336_), .A3(new_n812_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n826_), .A2(new_n837_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n843_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT58), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT58), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n843_), .B(new_n849_), .C1(new_n845_), .C2(new_n846_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n848_), .A2(new_n718_), .A3(new_n850_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n377_), .B1(new_n842_), .B2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT54), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n758_), .A2(new_n853_), .A3(new_n662_), .A4(new_n339_), .ZN(new_n854_));
  OAI21_X1  g653(.A(KEYINPUT54), .B1(new_n378_), .B2(new_n663_), .ZN(new_n855_));
  AND2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n617_), .B(new_n807_), .C1(new_n852_), .C2(new_n856_), .ZN(new_n857_));
  NOR2_X1   g656(.A1(new_n857_), .A2(new_n662_), .ZN(new_n858_));
  OR3_X1    g657(.A1(new_n858_), .A2(KEYINPUT116), .A3(G113gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(KEYINPUT116), .B1(new_n858_), .B2(G113gat), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n857_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n839_), .A2(new_n677_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT57), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n839_), .A2(new_n677_), .A3(KEYINPUT57), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n851_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n757_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n854_), .A2(new_n855_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n870_), .A2(KEYINPUT59), .A3(new_n617_), .A4(new_n807_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n862_), .A2(new_n871_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n663_), .A2(G113gat), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n859_), .A2(new_n860_), .B1(new_n872_), .B2(new_n873_), .ZN(G1340gat));
  NOR2_X1   g673(.A1(new_n339_), .A2(KEYINPUT60), .ZN(new_n875_));
  INV_X1    g674(.A(G120gat), .ZN(new_n876_));
  MUX2_X1   g675(.A(KEYINPUT60), .B(new_n875_), .S(new_n876_), .Z(new_n877_));
  NAND4_X1  g676(.A1(new_n870_), .A2(new_n617_), .A3(new_n807_), .A4(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT117), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n618_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n881_), .A2(KEYINPUT117), .A3(new_n807_), .A4(new_n877_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n339_), .B1(new_n862_), .B2(new_n871_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n883_), .B1(new_n884_), .B2(new_n876_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT118), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT118), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n883_), .B(new_n887_), .C1(new_n884_), .C2(new_n876_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(G1341gat));
  INV_X1    g688(.A(new_n857_), .ZN(new_n890_));
  INV_X1    g689(.A(G127gat), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(new_n891_), .A3(new_n377_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n757_), .B1(new_n862_), .B2(new_n871_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n893_), .B2(new_n891_), .ZN(G1342gat));
  INV_X1    g693(.A(G134gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n890_), .A2(new_n895_), .A3(new_n678_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n279_), .B1(new_n862_), .B2(new_n871_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n896_), .B1(new_n897_), .B2(new_n895_), .ZN(G1343gat));
  NAND2_X1  g697(.A1(new_n870_), .A2(new_n617_), .ZN(new_n899_));
  NOR3_X1   g698(.A1(new_n696_), .A2(new_n608_), .A3(new_n642_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n899_), .A2(new_n901_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n663_), .ZN(new_n903_));
  XOR2_X1   g702(.A(KEYINPUT119), .B(G141gat), .Z(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1344gat));
  NAND2_X1  g704(.A1(new_n902_), .A2(new_n715_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT120), .B(G148gat), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1345gat));
  NAND3_X1  g707(.A1(new_n881_), .A2(new_n377_), .A3(new_n900_), .ZN(new_n909_));
  OR2_X1    g708(.A1(new_n909_), .A2(KEYINPUT121), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(KEYINPUT121), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT61), .B(G155gat), .ZN(new_n912_));
  AND3_X1   g711(.A1(new_n910_), .A2(new_n911_), .A3(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n910_), .B2(new_n911_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(new_n914_), .ZN(G1346gat));
  NAND4_X1  g714(.A1(new_n881_), .A2(new_n464_), .A3(new_n678_), .A4(new_n900_), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n899_), .A2(new_n279_), .A3(new_n901_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n917_), .B2(new_n464_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT122), .ZN(G1347gat));
  NOR2_X1   g718(.A1(new_n644_), .A2(new_n613_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT123), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n616_), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n870_), .A2(new_n922_), .A3(new_n396_), .A4(new_n663_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n923_), .A2(KEYINPUT62), .A3(new_n397_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n923_), .A2(KEYINPUT62), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n870_), .A2(new_n922_), .A3(new_n926_), .A4(new_n663_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(G169gat), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n924_), .B1(new_n925_), .B2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(KEYINPUT124), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT124), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n931_), .B(new_n924_), .C1(new_n925_), .C2(new_n928_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(G1348gat));
  NAND2_X1  g732(.A1(new_n870_), .A2(new_n922_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n339_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(new_n398_), .ZN(G1349gat));
  INV_X1    g735(.A(new_n934_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n574_), .B1(new_n938_), .B2(G183gat), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n937_), .A2(new_n377_), .A3(new_n939_), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n938_), .B(new_n413_), .C1(new_n934_), .C2(new_n757_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n940_), .A2(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT126), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n942_), .B(new_n943_), .ZN(G1350gat));
  OAI21_X1  g743(.A(G190gat), .B1(new_n934_), .B2(new_n279_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n678_), .A2(new_n575_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n945_), .B1(new_n934_), .B2(new_n946_), .ZN(G1351gat));
  NOR3_X1   g746(.A1(new_n696_), .A2(new_n613_), .A3(new_n551_), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n870_), .A2(new_n948_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n949_), .A2(new_n663_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g750(.A1(new_n949_), .A2(new_n715_), .ZN(new_n952_));
  XNOR2_X1  g751(.A(new_n952_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g752(.A1(new_n949_), .A2(new_n377_), .ZN(new_n954_));
  NOR2_X1   g753(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n955_));
  AND2_X1   g754(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n956_));
  NOR3_X1   g755(.A1(new_n954_), .A2(new_n955_), .A3(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n957_), .B1(new_n954_), .B2(new_n955_), .ZN(G1354gat));
  AOI21_X1  g757(.A(G218gat), .B1(new_n949_), .B2(new_n678_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n718_), .A2(G218gat), .ZN(new_n960_));
  XOR2_X1   g759(.A(new_n960_), .B(KEYINPUT127), .Z(new_n961_));
  AOI21_X1  g760(.A(new_n959_), .B1(new_n949_), .B2(new_n961_), .ZN(G1355gat));
endmodule


