//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n563_,
    new_n564_, new_n565_, new_n566_, new_n567_, new_n568_, new_n569_,
    new_n570_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n671_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n819_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n843_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n858_, new_n859_, new_n860_;
  XOR2_X1   g000(.A(G29gat), .B(G36gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT15), .Z(new_n205_));
  XNOR2_X1  g004(.A(G15gat), .B(G22gat), .ZN(new_n206_));
  INV_X1    g005(.A(G1gat), .ZN(new_n207_));
  INV_X1    g006(.A(G8gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT14), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G1gat), .B(G8gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n205_), .A2(new_n212_), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n212_), .A2(new_n204_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G229gat), .A2(G233gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n212_), .B(new_n204_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n215_), .ZN(new_n218_));
  AOI22_X1  g017(.A1(new_n213_), .A2(new_n216_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(G113gat), .B(G141gat), .Z(new_n220_));
  XNOR2_X1  g019(.A(G169gat), .B(G197gat), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n220_), .B(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n219_), .A2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n219_), .A2(new_n222_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G227gat), .A2(G233gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT77), .ZN(new_n227_));
  XOR2_X1   g026(.A(G71gat), .B(G99gat), .Z(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G15gat), .B(G43gat), .ZN(new_n230_));
  XNOR2_X1  g029(.A(KEYINPUT76), .B(KEYINPUT78), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n230_), .B(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n229_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT22), .B(G169gat), .ZN(new_n234_));
  INV_X1    g033(.A(G176gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G169gat), .A2(G176gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT74), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n236_), .A2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  INV_X1    g039(.A(G183gat), .ZN(new_n241_));
  INV_X1    g040(.A(G190gat), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT23), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT23), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n244_), .A2(G183gat), .A3(G190gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n243_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n239_), .B1(new_n240_), .B2(new_n247_), .ZN(new_n248_));
  OR2_X1    g047(.A1(G169gat), .A2(G176gat), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n238_), .A2(KEYINPUT24), .A3(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT25), .B(G183gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT26), .B(G190gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n250_), .B(new_n253_), .C1(KEYINPUT24), .C2(new_n249_), .ZN(new_n254_));
  XOR2_X1   g053(.A(new_n245_), .B(KEYINPUT75), .Z(new_n255_));
  AND2_X1   g054(.A1(new_n255_), .A2(new_n243_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n248_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(KEYINPUT30), .Z(new_n258_));
  AND2_X1   g057(.A1(new_n258_), .A2(KEYINPUT79), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(KEYINPUT79), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n233_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n261_), .B1(new_n259_), .B2(new_n233_), .ZN(new_n262_));
  XOR2_X1   g061(.A(G127gat), .B(G134gat), .Z(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(KEYINPUT80), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G113gat), .B(G120gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n266_), .B(KEYINPUT31), .Z(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n262_), .A2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n262_), .A2(new_n268_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G155gat), .A2(G162gat), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n273_), .A2(KEYINPUT1), .ZN(new_n274_));
  NOR2_X1   g073(.A1(G155gat), .A2(G162gat), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n273_), .B1(new_n275_), .B2(KEYINPUT1), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT81), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n274_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(new_n277_), .B2(new_n276_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G141gat), .A2(G148gat), .ZN(new_n280_));
  INV_X1    g079(.A(G141gat), .ZN(new_n281_));
  INV_X1    g080(.A(G148gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n279_), .A2(new_n280_), .A3(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G155gat), .B(G162gat), .Z(new_n285_));
  XNOR2_X1  g084(.A(new_n285_), .B(KEYINPUT84), .ZN(new_n286_));
  NAND3_X1  g085(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT83), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n281_), .A2(new_n282_), .A3(KEYINPUT82), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT2), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n289_), .A2(KEYINPUT3), .B1(new_n290_), .B2(new_n280_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n288_), .B(new_n291_), .C1(KEYINPUT3), .C2(new_n289_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n286_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n284_), .A2(new_n293_), .ZN(new_n294_));
  AND2_X1   g093(.A1(new_n294_), .A2(KEYINPUT29), .ZN(new_n295_));
  INV_X1    g094(.A(G204gat), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(KEYINPUT86), .A3(G197gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G197gat), .B(G204gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  OAI211_X1 g098(.A(KEYINPUT21), .B(new_n297_), .C1(new_n299_), .C2(KEYINPUT86), .ZN(new_n300_));
  XOR2_X1   g099(.A(G211gat), .B(G218gat), .Z(new_n301_));
  INV_X1    g100(.A(KEYINPUT21), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n301_), .B1(new_n302_), .B2(new_n298_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n298_), .A2(new_n302_), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n300_), .A2(new_n303_), .B1(new_n301_), .B2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n295_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(G228gat), .A2(G233gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n305_), .B(KEYINPUT87), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(new_n307_), .ZN(new_n309_));
  OAI22_X1  g108(.A1(new_n306_), .A2(new_n307_), .B1(new_n309_), .B2(new_n295_), .ZN(new_n310_));
  XOR2_X1   g109(.A(G78gat), .B(G106gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n294_), .A2(KEYINPUT29), .ZN(new_n313_));
  XOR2_X1   g112(.A(G22gat), .B(G50gat), .Z(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  XOR2_X1   g114(.A(KEYINPUT85), .B(KEYINPUT28), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  OR2_X1    g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n312_), .A2(new_n317_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n318_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n272_), .A2(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(G1gat), .B(G29gat), .Z(new_n323_));
  XNOR2_X1  g122(.A(G57gat), .B(G85gat), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n326_));
  XOR2_X1   g125(.A(new_n325_), .B(new_n326_), .Z(new_n327_));
  INV_X1    g126(.A(new_n294_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(new_n266_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT4), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT4), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n266_), .A2(new_n331_), .A3(new_n294_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n330_), .A2(new_n332_), .ZN(new_n333_));
  AND2_X1   g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NOR2_X1   g134(.A1(new_n329_), .A2(new_n334_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n327_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT33), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n327_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n329_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n341_), .A2(KEYINPUT98), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT98), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n334_), .B1(new_n329_), .B2(new_n343_), .ZN(new_n344_));
  OAI221_X1 g143(.A(new_n340_), .B1(new_n342_), .B2(new_n344_), .C1(new_n334_), .C2(new_n333_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n337_), .A2(new_n338_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n339_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT95), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT20), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n308_), .B2(new_n257_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G226gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT90), .B(KEYINPUT24), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n355_), .A2(new_n249_), .ZN(new_n356_));
  AND3_X1   g155(.A1(new_n356_), .A2(new_n246_), .A3(new_n253_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n237_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT91), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT91), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n355_), .A2(new_n360_), .A3(new_n237_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n249_), .A3(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n357_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT92), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n239_), .B(KEYINPUT93), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(new_n240_), .B2(new_n256_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n305_), .ZN(new_n368_));
  OAI211_X1 g167(.A(new_n350_), .B(new_n354_), .C1(new_n365_), .C2(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n364_), .A2(new_n367_), .ZN(new_n370_));
  OAI221_X1 g169(.A(KEYINPUT20), .B1(new_n257_), .B2(new_n308_), .C1(new_n370_), .C2(new_n305_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT94), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n353_), .B(KEYINPUT89), .Z(new_n373_));
  AND3_X1   g172(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n372_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n369_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G8gat), .B(G36gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT18), .ZN(new_n378_));
  XNOR2_X1  g177(.A(G64gat), .B(G92gat), .ZN(new_n379_));
  XOR2_X1   g178(.A(new_n378_), .B(new_n379_), .Z(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n348_), .B1(new_n376_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n371_), .A2(new_n373_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT94), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n371_), .A2(new_n372_), .A3(new_n373_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND4_X1  g185(.A1(new_n386_), .A2(KEYINPUT95), .A3(new_n380_), .A4(new_n369_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n376_), .A2(new_n381_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n382_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT96), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT96), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n382_), .A2(new_n387_), .A3(new_n388_), .A4(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n347_), .B1(new_n390_), .B2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n363_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n350_), .B1(new_n394_), .B2(new_n368_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n353_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n396_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n397_), .A2(KEYINPUT32), .A3(new_n380_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n376_), .B1(KEYINPUT32), .B2(new_n380_), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n335_), .A2(new_n327_), .A3(new_n336_), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n400_), .B(KEYINPUT100), .Z(new_n401_));
  XNOR2_X1  g200(.A(new_n337_), .B(KEYINPUT99), .ZN(new_n402_));
  AOI211_X1 g201(.A(new_n398_), .B(new_n399_), .C1(new_n401_), .C2(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n322_), .B1(new_n393_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n402_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n271_), .A2(new_n321_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n272_), .A2(new_n320_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n405_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT27), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n389_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n397_), .A2(new_n381_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(KEYINPUT101), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n412_), .B(KEYINPUT27), .C1(new_n381_), .C2(new_n376_), .ZN(new_n413_));
  AND2_X1   g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n408_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n225_), .B1(new_n404_), .B2(new_n415_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT66), .B(KEYINPUT12), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT64), .ZN(new_n418_));
  OAI22_X1  g217(.A1(new_n418_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT7), .ZN(new_n420_));
  INV_X1    g219(.A(G99gat), .ZN(new_n421_));
  INV_X1    g220(.A(G106gat), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .A4(KEYINPUT64), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT6), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n424_), .B1(G99gat), .B2(G106gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G99gat), .A2(G106gat), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n426_), .A2(KEYINPUT6), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n419_), .B(new_n423_), .C1(new_n425_), .C2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G85gat), .ZN(new_n429_));
  INV_X1    g228(.A(G92gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G85gat), .A2(G92gat), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  AND3_X1   g232(.A1(new_n428_), .A2(KEYINPUT8), .A3(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT8), .B1(new_n428_), .B2(new_n433_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n426_), .A2(KEYINPUT6), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n424_), .A2(G99gat), .A3(G106gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OR2_X1    g237(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n439_));
  NAND2_X1  g238(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n422_), .A3(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n431_), .A2(KEYINPUT9), .A3(new_n432_), .ZN(new_n442_));
  OR2_X1    g241(.A1(new_n432_), .A2(KEYINPUT9), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n438_), .A2(new_n441_), .A3(new_n442_), .A4(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n434_), .A2(new_n435_), .A3(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G57gat), .B(G64gat), .ZN(new_n447_));
  INV_X1    g246(.A(G78gat), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(G71gat), .ZN(new_n449_));
  INV_X1    g248(.A(G71gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(G78gat), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n447_), .A2(KEYINPUT11), .A3(new_n449_), .A4(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G64gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G57gat), .ZN(new_n454_));
  INV_X1    g253(.A(G57gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(G64gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n456_), .A3(KEYINPUT11), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n449_), .A2(new_n451_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n447_), .A2(KEYINPUT11), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n452_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n417_), .B1(new_n446_), .B2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n428_), .A2(new_n433_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT8), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n428_), .A2(KEYINPUT8), .A3(new_n433_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(new_n466_), .A3(new_n444_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT65), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n468_), .B(new_n452_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n461_), .A2(KEYINPUT65), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n467_), .A2(KEYINPUT12), .A3(new_n469_), .A4(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G230gat), .A2(G233gat), .ZN(new_n472_));
  NAND4_X1  g271(.A1(new_n465_), .A2(new_n461_), .A3(new_n466_), .A4(new_n444_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n462_), .A2(new_n471_), .A3(new_n472_), .A4(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n472_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n446_), .A2(new_n461_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n473_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n474_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G120gat), .B(G148gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT5), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G176gat), .B(G204gat), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n481_), .B(new_n482_), .Z(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n479_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT67), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT13), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n485_), .A2(KEYINPUT67), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(KEYINPUT67), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n489_), .A2(KEYINPUT13), .A3(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G127gat), .B(G155gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT16), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G183gat), .B(G211gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(KEYINPUT17), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n497_), .B(KEYINPUT72), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G231gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n212_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(new_n461_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(KEYINPUT65), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT71), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n498_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n504_), .B1(new_n503_), .B2(new_n502_), .ZN(new_n505_));
  OR2_X1    g304(.A1(new_n496_), .A2(KEYINPUT17), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n501_), .A2(new_n497_), .A3(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(G190gat), .B(G218gat), .Z(new_n510_));
  XNOR2_X1  g309(.A(new_n510_), .B(KEYINPUT69), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G134gat), .B(G162gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT36), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT70), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n467_), .A2(new_n204_), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n516_), .B(KEYINPUT68), .Z(new_n517_));
  NAND2_X1  g316(.A1(G232gat), .A2(G233gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT34), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT35), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  AOI22_X1  g322(.A1(new_n205_), .A2(new_n467_), .B1(new_n521_), .B2(new_n520_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n517_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n523_), .B1(new_n517_), .B2(new_n524_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n515_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n527_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n513_), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n530_), .A2(KEYINPUT36), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n529_), .A2(new_n531_), .A3(new_n525_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(KEYINPUT37), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n514_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n532_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n534_), .B1(KEYINPUT37), .B2(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n492_), .A2(new_n509_), .A3(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(new_n538_), .B(KEYINPUT73), .Z(new_n539_));
  AND2_X1   g338(.A1(new_n416_), .A2(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(new_n207_), .A3(new_n405_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT38), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n541_), .A2(new_n542_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n536_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(new_n404_), .B2(new_n415_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n492_), .ZN(new_n547_));
  NOR3_X1   g346(.A1(new_n547_), .A2(new_n225_), .A3(new_n508_), .ZN(new_n548_));
  AND2_X1   g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n207_), .B1(new_n549_), .B2(new_n405_), .ZN(new_n550_));
  NOR3_X1   g349(.A1(new_n543_), .A2(new_n544_), .A3(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT102), .ZN(G1324gat));
  INV_X1    g351(.A(new_n414_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n540_), .A2(new_n208_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT103), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n549_), .A2(new_n553_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT39), .ZN(new_n557_));
  AND4_X1   g356(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .A4(G8gat), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n208_), .B1(KEYINPUT103), .B2(KEYINPUT39), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n556_), .A2(new_n559_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n554_), .B1(new_n558_), .B2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(new_n561_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g361(.A1(new_n549_), .A2(new_n272_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(G15gat), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT41), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(G15gat), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n540_), .A2(new_n567_), .A3(new_n272_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT104), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n569_), .B(new_n570_), .ZN(G1326gat));
  INV_X1    g370(.A(G22gat), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n572_), .B1(new_n549_), .B2(new_n321_), .ZN(new_n573_));
  XOR2_X1   g372(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n540_), .A2(new_n572_), .A3(new_n321_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(G1327gat));
  NOR3_X1   g376(.A1(new_n547_), .A2(new_n509_), .A3(new_n536_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n416_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(G29gat), .B1(new_n579_), .B2(new_n405_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n404_), .A2(new_n415_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n536_), .A2(KEYINPUT37), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n582_), .B1(KEYINPUT37), .B2(new_n533_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT43), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT43), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n581_), .A2(new_n586_), .A3(new_n583_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n225_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n492_), .A2(new_n589_), .A3(new_n508_), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT106), .Z(new_n591_));
  NAND4_X1  g390(.A1(new_n588_), .A2(KEYINPUT107), .A3(KEYINPUT44), .A4(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n586_), .B1(new_n581_), .B2(new_n583_), .ZN(new_n593_));
  AOI211_X1 g392(.A(KEYINPUT43), .B(new_n537_), .C1(new_n404_), .C2(new_n415_), .ZN(new_n594_));
  OAI211_X1 g393(.A(KEYINPUT44), .B(new_n591_), .C1(new_n593_), .C2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT107), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n588_), .A2(new_n591_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT44), .ZN(new_n599_));
  AOI22_X1  g398(.A1(new_n592_), .A2(new_n597_), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  AND2_X1   g399(.A1(new_n405_), .A2(G29gat), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n580_), .B1(new_n600_), .B2(new_n601_), .ZN(G1328gat));
  INV_X1    g401(.A(KEYINPUT46), .ZN(new_n603_));
  INV_X1    g402(.A(G36gat), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n600_), .B2(new_n553_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n579_), .A2(new_n604_), .A3(new_n553_), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n606_), .B(KEYINPUT45), .Z(new_n607_));
  OAI21_X1  g406(.A(new_n603_), .B1(new_n605_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n607_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n592_), .A2(new_n597_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n598_), .A2(new_n599_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n610_), .A2(new_n553_), .A3(new_n611_), .ZN(new_n612_));
  OAI211_X1 g411(.A(KEYINPUT46), .B(new_n609_), .C1(new_n612_), .C2(new_n604_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n608_), .A2(new_n613_), .ZN(G1329gat));
  NAND4_X1  g413(.A1(new_n610_), .A2(G43gat), .A3(new_n272_), .A4(new_n611_), .ZN(new_n615_));
  INV_X1    g414(.A(G43gat), .ZN(new_n616_));
  INV_X1    g415(.A(new_n579_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n616_), .B1(new_n617_), .B2(new_n271_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n615_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(KEYINPUT47), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT47), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n615_), .A2(new_n621_), .A3(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(G1330gat));
  AOI21_X1  g422(.A(G50gat), .B1(new_n579_), .B2(new_n321_), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n321_), .A2(G50gat), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n600_), .B2(new_n625_), .ZN(G1331gat));
  NOR3_X1   g425(.A1(new_n492_), .A2(new_n589_), .A3(new_n508_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n546_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n405_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G57gat), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n589_), .B1(new_n404_), .B2(new_n415_), .ZN(new_n632_));
  AND4_X1   g431(.A1(new_n547_), .A2(new_n632_), .A3(new_n509_), .A4(new_n537_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n633_), .A2(new_n455_), .A3(new_n405_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n634_), .ZN(G1332gat));
  NAND2_X1  g434(.A1(new_n553_), .A2(new_n453_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT108), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(G64gat), .B1(new_n629_), .B2(new_n414_), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n639_), .A2(KEYINPUT48), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(KEYINPUT48), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n638_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT109), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(G1333gat));
  AOI21_X1  g443(.A(new_n450_), .B1(new_n628_), .B2(new_n272_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT49), .Z(new_n646_));
  NAND3_X1  g445(.A1(new_n633_), .A2(new_n450_), .A3(new_n272_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1334gat));
  AOI21_X1  g447(.A(new_n448_), .B1(new_n628_), .B2(new_n321_), .ZN(new_n649_));
  XOR2_X1   g448(.A(new_n649_), .B(KEYINPUT50), .Z(new_n650_));
  NAND3_X1  g449(.A1(new_n633_), .A2(new_n448_), .A3(new_n321_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(G1335gat));
  NAND4_X1  g451(.A1(new_n632_), .A2(new_n547_), .A3(new_n508_), .A4(new_n545_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT110), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(new_n429_), .A3(new_n405_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n492_), .A2(new_n589_), .A3(new_n509_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n657_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n405_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n655_), .B1(new_n660_), .B2(new_n429_), .ZN(G1336gat));
  NAND3_X1  g460(.A1(new_n654_), .A2(new_n430_), .A3(new_n553_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n658_), .A2(new_n553_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n662_), .B1(new_n664_), .B2(new_n430_), .ZN(G1337gat));
  NAND4_X1  g464(.A1(new_n654_), .A2(new_n272_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n658_), .A2(new_n272_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(G99gat), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g469(.A1(new_n654_), .A2(new_n422_), .A3(new_n321_), .ZN(new_n671_));
  AOI211_X1 g470(.A(KEYINPUT52), .B(new_n422_), .C1(new_n658_), .C2(new_n321_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT52), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n658_), .A2(new_n321_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(G106gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n671_), .B1(new_n672_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT53), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT53), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n671_), .B(new_n678_), .C1(new_n672_), .C2(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1339gat));
  NOR2_X1   g479(.A1(new_n553_), .A2(new_n630_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n407_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(KEYINPUT59), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n474_), .A2(new_n478_), .A3(new_n484_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n589_), .A2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT56), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT111), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT55), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n474_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n474_), .B2(new_n689_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n470_), .A2(KEYINPUT12), .A3(new_n469_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n473_), .B1(new_n693_), .B2(new_n446_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n417_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n461_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n695_), .B1(new_n467_), .B2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n475_), .B1(new_n694_), .B2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n698_), .B1(new_n474_), .B2(new_n689_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT112), .B1(new_n692_), .B2(new_n699_), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n694_), .A2(new_n475_), .A3(new_n697_), .ZN(new_n701_));
  OAI21_X1  g500(.A(KEYINPUT111), .B1(new_n701_), .B2(KEYINPUT55), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n474_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT112), .ZN(new_n705_));
  INV_X1    g504(.A(new_n699_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n704_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  AOI211_X1 g506(.A(new_n687_), .B(new_n484_), .C1(new_n700_), .C2(new_n707_), .ZN(new_n708_));
  AOI211_X1 g507(.A(KEYINPUT112), .B(new_n699_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n705_), .B1(new_n704_), .B2(new_n706_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n483_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n687_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT113), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n708_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(KEYINPUT113), .A3(new_n687_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n686_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n213_), .A2(new_n214_), .A3(new_n218_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n222_), .B1(new_n217_), .B2(new_n215_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n223_), .B1(new_n717_), .B2(new_n718_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n486_), .A2(new_n719_), .ZN(new_n720_));
  OAI211_X1 g519(.A(KEYINPUT57), .B(new_n536_), .C1(new_n716_), .C2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT57), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n484_), .B1(new_n700_), .B2(new_n707_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n713_), .B1(new_n723_), .B2(KEYINPUT56), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(KEYINPUT56), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n724_), .A2(new_n715_), .A3(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n686_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n720_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n722_), .B1(new_n728_), .B2(new_n545_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT114), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(KEYINPUT58), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n719_), .A2(new_n685_), .ZN(new_n732_));
  AOI211_X1 g531(.A(new_n731_), .B(new_n732_), .C1(new_n712_), .C2(new_n725_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n712_), .B2(new_n725_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n731_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n583_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n721_), .B(new_n729_), .C1(new_n733_), .C2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(new_n508_), .ZN(new_n738_));
  NAND4_X1  g537(.A1(new_n492_), .A2(new_n225_), .A3(new_n509_), .A4(new_n537_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT54), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n739_), .B(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n738_), .A2(new_n742_), .ZN(new_n743_));
  AND2_X1   g542(.A1(new_n684_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(G113gat), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n225_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(KEYINPUT115), .B1(new_n736_), .B2(new_n733_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n723_), .A2(KEYINPUT56), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n749_), .A2(new_n708_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n731_), .B1(new_n750_), .B2(new_n732_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT115), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n734_), .A2(new_n735_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n751_), .A2(new_n752_), .A3(new_n753_), .A4(new_n583_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n721_), .A2(new_n729_), .A3(new_n748_), .A4(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(new_n508_), .ZN(new_n756_));
  AOI21_X1  g555(.A(KEYINPUT116), .B1(new_n756_), .B2(new_n742_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT116), .ZN(new_n758_));
  AOI211_X1 g557(.A(new_n758_), .B(new_n741_), .C1(new_n755_), .C2(new_n508_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n757_), .A2(new_n759_), .A3(new_n683_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT59), .ZN(new_n761_));
  OAI21_X1  g560(.A(KEYINPUT118), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n756_), .A2(new_n742_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(new_n758_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n756_), .A2(KEYINPUT116), .A3(new_n742_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n683_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n764_), .A2(new_n765_), .A3(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT118), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n768_), .A3(KEYINPUT59), .ZN(new_n769_));
  AOI211_X1 g568(.A(new_n744_), .B(new_n747_), .C1(new_n762_), .C2(new_n769_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n757_), .A2(new_n759_), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT117), .B1(new_n771_), .B2(new_n766_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT117), .ZN(new_n773_));
  NOR4_X1   g572(.A1(new_n757_), .A2(new_n759_), .A3(new_n773_), .A4(new_n683_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(G113gat), .B1(new_n775_), .B2(new_n589_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT119), .B1(new_n770_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n762_), .A2(new_n769_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n744_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n778_), .A2(new_n779_), .A3(new_n746_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT119), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n760_), .A2(KEYINPUT117), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n767_), .A2(new_n773_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n745_), .B1(new_n784_), .B2(new_n225_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n780_), .A2(new_n781_), .A3(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n777_), .A2(new_n786_), .ZN(G1340gat));
  INV_X1    g586(.A(G120gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n492_), .B2(KEYINPUT60), .ZN(new_n789_));
  OAI211_X1 g588(.A(new_n775_), .B(new_n789_), .C1(KEYINPUT60), .C2(new_n788_), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n492_), .B(new_n744_), .C1(new_n762_), .C2(new_n769_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(new_n788_), .ZN(G1341gat));
  INV_X1    g591(.A(G127gat), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n775_), .A2(new_n793_), .A3(new_n509_), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n508_), .B(new_n744_), .C1(new_n762_), .C2(new_n769_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n794_), .B1(new_n795_), .B2(new_n793_), .ZN(G1342gat));
  INV_X1    g595(.A(G134gat), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n775_), .A2(new_n797_), .A3(new_n545_), .ZN(new_n798_));
  AOI211_X1 g597(.A(new_n537_), .B(new_n744_), .C1(new_n762_), .C2(new_n769_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n797_), .ZN(G1343gat));
  NAND2_X1  g599(.A1(new_n764_), .A2(new_n765_), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n553_), .A2(new_n630_), .A3(new_n406_), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n802_), .B(KEYINPUT120), .Z(new_n803_));
  NOR2_X1   g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n589_), .ZN(new_n805_));
  XNOR2_X1  g604(.A(new_n805_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n547_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g607(.A1(new_n804_), .A2(new_n509_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT121), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT121), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n804_), .A2(new_n811_), .A3(new_n509_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(KEYINPUT61), .B(G155gat), .ZN(new_n813_));
  AND3_X1   g612(.A1(new_n810_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n813_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n814_), .A2(new_n815_), .ZN(G1346gat));
  AOI21_X1  g615(.A(G162gat), .B1(new_n804_), .B2(new_n545_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n583_), .A2(G162gat), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(KEYINPUT122), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n817_), .B1(new_n804_), .B2(new_n819_), .ZN(G1347gat));
  NAND2_X1  g619(.A1(new_n553_), .A2(new_n630_), .ZN(new_n821_));
  NOR3_X1   g620(.A1(new_n821_), .A2(new_n271_), .A3(new_n225_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n321_), .B1(new_n822_), .B2(KEYINPUT123), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(KEYINPUT123), .B2(new_n822_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n743_), .ZN(new_n825_));
  OAI21_X1  g624(.A(G169gat), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(KEYINPUT62), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n821_), .A2(new_n407_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n743_), .A2(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n589_), .A2(new_n234_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n827_), .B1(new_n829_), .B2(new_n830_), .ZN(G1348gat));
  NOR2_X1   g630(.A1(new_n801_), .A2(new_n321_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n821_), .A2(new_n271_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n832_), .A2(G176gat), .A3(new_n547_), .A4(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n235_), .B1(new_n829_), .B2(new_n492_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n834_), .A2(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(KEYINPUT124), .ZN(G1349gat));
  NOR3_X1   g636(.A1(new_n829_), .A2(new_n251_), .A3(new_n508_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n832_), .A2(new_n509_), .A3(new_n833_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n838_), .B1(new_n839_), .B2(new_n241_), .ZN(G1350gat));
  OAI21_X1  g639(.A(G190gat), .B1(new_n829_), .B2(new_n537_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n545_), .A2(new_n252_), .ZN(new_n842_));
  XOR2_X1   g641(.A(new_n842_), .B(KEYINPUT125), .Z(new_n843_));
  OAI21_X1  g642(.A(new_n841_), .B1(new_n829_), .B2(new_n843_), .ZN(G1351gat));
  NOR3_X1   g643(.A1(new_n801_), .A2(new_n406_), .A3(new_n821_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n589_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT126), .B(G197gat), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n846_), .B2(new_n849_), .ZN(G1352gat));
  NAND2_X1  g649(.A1(new_n845_), .A2(new_n547_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g651(.A1(new_n845_), .A2(new_n509_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n854_));
  AND2_X1   g653(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n853_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n853_), .B2(new_n854_), .ZN(G1354gat));
  NAND2_X1  g656(.A1(new_n845_), .A2(new_n545_), .ZN(new_n858_));
  XOR2_X1   g657(.A(KEYINPUT127), .B(G218gat), .Z(new_n859_));
  NOR2_X1   g658(.A1(new_n537_), .A2(new_n859_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n858_), .A2(new_n859_), .B1(new_n845_), .B2(new_n860_), .ZN(G1355gat));
endmodule


