//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 0 0 1 0 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:24 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n758_, new_n759_, new_n760_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n939_, new_n941_, new_n942_, new_n943_,
    new_n945_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n953_, new_n954_, new_n955_, new_n956_;
  AND3_X1   g000(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n202_));
  AOI21_X1  g001(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n203_));
  NOR2_X1   g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT10), .B(G99gat), .ZN(new_n205_));
  AOI21_X1  g004(.A(KEYINPUT64), .B1(G85gat), .B2(G92gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT9), .ZN(new_n207_));
  OAI22_X1  g006(.A1(new_n206_), .A2(new_n207_), .B1(G85gat), .B2(G92gat), .ZN(new_n208_));
  AND2_X1   g007(.A1(new_n206_), .A2(new_n207_), .ZN(new_n209_));
  OAI221_X1 g008(.A(new_n204_), .B1(G106gat), .B2(new_n205_), .C1(new_n208_), .C2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT8), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NOR3_X1   g012(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT6), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT65), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT65), .B1(new_n202_), .B2(new_n203_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n215_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  XOR2_X1   g022(.A(G85gat), .B(G92gat), .Z(new_n224_));
  AOI21_X1  g023(.A(new_n211_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n211_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n226_), .B1(new_n204_), .B2(new_n215_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n210_), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT66), .B(KEYINPUT67), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(G50gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G43gat), .ZN(new_n232_));
  INV_X1    g031(.A(G43gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(G50gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n232_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G29gat), .B(G36gat), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(G36gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(G29gat), .ZN(new_n239_));
  INV_X1    g038(.A(G29gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(G36gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n230_), .B1(new_n237_), .B2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n243_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n235_), .A2(new_n236_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n246_), .A2(new_n247_), .A3(new_n229_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n245_), .A2(new_n248_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n228_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G232gat), .A2(G233gat), .ZN(new_n251_));
  XOR2_X1   g050(.A(new_n251_), .B(KEYINPUT34), .Z(new_n252_));
  INV_X1    g051(.A(KEYINPUT35), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT70), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n256_), .B1(new_n253_), .B2(new_n252_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT15), .ZN(new_n258_));
  AND3_X1   g057(.A1(new_n246_), .A2(new_n247_), .A3(new_n229_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n229_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n258_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n245_), .A2(KEYINPUT15), .A3(new_n248_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  AND3_X1   g062(.A1(new_n263_), .A2(KEYINPUT68), .A3(new_n228_), .ZN(new_n264_));
  AOI21_X1  g063(.A(KEYINPUT68), .B1(new_n263_), .B2(new_n228_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n257_), .A2(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT69), .B1(new_n264_), .B2(new_n265_), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n259_), .A2(new_n260_), .A3(new_n258_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT15), .B1(new_n245_), .B2(new_n248_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n228_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n263_), .A2(KEYINPUT68), .A3(new_n228_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n268_), .A2(new_n276_), .A3(new_n256_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n252_), .A2(new_n253_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n277_), .A2(KEYINPUT71), .A3(new_n278_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n267_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G190gat), .B(G218gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G134gat), .B(G162gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(new_n286_), .B(KEYINPUT36), .Z(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n283_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n286_), .A2(KEYINPUT36), .ZN(new_n290_));
  INV_X1    g089(.A(new_n267_), .ZN(new_n291_));
  AND3_X1   g090(.A1(new_n277_), .A2(KEYINPUT71), .A3(new_n278_), .ZN(new_n292_));
  AOI21_X1  g091(.A(KEYINPUT71), .B1(new_n277_), .B2(new_n278_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n290_), .B(new_n291_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT37), .ZN(new_n295_));
  OR2_X1    g094(.A1(new_n289_), .A2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n288_), .B1(new_n297_), .B2(KEYINPUT72), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n299_), .B(new_n291_), .C1(new_n292_), .C2(new_n293_), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n298_), .A2(new_n300_), .B1(new_n290_), .B2(new_n283_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n296_), .B1(new_n301_), .B2(KEYINPUT37), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G127gat), .B(G155gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G183gat), .B(G211gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G71gat), .B(G78gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(G57gat), .B(G64gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n308_), .B1(KEYINPUT11), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(KEYINPUT11), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G15gat), .B(G22gat), .ZN(new_n314_));
  INV_X1    g113(.A(G1gat), .ZN(new_n315_));
  INV_X1    g114(.A(G8gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT14), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n314_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G1gat), .B(G8gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT73), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(KEYINPUT73), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G231gat), .A2(G233gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n325_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n313_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n328_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(new_n326_), .A3(new_n312_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n307_), .B1(new_n332_), .B2(KEYINPUT17), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT75), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n329_), .A2(new_n331_), .A3(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n307_), .A2(KEYINPUT17), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n333_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n335_), .B1(new_n333_), .B2(new_n336_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n302_), .A2(new_n340_), .ZN(new_n341_));
  OR2_X1    g140(.A1(new_n341_), .A2(KEYINPUT76), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(KEYINPUT76), .ZN(new_n343_));
  AND2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G127gat), .B(G134gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT87), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT88), .ZN(new_n348_));
  XOR2_X1   g147(.A(G113gat), .B(G120gat), .Z(new_n349_));
  NAND3_X1  g148(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n347_), .B(new_n349_), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n350_), .B1(new_n351_), .B2(new_n348_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G155gat), .A2(G162gat), .ZN(new_n353_));
  XOR2_X1   g152(.A(new_n353_), .B(KEYINPUT1), .Z(new_n354_));
  NOR2_X1   g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT90), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G141gat), .ZN(new_n358_));
  INV_X1    g157(.A(G148gat), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n359_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n357_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT2), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n364_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n366_));
  OAI211_X1 g165(.A(new_n365_), .B(new_n366_), .C1(KEYINPUT3), .C2(new_n362_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n362_), .A2(KEYINPUT3), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT91), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT91), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n362_), .A2(new_n370_), .A3(KEYINPUT3), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n367_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n356_), .A2(new_n353_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n363_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n352_), .A2(new_n374_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n351_), .B(new_n363_), .C1(new_n372_), .C2(new_n373_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n375_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G225gat), .A2(G233gat), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n375_), .A2(KEYINPUT4), .A3(new_n376_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(KEYINPUT100), .B(KEYINPUT4), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n352_), .A2(new_n374_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n378_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G1gat), .B(G29gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT0), .ZN(new_n386_));
  INV_X1    g185(.A(G57gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n386_), .B(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(G85gat), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n380_), .A2(new_n384_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n393_), .A2(KEYINPUT103), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n391_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT103), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n395_), .B1(new_n392_), .B2(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n394_), .A2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT104), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G226gat), .A2(G233gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT19), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT96), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G211gat), .B(G218gat), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT95), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G197gat), .A2(G204gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT93), .B(G197gat), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n407_), .B1(new_n408_), .B2(G204gat), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT21), .ZN(new_n411_));
  NOR3_X1   g210(.A1(new_n406_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G204gat), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(G197gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n408_), .A2(new_n413_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n414_), .B1(new_n415_), .B2(KEYINPUT94), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT94), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n408_), .A2(new_n417_), .A3(new_n413_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT21), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n404_), .B(KEYINPUT95), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(new_n411_), .B2(new_n410_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n412_), .B1(new_n420_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G183gat), .A2(G190gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT23), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT24), .ZN(new_n426_));
  INV_X1    g225(.A(G169gat), .ZN(new_n427_));
  INV_X1    g226(.A(G176gat), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT25), .B(G183gat), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT79), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(G190gat), .ZN(new_n434_));
  OR3_X1    g233(.A1(new_n434_), .A2(KEYINPUT80), .A3(KEYINPUT26), .ZN(new_n435_));
  INV_X1    g234(.A(G183gat), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n432_), .B1(new_n436_), .B2(KEYINPUT25), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT26), .B1(new_n434_), .B2(KEYINPUT80), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n435_), .A2(new_n437_), .A3(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G169gat), .A2(G176gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT81), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT82), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n441_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT81), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n440_), .B(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n443_), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT82), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  OAI221_X1 g247(.A(new_n430_), .B1(new_n433_), .B2(new_n439_), .C1(new_n444_), .C2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(KEYINPUT83), .B(G176gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT22), .B(G169gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n446_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT84), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n446_), .A3(KEYINPUT84), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n425_), .B1(G183gat), .B2(G190gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n423_), .A2(new_n449_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT20), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n421_), .A2(KEYINPUT21), .A3(new_n409_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n411_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n406_), .B1(KEYINPUT21), .B2(new_n409_), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n461_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT26), .B(G190gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n431_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT97), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n447_), .A2(new_n440_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n467_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n430_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n451_), .B(KEYINPUT98), .ZN(new_n472_));
  INV_X1    g271(.A(new_n450_), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n446_), .B(new_n457_), .C1(new_n472_), .C2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(new_n474_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n460_), .B1(new_n464_), .B2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n403_), .B1(new_n459_), .B2(new_n476_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n401_), .A2(new_n460_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n478_), .B1(new_n464_), .B2(new_n475_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n420_), .A2(new_n422_), .ZN(new_n480_));
  AOI22_X1  g279(.A1(new_n480_), .A2(new_n461_), .B1(new_n449_), .B2(new_n458_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G8gat), .B(G36gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT18), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(G64gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(G92gat), .ZN(new_n486_));
  NOR3_X1   g285(.A1(new_n477_), .A2(new_n482_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT99), .ZN(new_n488_));
  OAI21_X1  g287(.A(new_n486_), .B1(new_n477_), .B2(new_n482_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  OAI211_X1 g289(.A(KEYINPUT99), .B(new_n486_), .C1(new_n477_), .C2(new_n482_), .ZN(new_n491_));
  AOI21_X1  g290(.A(KEYINPUT27), .B1(new_n490_), .B2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT27), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n487_), .A2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT102), .B(KEYINPUT20), .Z(new_n495_));
  OAI21_X1  g294(.A(new_n495_), .B1(new_n464_), .B2(new_n475_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n401_), .B1(new_n496_), .B2(new_n481_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n459_), .A2(new_n476_), .A3(new_n403_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n486_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n494_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n399_), .B1(new_n492_), .B2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n487_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n489_), .A2(new_n488_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n505_), .A3(new_n491_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n493_), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(KEYINPUT104), .A3(new_n501_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G22gat), .B(G50gat), .ZN(new_n509_));
  XOR2_X1   g308(.A(new_n509_), .B(KEYINPUT28), .Z(new_n510_));
  NAND2_X1  g309(.A1(new_n374_), .A2(KEYINPUT29), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G78gat), .B(G106gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n464_), .A3(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n512_), .B1(new_n511_), .B2(new_n464_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n510_), .B1(new_n514_), .B2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n515_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n510_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n513_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n516_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G228gat), .A2(G233gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n521_), .B1(new_n423_), .B2(KEYINPUT92), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n374_), .A2(KEYINPUT29), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n523_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n520_), .A2(new_n526_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n516_), .A2(new_n519_), .A3(new_n524_), .A4(new_n525_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT31), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n352_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT89), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G227gat), .A2(G233gat), .ZN(new_n534_));
  XNOR2_X1  g333(.A(new_n534_), .B(KEYINPUT86), .ZN(new_n535_));
  XOR2_X1   g334(.A(G71gat), .B(G99gat), .Z(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT85), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n449_), .A2(new_n539_), .A3(new_n458_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n539_), .B1(new_n449_), .B2(new_n458_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G15gat), .B(G43gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT30), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n542_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n540_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n545_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n538_), .B1(new_n546_), .B2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n546_), .A2(new_n550_), .A3(new_n538_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n533_), .A2(new_n552_), .A3(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n553_), .ZN(new_n555_));
  OAI22_X1  g354(.A1(new_n555_), .A2(new_n551_), .B1(new_n532_), .B2(new_n531_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n529_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n503_), .A2(new_n508_), .A3(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n554_), .A2(new_n556_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n560_), .A2(new_n529_), .A3(new_n507_), .A4(new_n501_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n398_), .B1(new_n558_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n529_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n560_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n506_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n390_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n566_));
  AND2_X1   g365(.A1(new_n381_), .A2(new_n383_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n567_), .B2(new_n378_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT33), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n395_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n395_), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT101), .B1(new_n571_), .B2(KEYINPUT33), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT101), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n395_), .A2(new_n573_), .A3(new_n569_), .ZN(new_n574_));
  OAI211_X1 g373(.A(new_n565_), .B(new_n570_), .C1(new_n572_), .C2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT32), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n486_), .A2(new_n576_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n577_), .A2(new_n477_), .A3(new_n482_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n578_), .B1(new_n499_), .B2(new_n577_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n579_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n564_), .B1(new_n575_), .B2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n562_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G230gat), .A2(G233gat), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  OR2_X1    g383(.A1(new_n228_), .A2(new_n312_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n228_), .A2(new_n312_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n585_), .A2(KEYINPUT12), .A3(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT12), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n228_), .A2(new_n588_), .A3(new_n312_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n584_), .B1(new_n587_), .B2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n583_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(G120gat), .B(G148gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(new_n413_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT5), .B(G176gat), .ZN(new_n595_));
  XOR2_X1   g394(.A(new_n594_), .B(new_n595_), .Z(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  OR3_X1    g396(.A1(new_n591_), .A2(new_n592_), .A3(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n597_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT13), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n598_), .A2(KEYINPUT13), .A3(new_n599_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n263_), .A2(new_n320_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n321_), .A2(new_n248_), .A3(new_n245_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(G229gat), .A2(G233gat), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n605_), .A2(new_n606_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT77), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n249_), .A2(new_n320_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n606_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n607_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n609_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  AOI211_X1 g412(.A(KEYINPUT77), .B(new_n607_), .C1(new_n606_), .C2(new_n610_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n608_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G113gat), .B(G141gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(G197gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(KEYINPUT78), .B(G169gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n617_), .B(new_n618_), .Z(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n608_), .B(new_n621_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n604_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n582_), .A2(new_n626_), .ZN(new_n627_));
  AND2_X1   g426(.A1(new_n344_), .A2(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n315_), .A3(new_n398_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT38), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(KEYINPUT106), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT106), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n631_), .B1(new_n632_), .B2(KEYINPUT38), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n629_), .A2(KEYINPUT106), .A3(new_n630_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT105), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n635_), .B1(new_n582_), .B2(new_n301_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n287_), .B1(new_n283_), .B2(new_n299_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n300_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n294_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  OAI211_X1 g438(.A(KEYINPUT105), .B(new_n639_), .C1(new_n562_), .C2(new_n581_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n625_), .A2(new_n339_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n394_), .A2(new_n397_), .ZN(new_n645_));
  OAI21_X1  g444(.A(G1gat), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n633_), .A2(new_n634_), .A3(new_n646_), .ZN(G1324gat));
  XNOR2_X1  g446(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT108), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n503_), .A2(new_n508_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  AOI211_X1 g451(.A(new_n652_), .B(new_n642_), .C1(new_n636_), .C2(new_n640_), .ZN(new_n653_));
  OAI21_X1  g452(.A(KEYINPUT39), .B1(new_n653_), .B2(new_n316_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n641_), .A2(new_n651_), .A3(new_n643_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(G8gat), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n652_), .A2(G8gat), .ZN(new_n659_));
  AND4_X1   g458(.A1(new_n342_), .A2(new_n343_), .A3(new_n627_), .A4(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n650_), .B1(new_n658_), .B2(new_n661_), .ZN(new_n662_));
  AOI211_X1 g461(.A(KEYINPUT108), .B(new_n660_), .C1(new_n654_), .C2(new_n657_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n649_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n653_), .A2(KEYINPUT39), .A3(new_n316_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n656_), .B1(new_n655_), .B2(G8gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n661_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT108), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n658_), .A2(new_n650_), .A3(new_n661_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n648_), .A3(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n664_), .A2(new_n670_), .ZN(G1325gat));
  OAI21_X1  g470(.A(G15gat), .B1(new_n644_), .B2(new_n560_), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT41), .Z(new_n673_));
  INV_X1    g472(.A(G15gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n628_), .A2(new_n674_), .A3(new_n559_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(G1326gat));
  OAI21_X1  g475(.A(G22gat), .B1(new_n644_), .B2(new_n563_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT42), .ZN(new_n678_));
  INV_X1    g477(.A(G22gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n628_), .A2(new_n679_), .A3(new_n529_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1327gat));
  INV_X1    g480(.A(KEYINPUT109), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n289_), .A2(new_n295_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT37), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n639_), .B2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n682_), .B1(new_n582_), .B2(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n686_), .A2(KEYINPUT43), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n682_), .B(new_n688_), .C1(new_n582_), .C2(new_n685_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n626_), .A2(new_n339_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(KEYINPUT44), .A3(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n687_), .A2(new_n689_), .A3(new_n691_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  AND3_X1   g494(.A1(new_n692_), .A2(new_n398_), .A3(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n582_), .A2(new_n639_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(new_n691_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n645_), .A2(G29gat), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT110), .ZN(new_n700_));
  OAI22_X1  g499(.A1(new_n696_), .A2(new_n240_), .B1(new_n698_), .B2(new_n700_), .ZN(G1328gat));
  NAND2_X1  g500(.A1(new_n695_), .A2(new_n651_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n693_), .A2(new_n694_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G36gat), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n698_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n705_), .A2(new_n238_), .A3(new_n651_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT45), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n704_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT46), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n704_), .A2(new_n707_), .A3(KEYINPUT46), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(G1329gat));
  OAI21_X1  g511(.A(new_n233_), .B1(new_n698_), .B2(new_n560_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT111), .Z(new_n714_));
  NAND4_X1  g513(.A1(new_n692_), .A2(G43gat), .A3(new_n559_), .A4(new_n695_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(KEYINPUT47), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n714_), .A2(new_n715_), .A3(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n717_), .A2(new_n719_), .ZN(G1330gat));
  AOI21_X1  g519(.A(G50gat), .B1(new_n705_), .B2(new_n529_), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n231_), .B(new_n563_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(new_n692_), .ZN(G1331gat));
  INV_X1    g522(.A(new_n604_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(new_n623_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n582_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n344_), .A2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(new_n387_), .A3(new_n398_), .ZN(new_n730_));
  AOI211_X1 g529(.A(new_n340_), .B(new_n726_), .C1(new_n636_), .C2(new_n640_), .ZN(new_n731_));
  AND2_X1   g530(.A1(new_n731_), .A2(new_n398_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n730_), .B1(new_n732_), .B2(new_n387_), .ZN(G1332gat));
  INV_X1    g532(.A(G64gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n731_), .B2(new_n651_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT48), .Z(new_n736_));
  NAND2_X1  g535(.A1(new_n651_), .A2(new_n734_), .ZN(new_n737_));
  XOR2_X1   g536(.A(new_n737_), .B(KEYINPUT112), .Z(new_n738_));
  OAI21_X1  g537(.A(new_n736_), .B1(new_n728_), .B2(new_n738_), .ZN(G1333gat));
  INV_X1    g538(.A(G71gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(new_n731_), .B2(new_n559_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT49), .Z(new_n742_));
  NAND3_X1  g541(.A1(new_n729_), .A2(new_n740_), .A3(new_n559_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(G1334gat));
  INV_X1    g543(.A(G78gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n731_), .B2(new_n529_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT50), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n729_), .A2(new_n745_), .A3(new_n529_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1335gat));
  NAND2_X1  g548(.A1(new_n725_), .A2(new_n340_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT114), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n690_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n645_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n697_), .A2(new_n340_), .A3(new_n725_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT113), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n389_), .A3(new_n398_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n756_), .ZN(G1336gat));
  OAI21_X1  g556(.A(G92gat), .B1(new_n752_), .B2(new_n652_), .ZN(new_n758_));
  INV_X1    g557(.A(G92gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n755_), .A2(new_n759_), .A3(new_n651_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(G1337gat));
  OAI21_X1  g560(.A(G99gat), .B1(new_n752_), .B2(new_n560_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n205_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n755_), .A2(new_n763_), .A3(new_n559_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g565(.A1(new_n687_), .A2(new_n751_), .A3(new_n529_), .A4(new_n689_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(G106gat), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT115), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771_));
  AOI21_X1  g570(.A(KEYINPUT115), .B1(new_n767_), .B2(G106gat), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n770_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n563_), .A2(G106gat), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n755_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n768_), .A2(new_n769_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(KEYINPUT52), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT53), .B1(new_n773_), .B2(new_n777_), .ZN(new_n778_));
  AOI22_X1  g577(.A1(new_n772_), .A2(new_n771_), .B1(new_n755_), .B2(new_n774_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT53), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n776_), .A2(KEYINPUT52), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n779_), .B(new_n780_), .C1(new_n781_), .C2(new_n770_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n778_), .A2(new_n782_), .ZN(G1339gat));
  INV_X1    g582(.A(KEYINPUT56), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n591_), .A2(new_n785_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n228_), .A2(new_n312_), .ZN(new_n787_));
  OAI21_X1  g586(.A(KEYINPUT12), .B1(new_n228_), .B2(new_n312_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n583_), .B1(new_n789_), .B2(new_n589_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT55), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n789_), .A2(new_n589_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n786_), .A2(new_n791_), .B1(new_n584_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n784_), .B1(new_n793_), .B2(new_n596_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n584_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n591_), .A2(new_n785_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n790_), .A2(KEYINPUT55), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n798_), .A2(KEYINPUT56), .A3(new_n597_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n794_), .A2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n622_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n621_), .B1(new_n611_), .B2(new_n607_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n605_), .A2(new_n606_), .A3(new_n612_), .ZN(new_n803_));
  AND2_X1   g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n801_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n598_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(KEYINPUT58), .B1(new_n800_), .B2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT58), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n809_), .B(new_n806_), .C1(new_n794_), .C2(new_n799_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n600_), .A2(new_n805_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n784_), .A2(KEYINPUT117), .ZN(new_n813_));
  INV_X1    g612(.A(new_n813_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n798_), .A2(new_n597_), .A3(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(new_n598_), .A3(new_n623_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n813_), .B1(new_n793_), .B2(new_n596_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n812_), .B1(new_n816_), .B2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n639_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n302_), .A2(new_n811_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n820_), .A2(new_n821_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n822_), .A2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826_));
  NAND4_X1  g625(.A1(new_n724_), .A2(new_n826_), .A3(new_n339_), .A4(new_n624_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n339_), .A2(new_n624_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT116), .B1(new_n828_), .B2(new_n604_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n685_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT54), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT54), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n685_), .A2(new_n830_), .A3(new_n833_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n825_), .A2(new_n340_), .B1(new_n832_), .B2(new_n834_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n835_), .A2(new_n558_), .A3(new_n645_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT59), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n823_), .B1(new_n822_), .B2(KEYINPUT118), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n302_), .A2(new_n811_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n598_), .A2(new_n623_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n786_), .A2(new_n791_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n596_), .B1(new_n841_), .B2(new_n795_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n840_), .B1(new_n842_), .B2(new_n814_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n843_), .A2(new_n817_), .B1(new_n600_), .B2(new_n805_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n821_), .B1(new_n301_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n839_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT118), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n339_), .B1(new_n838_), .B2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n832_), .A2(new_n834_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n652_), .A2(new_n837_), .A3(new_n557_), .A4(new_n398_), .ZN(new_n853_));
  OAI22_X1  g652(.A1(new_n836_), .A2(new_n837_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  OAI21_X1  g653(.A(G113gat), .B1(new_n854_), .B2(new_n624_), .ZN(new_n855_));
  INV_X1    g654(.A(G113gat), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n836_), .A2(new_n856_), .A3(new_n623_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(G1340gat));
  NOR2_X1   g657(.A1(new_n724_), .A2(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n836_), .B1(KEYINPUT60), .B2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n604_), .ZN(new_n861_));
  OAI21_X1  g660(.A(G120gat), .B1(new_n861_), .B2(new_n854_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n862_), .B1(KEYINPUT60), .B2(new_n860_), .ZN(G1341gat));
  OAI21_X1  g662(.A(G127gat), .B1(new_n854_), .B2(new_n340_), .ZN(new_n864_));
  INV_X1    g663(.A(G127gat), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n836_), .A2(new_n865_), .A3(new_n339_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1342gat));
  XNOR2_X1  g666(.A(KEYINPUT120), .B(G134gat), .ZN(new_n868_));
  NOR3_X1   g667(.A1(new_n854_), .A2(new_n685_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(G134gat), .B1(new_n836_), .B2(new_n301_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n870_), .A2(KEYINPUT119), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(KEYINPUT119), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n869_), .A2(new_n871_), .A3(new_n872_), .ZN(G1343gat));
  NAND4_X1  g672(.A1(new_n652_), .A2(new_n560_), .A3(new_n529_), .A4(new_n398_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(KEYINPUT121), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n835_), .A2(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n623_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT122), .B(G141gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1344gat));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n604_), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n880_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g680(.A(KEYINPUT123), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n876_), .B2(new_n339_), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n835_), .A2(KEYINPUT123), .A3(new_n340_), .A4(new_n875_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT61), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n825_), .A2(new_n340_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n886_), .A2(new_n850_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n875_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(KEYINPUT123), .B1(new_n889_), .B2(new_n340_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT61), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n876_), .A2(new_n882_), .A3(new_n339_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n890_), .A2(new_n891_), .A3(new_n892_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n885_), .A2(new_n893_), .A3(G155gat), .ZN(new_n894_));
  AOI21_X1  g693(.A(G155gat), .B1(new_n885_), .B2(new_n893_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1346gat));
  OR3_X1    g695(.A1(new_n889_), .A2(G162gat), .A3(new_n639_), .ZN(new_n897_));
  OAI21_X1  g696(.A(G162gat), .B1(new_n889_), .B2(new_n685_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1347gat));
  NAND3_X1  g698(.A1(new_n651_), .A2(new_n559_), .A3(new_n645_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n900_), .A2(KEYINPUT124), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n900_), .A2(KEYINPUT124), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n563_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n793_), .A2(new_n784_), .A3(new_n596_), .ZN(new_n906_));
  AOI21_X1  g705(.A(KEYINPUT56), .B1(new_n798_), .B2(new_n597_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n807_), .B1(new_n906_), .B2(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n809_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n800_), .A2(KEYINPUT58), .A3(new_n807_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  OAI211_X1 g710(.A(KEYINPUT118), .B(new_n845_), .C1(new_n685_), .C2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n824_), .ZN(new_n913_));
  AOI21_X1  g712(.A(KEYINPUT118), .B1(new_n839_), .B2(new_n845_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n340_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n905_), .B1(new_n915_), .B2(new_n850_), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n427_), .B1(new_n916_), .B2(new_n623_), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n917_), .A2(KEYINPUT62), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(KEYINPUT62), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n916_), .A2(new_n623_), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n918_), .B(new_n919_), .C1(new_n472_), .C2(new_n920_), .ZN(G1348gat));
  NOR3_X1   g720(.A1(new_n903_), .A2(new_n428_), .A3(new_n724_), .ZN(new_n922_));
  NAND3_X1  g721(.A1(new_n887_), .A2(new_n563_), .A3(new_n922_), .ZN(new_n923_));
  INV_X1    g722(.A(KEYINPUT125), .ZN(new_n924_));
  AOI211_X1 g723(.A(new_n924_), .B(new_n473_), .C1(new_n916_), .C2(new_n604_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n903_), .A2(new_n529_), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n604_), .B(new_n926_), .C1(new_n849_), .C2(new_n851_), .ZN(new_n927_));
  AOI21_X1  g726(.A(KEYINPUT125), .B1(new_n927_), .B2(new_n450_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n923_), .B1(new_n925_), .B2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(KEYINPUT126), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT126), .ZN(new_n931_));
  OAI211_X1 g730(.A(new_n931_), .B(new_n923_), .C1(new_n925_), .C2(new_n928_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n930_), .A2(new_n932_), .ZN(G1349gat));
  OAI21_X1  g732(.A(new_n926_), .B1(new_n849_), .B2(new_n851_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n934_), .A2(new_n340_), .A3(new_n431_), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n887_), .A2(new_n339_), .A3(new_n563_), .A4(new_n904_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n935_), .B1(new_n436_), .B2(new_n936_), .ZN(G1350gat));
  OAI21_X1  g736(.A(G190gat), .B1(new_n934_), .B2(new_n685_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n916_), .A2(new_n301_), .A3(new_n465_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1351gat));
  NOR4_X1   g739(.A1(new_n652_), .A2(new_n559_), .A3(new_n398_), .A4(new_n563_), .ZN(new_n941_));
  AND2_X1   g740(.A1(new_n887_), .A2(new_n941_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n942_), .A2(new_n623_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g743(.A1(new_n887_), .A2(new_n941_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n724_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(new_n413_), .ZN(G1353gat));
  NAND2_X1  g746(.A1(new_n942_), .A2(new_n339_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n949_));
  AND2_X1   g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n948_), .A2(new_n949_), .A3(new_n950_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n951_), .B1(new_n948_), .B2(new_n949_), .ZN(G1354gat));
  INV_X1    g751(.A(G218gat), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n942_), .A2(new_n953_), .A3(new_n301_), .ZN(new_n954_));
  OAI21_X1  g753(.A(G218gat), .B1(new_n945_), .B2(new_n685_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n954_), .A2(new_n955_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


