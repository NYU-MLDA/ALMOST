//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n794_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n923_, new_n924_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n940_,
    new_n941_, new_n942_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n951_, new_n952_, new_n953_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n960_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  XOR2_X1   g001(.A(G113gat), .B(G120gat), .Z(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  OAI21_X1  g003(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT88), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR2_X1   g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n210_));
  AOI22_X1  g009(.A1(new_n208_), .A2(KEYINPUT2), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT85), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n207_), .B(new_n212_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n206_), .B(new_n211_), .C1(KEYINPUT2), .C2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G155gat), .ZN(new_n215_));
  INV_X1    g014(.A(G162gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(KEYINPUT86), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT86), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(G155gat), .B2(G162gat), .ZN(new_n219_));
  AOI22_X1  g018(.A1(new_n217_), .A2(new_n219_), .B1(G155gat), .B2(G162gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n214_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n213_), .A2(new_n209_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G155gat), .A2(G162gat), .ZN(new_n225_));
  AOI22_X1  g024(.A1(new_n217_), .A2(new_n219_), .B1(KEYINPUT1), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT87), .ZN(new_n227_));
  OR2_X1    g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(new_n225_), .A2(KEYINPUT1), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n229_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n224_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n204_), .B1(new_n222_), .B2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n228_), .A2(new_n230_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(new_n223_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n204_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(new_n221_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n232_), .A2(KEYINPUT4), .A3(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G225gat), .A2(G233gat), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n234_), .A2(new_n221_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(new_n241_), .A3(new_n204_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n237_), .A2(new_n239_), .A3(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n232_), .A2(new_n236_), .A3(new_n238_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G1gat), .B(G29gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n246_), .B(G85gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT0), .B(G57gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n247_), .B(new_n248_), .Z(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n245_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n243_), .A2(new_n244_), .A3(new_n249_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NOR2_X1   g053(.A1(new_n254_), .A2(G1gat), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT97), .ZN(new_n256_));
  XNOR2_X1  g055(.A(G8gat), .B(G36gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n257_), .B(KEYINPUT18), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G64gat), .B(G92gat), .ZN(new_n259_));
  XOR2_X1   g058(.A(new_n258_), .B(new_n259_), .Z(new_n260_));
  INV_X1    g059(.A(KEYINPUT20), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT25), .B(G183gat), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT26), .B(G190gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT81), .B(KEYINPUT23), .ZN(new_n265_));
  NAND2_X1  g064(.A1(G183gat), .A2(G190gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(new_n267_), .A2(KEYINPUT23), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n264_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G169gat), .ZN(new_n271_));
  INV_X1    g070(.A(G176gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n273_), .A2(KEYINPUT24), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(KEYINPUT24), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n274_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n270_), .A2(new_n278_), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT22), .B(G169gat), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n272_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n266_), .A2(KEYINPUT23), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n282_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284_));
  OAI211_X1 g083(.A(new_n275_), .B(new_n281_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n279_), .A2(new_n285_), .ZN(new_n286_));
  XOR2_X1   g085(.A(G211gat), .B(G218gat), .Z(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT92), .ZN(new_n288_));
  INV_X1    g087(.A(G197gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G204gat), .ZN(new_n290_));
  INV_X1    g089(.A(G204gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(G197gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n290_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G211gat), .B(G218gat), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT92), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n288_), .A2(KEYINPUT21), .A3(new_n293_), .A4(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(new_n290_), .A3(new_n292_), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n290_), .A2(new_n292_), .A3(KEYINPUT90), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT21), .B1(new_n290_), .B2(KEYINPUT90), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n299_), .B(new_n294_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n297_), .A2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n261_), .B1(new_n286_), .B2(new_n303_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n297_), .A2(new_n302_), .A3(KEYINPUT93), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT93), .B1(new_n297_), .B2(new_n302_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n277_), .A2(new_n283_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT25), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT79), .B1(new_n309_), .B2(G183gat), .ZN(new_n310_));
  OAI211_X1 g109(.A(new_n310_), .B(new_n263_), .C1(new_n262_), .C2(KEYINPUT79), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NOR2_X1   g112(.A1(new_n311_), .A2(new_n312_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n308_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT22), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT82), .B1(new_n316_), .B2(G169gat), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n272_), .B(new_n317_), .C1(new_n280_), .C2(KEYINPUT82), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n268_), .A2(new_n269_), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n275_), .B(new_n318_), .C1(new_n319_), .C2(new_n284_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n304_), .B1(new_n307_), .B2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT19), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n324_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n286_), .A2(new_n303_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n327_), .A2(new_n261_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n307_), .A2(new_n321_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n326_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  OAI211_X1 g129(.A(KEYINPUT32), .B(new_n260_), .C1(new_n325_), .C2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n322_), .A2(new_n324_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n303_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT94), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(new_n285_), .A4(new_n279_), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT94), .B1(new_n286_), .B2(new_n303_), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n324_), .A2(new_n261_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n329_), .A2(new_n335_), .A3(new_n336_), .A4(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n260_), .A2(KEYINPUT32), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n332_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n253_), .A2(new_n331_), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n260_), .B1(new_n332_), .B2(new_n338_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n332_), .A2(new_n338_), .A3(new_n260_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n342_), .B1(KEYINPUT95), .B2(new_n343_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(KEYINPUT96), .A2(KEYINPUT33), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n243_), .A2(new_n244_), .A3(new_n249_), .A4(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT95), .ZN(new_n348_));
  NAND4_X1  g147(.A1(new_n332_), .A2(new_n338_), .A3(new_n348_), .A4(new_n260_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n237_), .A2(new_n238_), .A3(new_n242_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n232_), .A2(new_n236_), .A3(new_n239_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n250_), .A3(new_n351_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n344_), .A2(new_n347_), .A3(new_n349_), .A4(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n252_), .A2(new_n345_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n341_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT29), .B1(new_n222_), .B2(new_n231_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT89), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G228gat), .A2(G233gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT89), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n240_), .A2(new_n360_), .A3(KEYINPUT29), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n358_), .A2(new_n359_), .A3(new_n361_), .A4(new_n307_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n357_), .A2(new_n303_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n363_), .A2(G228gat), .A3(G233gat), .ZN(new_n364_));
  XOR2_X1   g163(.A(G78gat), .B(G106gat), .Z(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n362_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n366_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT28), .B1(new_n240_), .B2(KEYINPUT29), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT28), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT29), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n234_), .A2(new_n371_), .A3(new_n372_), .A4(new_n221_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G22gat), .B(G50gat), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n370_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n375_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n377_));
  OAI22_X1  g176(.A1(new_n368_), .A2(new_n369_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n369_), .ZN(new_n379_));
  NOR2_X1   g178(.A1(new_n376_), .A2(new_n377_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n379_), .A2(new_n380_), .A3(new_n367_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n378_), .A2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n343_), .A2(KEYINPUT95), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n332_), .A2(new_n338_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n260_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n384_), .A2(new_n349_), .A3(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT27), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n386_), .B1(new_n325_), .B2(new_n330_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n343_), .A2(KEYINPUT27), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n388_), .A2(new_n389_), .B1(new_n390_), .B2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n253_), .B1(new_n378_), .B2(new_n381_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n356_), .A2(new_n383_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n321_), .B(KEYINPUT30), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G227gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(G15gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n396_), .B(new_n397_), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(G71gat), .ZN(new_n399_));
  INV_X1    g198(.A(G99gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n395_), .B(new_n401_), .ZN(new_n402_));
  XOR2_X1   g201(.A(KEYINPUT84), .B(KEYINPUT31), .Z(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT83), .B(G43gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n204_), .B(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n402_), .A2(new_n404_), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n405_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n407_), .B1(new_n405_), .B2(new_n408_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n256_), .B1(new_n394_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n392_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(new_n382_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n411_), .A2(new_n254_), .A3(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n409_), .A2(new_n410_), .ZN(new_n416_));
  AND3_X1   g215(.A1(new_n384_), .A2(new_n349_), .A3(new_n387_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n417_), .A2(new_n354_), .A3(new_n347_), .A4(new_n352_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n382_), .B1(new_n418_), .B2(new_n341_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n393_), .A2(new_n392_), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n416_), .B(KEYINPUT97), .C1(new_n419_), .C2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n412_), .A2(new_n415_), .A3(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G113gat), .B(G141gat), .Z(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT78), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G169gat), .B(G197gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n424_), .B(new_n425_), .Z(new_n426_));
  NAND2_X1  g225(.A1(G229gat), .A2(G233gat), .ZN(new_n427_));
  XOR2_X1   g226(.A(G15gat), .B(G22gat), .Z(new_n428_));
  NAND2_X1  g227(.A1(G1gat), .A2(G8gat), .ZN(new_n429_));
  AND2_X1   g228(.A1(new_n429_), .A2(KEYINPUT14), .ZN(new_n430_));
  OR3_X1    g229(.A1(new_n428_), .A2(KEYINPUT75), .A3(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n429_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(G1gat), .A2(G8gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  OAI21_X1  g233(.A(KEYINPUT75), .B1(new_n428_), .B2(new_n430_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n431_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n434_), .B1(new_n431_), .B2(new_n435_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G29gat), .B(G36gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G43gat), .B(G50gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n439_), .B(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n438_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n441_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n443_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT77), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n442_), .A2(KEYINPUT77), .A3(new_n444_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n427_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n441_), .B(KEYINPUT15), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n442_), .A2(new_n450_), .A3(new_n427_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n426_), .B1(new_n448_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n426_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n447_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n455_), .A2(new_n445_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n451_), .B(new_n454_), .C1(new_n456_), .C2(new_n427_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n422_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G232gat), .A2(G233gat), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(KEYINPUT34), .Z(new_n461_));
  INV_X1    g260(.A(KEYINPUT35), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n462_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT71), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT72), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G92gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n470_), .A2(KEYINPUT9), .ZN(new_n471_));
  AND2_X1   g270(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n471_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(G85gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n470_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G85gat), .A2(G92gat), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n476_), .A2(KEYINPUT9), .A3(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(KEYINPUT66), .B1(new_n474_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n474_), .A2(new_n478_), .A3(KEYINPUT66), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT6), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT6), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n485_), .A2(G99gat), .A3(G106gat), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  OR2_X1    g286(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT64), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n488_), .A2(KEYINPUT64), .A3(new_n489_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G106gat), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n487_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT67), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n476_), .A2(new_n497_), .A3(new_n477_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT7), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n499_), .A2(new_n400_), .A3(new_n495_), .ZN(new_n500_));
  OAI21_X1  g299(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n498_), .B1(new_n487_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT8), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n484_), .A2(new_n486_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(new_n501_), .A3(new_n500_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT8), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n507_), .A3(new_n498_), .ZN(new_n508_));
  AOI22_X1  g307(.A1(new_n482_), .A2(new_n496_), .B1(new_n504_), .B2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(KEYINPUT70), .B1(new_n509_), .B2(new_n441_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n504_), .A2(new_n508_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n488_), .A2(KEYINPUT64), .A3(new_n489_), .ZN(new_n512_));
  AOI21_X1  g311(.A(KEYINPUT64), .B1(new_n488_), .B2(new_n489_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n495_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n474_), .A2(KEYINPUT66), .A3(new_n478_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n514_), .B(new_n505_), .C1(new_n515_), .C2(new_n479_), .ZN(new_n516_));
  AND4_X1   g315(.A1(KEYINPUT70), .A2(new_n511_), .A3(new_n441_), .A4(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n469_), .B1(new_n510_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n449_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT69), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n476_), .A2(new_n497_), .A3(new_n477_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n500_), .A2(new_n501_), .ZN(new_n522_));
  AOI211_X1 g321(.A(KEYINPUT8), .B(new_n521_), .C1(new_n522_), .C2(new_n505_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n507_), .B1(new_n506_), .B2(new_n498_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n520_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n504_), .A2(KEYINPUT69), .A3(new_n508_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n519_), .B1(new_n527_), .B2(new_n516_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n463_), .B1(new_n518_), .B2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G190gat), .B(G218gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G134gat), .B(G162gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(KEYINPUT36), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT70), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n515_), .A2(new_n479_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n514_), .A2(new_n505_), .ZN(new_n536_));
  OAI22_X1  g335(.A1(new_n535_), .A2(new_n536_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n534_), .B1(new_n537_), .B2(new_n443_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n509_), .A2(KEYINPUT70), .A3(new_n441_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n468_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(new_n463_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n527_), .A2(new_n516_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n449_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n540_), .A2(new_n541_), .A3(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n529_), .A2(new_n533_), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT73), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n529_), .A2(KEYINPUT73), .A3(new_n544_), .A4(new_n533_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n532_), .B(KEYINPUT36), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n550_), .B1(new_n529_), .B2(new_n544_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT74), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n554_), .A2(KEYINPUT37), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(KEYINPUT37), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n553_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT17), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n438_), .B(new_n560_), .Z(new_n561_));
  INV_X1    g360(.A(KEYINPUT11), .ZN(new_n562_));
  INV_X1    g361(.A(G57gat), .ZN(new_n563_));
  NOR2_X1   g362(.A1(new_n563_), .A2(G64gat), .ZN(new_n564_));
  INV_X1    g363(.A(G64gat), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n565_), .A2(G57gat), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n562_), .B1(new_n564_), .B2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(G57gat), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n563_), .A2(G64gat), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(KEYINPUT11), .ZN(new_n570_));
  INV_X1    g369(.A(G78gat), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(G71gat), .ZN(new_n572_));
  INV_X1    g371(.A(G71gat), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(G78gat), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n567_), .A2(new_n570_), .A3(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G57gat), .B(G64gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G71gat), .B(G78gat), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(KEYINPUT11), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n561_), .A2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n561_), .A2(new_n580_), .ZN(new_n582_));
  XOR2_X1   g381(.A(G127gat), .B(G155gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(G183gat), .B(G211gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n583_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  OR4_X1    g386(.A1(new_n559_), .A2(new_n581_), .A3(new_n582_), .A4(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n580_), .A2(KEYINPUT68), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT68), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n570_), .A2(new_n575_), .ZN(new_n591_));
  AOI21_X1  g390(.A(KEYINPUT11), .B1(new_n568_), .B2(new_n569_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n590_), .B(new_n579_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n589_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n561_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n587_), .B(KEYINPUT17), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n588_), .A2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n551_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(new_n554_), .A3(KEYINPUT37), .ZN(new_n600_));
  INV_X1    g399(.A(new_n593_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n590_), .B1(new_n576_), .B2(new_n579_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT12), .B1(new_n537_), .B2(new_n603_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n537_), .A2(new_n603_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n576_), .A2(KEYINPUT12), .A3(new_n579_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n542_), .A2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n606_), .A2(new_n609_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n610_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n509_), .A2(new_n594_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n612_), .B1(new_n613_), .B2(new_n605_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT5), .ZN(new_n617_));
  XNOR2_X1  g416(.A(G176gat), .B(G204gat), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n617_), .B(new_n618_), .Z(new_n619_));
  NAND2_X1  g418(.A1(new_n615_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n619_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n611_), .A2(new_n614_), .A3(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT13), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n558_), .A2(new_n598_), .A3(new_n600_), .A4(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n459_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT98), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n459_), .A2(new_n629_), .A3(new_n626_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n628_), .A2(KEYINPUT99), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(KEYINPUT99), .B1(new_n628_), .B2(new_n630_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n255_), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT38), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  OAI211_X1 g435(.A(KEYINPUT38), .B(new_n255_), .C1(new_n632_), .C2(new_n633_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n624_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n458_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n598_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT100), .Z(new_n642_));
  NAND3_X1  g441(.A1(new_n642_), .A2(new_n422_), .A3(new_n553_), .ZN(new_n643_));
  OAI21_X1  g442(.A(G1gat), .B1(new_n643_), .B2(new_n254_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT101), .Z(new_n645_));
  NAND3_X1  g444(.A1(new_n636_), .A2(new_n637_), .A3(new_n645_), .ZN(G1324gat));
  INV_X1    g445(.A(KEYINPUT40), .ZN(new_n647_));
  OAI21_X1  g446(.A(G8gat), .B1(new_n643_), .B2(new_n392_), .ZN(new_n648_));
  XOR2_X1   g447(.A(new_n648_), .B(KEYINPUT39), .Z(new_n649_));
  OR2_X1    g448(.A1(new_n392_), .A2(G8gat), .ZN(new_n650_));
  INV_X1    g449(.A(new_n633_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n651_), .B2(new_n631_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n647_), .B1(new_n649_), .B2(new_n652_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n648_), .B(KEYINPUT39), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n632_), .A2(new_n633_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n654_), .B(KEYINPUT40), .C1(new_n655_), .C2(new_n650_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n653_), .A2(new_n656_), .ZN(G1325gat));
  OAI21_X1  g456(.A(G15gat), .B1(new_n643_), .B2(new_n416_), .ZN(new_n658_));
  XOR2_X1   g457(.A(new_n658_), .B(KEYINPUT41), .Z(new_n659_));
  NAND4_X1  g458(.A1(new_n628_), .A2(new_n397_), .A3(new_n411_), .A4(new_n630_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT102), .ZN(new_n661_));
  OR2_X1    g460(.A1(new_n660_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n661_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n659_), .A2(new_n662_), .A3(new_n663_), .ZN(G1326gat));
  XNOR2_X1  g463(.A(new_n382_), .B(KEYINPUT103), .ZN(new_n665_));
  OAI21_X1  g464(.A(G22gat), .B1(new_n643_), .B2(new_n665_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT42), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n628_), .A2(new_n630_), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n665_), .A2(G22gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n667_), .B1(new_n668_), .B2(new_n669_), .ZN(G1327gat));
  INV_X1    g469(.A(new_n598_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n640_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n558_), .A2(new_n600_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(KEYINPUT43), .B1(new_n675_), .B2(KEYINPUT104), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n421_), .A2(new_n415_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n384_), .A2(new_n387_), .A3(new_n349_), .A4(new_n352_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n347_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n678_), .A2(new_n355_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n341_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n383_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n393_), .A2(new_n392_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT97), .B1(new_n684_), .B2(new_n416_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n674_), .B(new_n676_), .C1(new_n677_), .C2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n676_), .B1(new_n422_), .B2(new_n674_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT44), .B(new_n673_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT105), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n674_), .B1(new_n677_), .B2(new_n685_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n676_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(new_n686_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT105), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(KEYINPUT44), .A4(new_n673_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n690_), .A2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n694_), .A2(new_n673_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT44), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND4_X1  g499(.A1(new_n697_), .A2(G29gat), .A3(new_n253_), .A4(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n671_), .A2(new_n599_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n702_), .A2(new_n638_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n422_), .A2(new_n458_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G29gat), .B1(new_n705_), .B2(new_n253_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n701_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT106), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT106), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n701_), .A2(new_n710_), .A3(new_n707_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n709_), .A2(new_n711_), .ZN(G1328gat));
  OAI21_X1  g511(.A(KEYINPUT109), .B1(KEYINPUT108), .B2(KEYINPUT46), .ZN(new_n713_));
  INV_X1    g512(.A(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(G36gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n392_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n697_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n392_), .A2(G36gat), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n459_), .A2(new_n718_), .A3(new_n703_), .A4(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT45), .ZN(new_n721_));
  INV_X1    g520(.A(new_n719_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT107), .B1(new_n704_), .B2(new_n722_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n720_), .A2(new_n721_), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n721_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n726_));
  OAI22_X1  g525(.A1(new_n725_), .A2(new_n726_), .B1(KEYINPUT109), .B2(KEYINPUT46), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n714_), .B1(new_n717_), .B2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n720_), .A2(new_n723_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(KEYINPUT45), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(new_n731_), .B2(new_n724_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n672_), .B1(new_n693_), .B2(new_n686_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n413_), .B1(new_n733_), .B2(KEYINPUT44), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n734_), .B1(new_n690_), .B2(new_n696_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n732_), .B(new_n713_), .C1(new_n735_), .C2(new_n715_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n728_), .A2(new_n736_), .ZN(G1329gat));
  NAND4_X1  g536(.A1(new_n697_), .A2(G43gat), .A3(new_n411_), .A4(new_n700_), .ZN(new_n738_));
  AOI21_X1  g537(.A(G43gat), .B1(new_n705_), .B2(new_n411_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT47), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n738_), .A2(new_n743_), .A3(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(G1330gat));
  INV_X1    g544(.A(G50gat), .ZN(new_n746_));
  INV_X1    g545(.A(new_n665_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n705_), .A2(new_n746_), .A3(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT110), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n383_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n697_), .A2(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n751_), .B2(G50gat), .ZN(new_n752_));
  AOI211_X1 g551(.A(KEYINPUT110), .B(new_n746_), .C1(new_n697_), .C2(new_n750_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n748_), .B1(new_n752_), .B2(new_n753_), .ZN(G1331gat));
  AND2_X1   g553(.A1(new_n422_), .A2(new_n639_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n755_), .A2(new_n675_), .A3(new_n598_), .A4(new_n638_), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n756_), .B(KEYINPUT111), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n757_), .A2(new_n563_), .A3(new_n253_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n624_), .A2(new_n458_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n422_), .A2(new_n553_), .A3(new_n598_), .A4(new_n759_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT112), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(new_n253_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(G57gat), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n758_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n758_), .A2(KEYINPUT113), .A3(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1332gat));
  NAND3_X1  g567(.A1(new_n757_), .A2(new_n565_), .A3(new_n413_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n761_), .A2(new_n413_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(G64gat), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n771_), .A2(KEYINPUT48), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(KEYINPUT48), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(G1333gat));
  NAND3_X1  g573(.A1(new_n757_), .A2(new_n573_), .A3(new_n411_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n761_), .A2(new_n411_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(G71gat), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n777_), .A2(KEYINPUT49), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n777_), .A2(KEYINPUT49), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1334gat));
  NAND3_X1  g579(.A1(new_n757_), .A2(new_n571_), .A3(new_n747_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n761_), .A2(new_n747_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(G78gat), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n783_), .A2(KEYINPUT50), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(KEYINPUT50), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(G1335gat));
  NAND2_X1  g585(.A1(new_n759_), .A2(new_n671_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n693_), .B2(new_n686_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n472_), .A2(new_n473_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n254_), .A2(new_n789_), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n702_), .A2(new_n624_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n755_), .A2(new_n253_), .A3(new_n791_), .ZN(new_n792_));
  AOI22_X1  g591(.A1(new_n788_), .A2(new_n790_), .B1(new_n792_), .B2(new_n475_), .ZN(G1336gat));
  AND2_X1   g592(.A1(new_n788_), .A2(new_n413_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n755_), .A2(new_n791_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n413_), .A2(new_n470_), .ZN(new_n796_));
  OAI22_X1  g595(.A1(new_n794_), .A2(new_n470_), .B1(new_n795_), .B2(new_n796_), .ZN(G1337gat));
  INV_X1    g596(.A(new_n494_), .ZN(new_n798_));
  NOR3_X1   g597(.A1(new_n795_), .A2(new_n416_), .A3(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT114), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n400_), .B1(new_n788_), .B2(new_n411_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  OR3_X1    g602(.A1(new_n800_), .A2(new_n801_), .A3(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n803_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(G1338gat));
  AOI211_X1 g605(.A(KEYINPUT116), .B(new_n495_), .C1(new_n788_), .C2(new_n382_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n808_));
  INV_X1    g607(.A(new_n787_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n694_), .A2(new_n382_), .A3(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n808_), .B1(new_n810_), .B2(G106gat), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n807_), .A2(new_n811_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(G106gat), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n814_), .A2(KEYINPUT116), .A3(new_n812_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n795_), .A2(G106gat), .A3(new_n383_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT53), .B1(new_n813_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n816_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n811_), .A2(new_n812_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n820_), .B(new_n821_), .C1(new_n822_), .C2(new_n807_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n819_), .A2(new_n823_), .ZN(G1339gat));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n607_), .B1(new_n527_), .B2(new_n516_), .ZN(new_n826_));
  NOR4_X1   g625(.A1(new_n826_), .A2(new_n604_), .A3(new_n605_), .A4(new_n612_), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT12), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n828_), .B1(new_n509_), .B2(new_n594_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n509_), .A2(new_n594_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n612_), .B1(new_n831_), .B2(new_n826_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n827_), .B1(KEYINPUT55), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT55), .ZN(new_n834_));
  NOR4_X1   g633(.A1(new_n831_), .A2(new_n826_), .A3(new_n834_), .A4(new_n612_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n619_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT56), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT56), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n838_), .B(new_n619_), .C1(new_n833_), .C2(new_n835_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n837_), .A2(new_n458_), .A3(new_n622_), .A4(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n427_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n454_), .B1(new_n841_), .B2(new_n450_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n427_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n842_), .B1(new_n456_), .B2(new_n843_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n457_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(new_n623_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n840_), .A2(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n825_), .B1(new_n847_), .B2(new_n599_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n599_), .B1(new_n840_), .B2(new_n846_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(KEYINPUT57), .ZN(new_n850_));
  INV_X1    g649(.A(new_n622_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n836_), .B2(KEYINPUT56), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n852_), .A2(new_n845_), .A3(new_n839_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n852_), .A2(KEYINPUT58), .A3(new_n845_), .A4(new_n839_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n674_), .A3(new_n856_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n848_), .A2(new_n850_), .A3(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(KEYINPUT54), .B1(new_n625_), .B2(new_n458_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT54), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n626_), .A2(new_n860_), .A3(new_n639_), .ZN(new_n861_));
  AOI22_X1  g660(.A1(new_n858_), .A2(new_n671_), .B1(new_n859_), .B2(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n411_), .A2(new_n253_), .A3(new_n414_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT117), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  NAND4_X1  g664(.A1(new_n411_), .A2(KEYINPUT117), .A3(new_n253_), .A4(new_n414_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n862_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(G113gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n869_), .A3(new_n458_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n599_), .A2(new_n554_), .A3(KEYINPUT37), .ZN(new_n872_));
  INV_X1    g671(.A(new_n557_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n599_), .A2(new_n555_), .A3(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n856_), .B1(new_n872_), .B2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n610_), .B1(new_n606_), .B2(new_n609_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n611_), .B1(new_n876_), .B2(new_n834_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n835_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n621_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n622_), .B1(new_n879_), .B2(new_n838_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n839_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n880_), .A2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(KEYINPUT58), .B1(new_n882_), .B2(new_n845_), .ZN(new_n883_));
  OAI22_X1  g682(.A1(new_n875_), .A2(new_n883_), .B1(new_n849_), .B2(KEYINPUT57), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n849_), .A2(KEYINPUT57), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n671_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n861_), .A2(new_n859_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(new_n867_), .ZN(new_n889_));
  AOI21_X1  g688(.A(KEYINPUT59), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT59), .ZN(new_n891_));
  AOI211_X1 g690(.A(new_n891_), .B(new_n867_), .C1(new_n886_), .C2(new_n887_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n871_), .B1(new_n890_), .B2(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n891_), .B1(new_n862_), .B2(new_n867_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n888_), .A2(KEYINPUT59), .A3(new_n889_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n894_), .A2(new_n895_), .A3(KEYINPUT118), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n893_), .A2(new_n896_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n897_), .A2(new_n458_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n870_), .B1(new_n898_), .B2(new_n869_), .ZN(G1340gat));
  INV_X1    g698(.A(G120gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n900_), .B1(new_n624_), .B2(KEYINPUT60), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n868_), .B(new_n901_), .C1(KEYINPUT60), .C2(new_n900_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n624_), .B1(new_n894_), .B2(new_n895_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n902_), .B1(new_n903_), .B2(new_n900_), .ZN(G1341gat));
  NAND3_X1  g703(.A1(new_n893_), .A2(new_n598_), .A3(new_n896_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(G127gat), .ZN(new_n906_));
  INV_X1    g705(.A(G127gat), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n868_), .A2(new_n907_), .A3(new_n598_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n906_), .A2(KEYINPUT119), .A3(new_n908_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1342gat));
  AOI21_X1  g712(.A(G134gat), .B1(new_n868_), .B2(new_n599_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n674_), .A2(G134gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n915_), .B(KEYINPUT120), .ZN(new_n916_));
  AOI21_X1  g715(.A(new_n914_), .B1(new_n897_), .B2(new_n916_), .ZN(G1343gat));
  NAND4_X1  g716(.A1(new_n416_), .A2(new_n382_), .A3(new_n253_), .A4(new_n392_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(KEYINPUT121), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n888_), .A2(new_n919_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(new_n920_), .A2(new_n639_), .ZN(new_n921_));
  XOR2_X1   g720(.A(new_n921_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g721(.A1(new_n920_), .A2(new_n624_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(KEYINPUT122), .B(G148gat), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n923_), .B(new_n924_), .ZN(G1345gat));
  NOR2_X1   g724(.A1(new_n920_), .A2(new_n671_), .ZN(new_n926_));
  XOR2_X1   g725(.A(KEYINPUT61), .B(G155gat), .Z(new_n927_));
  XNOR2_X1  g726(.A(new_n926_), .B(new_n927_), .ZN(G1346gat));
  OAI21_X1  g727(.A(new_n216_), .B1(new_n920_), .B2(new_n553_), .ZN(new_n929_));
  XOR2_X1   g728(.A(new_n929_), .B(KEYINPUT123), .Z(new_n930_));
  NOR3_X1   g729(.A1(new_n920_), .A2(new_n216_), .A3(new_n675_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1347gat));
  NAND3_X1  g731(.A1(new_n411_), .A2(new_n254_), .A3(new_n413_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n862_), .A2(new_n747_), .A3(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n271_), .B1(new_n934_), .B2(new_n458_), .ZN(new_n935_));
  OR2_X1    g734(.A1(new_n935_), .A2(KEYINPUT62), .ZN(new_n936_));
  NAND3_X1  g735(.A1(new_n934_), .A2(new_n458_), .A3(new_n280_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n935_), .A2(KEYINPUT62), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n936_), .A2(new_n937_), .A3(new_n938_), .ZN(G1348gat));
  AOI21_X1  g738(.A(G176gat), .B1(new_n934_), .B2(new_n638_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n862_), .A2(new_n382_), .ZN(new_n941_));
  NOR3_X1   g740(.A1(new_n933_), .A2(new_n272_), .A3(new_n624_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n940_), .B1(new_n941_), .B2(new_n942_), .ZN(G1349gat));
  NOR2_X1   g742(.A1(new_n671_), .A2(new_n262_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n934_), .A2(new_n944_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n945_), .A2(KEYINPUT124), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n945_), .A2(KEYINPUT124), .ZN(new_n947_));
  NOR2_X1   g746(.A1(new_n933_), .A2(new_n671_), .ZN(new_n948_));
  AOI21_X1  g747(.A(G183gat), .B1(new_n941_), .B2(new_n948_), .ZN(new_n949_));
  NOR3_X1   g748(.A1(new_n946_), .A2(new_n947_), .A3(new_n949_), .ZN(G1350gat));
  NAND2_X1  g749(.A1(new_n934_), .A2(new_n674_), .ZN(new_n951_));
  AND2_X1   g750(.A1(new_n599_), .A2(new_n263_), .ZN(new_n952_));
  AOI22_X1  g751(.A1(new_n951_), .A2(G190gat), .B1(new_n934_), .B2(new_n952_), .ZN(new_n953_));
  XOR2_X1   g752(.A(new_n953_), .B(KEYINPUT125), .Z(G1351gat));
  NAND4_X1  g753(.A1(new_n888_), .A2(new_n416_), .A3(new_n413_), .A4(new_n393_), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT126), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n955_), .B(new_n956_), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n957_), .A2(new_n458_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g758(.A1(new_n957_), .A2(new_n638_), .ZN(new_n960_));
  XNOR2_X1  g759(.A(new_n960_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g760(.A(new_n955_), .B(KEYINPUT126), .ZN(new_n962_));
  NOR2_X1   g761(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n963_));
  AND2_X1   g762(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n964_));
  NOR4_X1   g763(.A1(new_n962_), .A2(new_n671_), .A3(new_n963_), .A4(new_n964_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n957_), .A2(new_n598_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n965_), .B1(new_n966_), .B2(new_n963_), .ZN(G1354gat));
  NOR3_X1   g766(.A1(new_n962_), .A2(G218gat), .A3(new_n553_), .ZN(new_n968_));
  INV_X1    g767(.A(G218gat), .ZN(new_n969_));
  AOI21_X1  g768(.A(new_n969_), .B1(new_n957_), .B2(new_n674_), .ZN(new_n970_));
  OAI21_X1  g769(.A(KEYINPUT127), .B1(new_n968_), .B2(new_n970_), .ZN(new_n971_));
  OAI21_X1  g770(.A(G218gat), .B1(new_n962_), .B2(new_n675_), .ZN(new_n972_));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n957_), .A2(new_n969_), .A3(new_n599_), .ZN(new_n974_));
  NAND3_X1  g773(.A1(new_n972_), .A2(new_n973_), .A3(new_n974_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n971_), .A2(new_n975_), .ZN(G1355gat));
endmodule


