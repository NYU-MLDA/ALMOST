//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n656_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n857_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n895_, new_n896_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n927_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT20), .ZN(new_n205_));
  INV_X1    g004(.A(G183gat), .ZN(new_n206_));
  INV_X1    g005(.A(G190gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT23), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT83), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G169gat), .ZN(new_n214_));
  INV_X1    g013(.A(G176gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT24), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n215_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT25), .B(G183gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT26), .B(G190gat), .ZN(new_n221_));
  AOI22_X1  g020(.A1(new_n218_), .A2(new_n219_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n217_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n213_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n208_), .A2(new_n212_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT22), .B(G169gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n216_), .B1(new_n229_), .B2(new_n215_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n224_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G204gat), .ZN(new_n233_));
  OR3_X1    g032(.A1(new_n233_), .A2(KEYINPUT90), .A3(G197gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(KEYINPUT90), .B1(new_n233_), .B2(G197gat), .ZN(new_n235_));
  INV_X1    g034(.A(G197gat), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n234_), .B(new_n235_), .C1(new_n236_), .C2(G204gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT21), .ZN(new_n238_));
  XNOR2_X1  g037(.A(G211gat), .B(G218gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT91), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n240_), .B1(G197gat), .B2(new_n233_), .ZN(new_n241_));
  NOR3_X1   g040(.A1(new_n236_), .A2(KEYINPUT91), .A3(G204gat), .ZN(new_n242_));
  OAI22_X1  g041(.A1(new_n241_), .A2(new_n242_), .B1(G197gat), .B2(new_n233_), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n238_), .B(new_n239_), .C1(new_n243_), .C2(KEYINPUT21), .ZN(new_n244_));
  INV_X1    g043(.A(new_n239_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(KEYINPUT21), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n205_), .B1(new_n232_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n225_), .A2(new_n223_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT94), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n249_), .B(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(new_n222_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT95), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n251_), .A2(KEYINPUT95), .A3(new_n222_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n213_), .A2(new_n227_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(new_n230_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n204_), .B(new_n248_), .C1(new_n259_), .C2(new_n247_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT20), .B1(new_n232_), .B2(new_n247_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n261_), .B1(new_n259_), .B2(new_n247_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n260_), .B1(new_n262_), .B2(new_n204_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G8gat), .B(G36gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT18), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G64gat), .B(G92gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n263_), .A2(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n260_), .B(new_n267_), .C1(new_n262_), .C2(new_n204_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT27), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n252_), .A2(new_n258_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n248_), .B1(new_n247_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n203_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n261_), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n254_), .A2(new_n255_), .B1(new_n230_), .B2(new_n257_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n247_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n277_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n276_), .B1(new_n280_), .B2(new_n203_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n268_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(new_n270_), .A3(KEYINPUT27), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT99), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285_));
  OR2_X1    g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT86), .ZN(new_n287_));
  OR4_X1    g086(.A1(new_n287_), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n288_));
  INV_X1    g087(.A(G141gat), .ZN(new_n289_));
  INV_X1    g088(.A(G148gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT87), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT2), .ZN(new_n292_));
  OAI22_X1  g091(.A1(new_n287_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n288_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n291_), .A2(KEYINPUT2), .ZN(new_n295_));
  OAI211_X1 g094(.A(new_n285_), .B(new_n286_), .C1(new_n294_), .C2(new_n295_), .ZN(new_n296_));
  AND3_X1   g095(.A1(new_n285_), .A2(KEYINPUT85), .A3(KEYINPUT1), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT85), .B1(new_n285_), .B2(KEYINPUT1), .ZN(new_n298_));
  OAI221_X1 g097(.A(new_n286_), .B1(KEYINPUT1), .B2(new_n285_), .C1(new_n297_), .C2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G141gat), .B(G148gat), .Z(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n296_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G127gat), .B(G134gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(G113gat), .B(G120gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n303_), .B(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n296_), .A2(new_n301_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT84), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n308_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n305_), .B2(new_n308_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(G225gat), .A2(G233gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n306_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT4), .B1(new_n307_), .B2(new_n310_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n306_), .A2(new_n311_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n314_), .B1(new_n315_), .B2(KEYINPUT4), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n312_), .B(KEYINPUT96), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n313_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(G1gat), .B(G29gat), .Z(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G57gat), .B(G85gat), .ZN(new_n323_));
  XOR2_X1   g122(.A(new_n322_), .B(new_n323_), .Z(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n319_), .A2(new_n325_), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n313_), .B(new_n324_), .C1(new_n316_), .C2(new_n318_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT99), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n282_), .A2(new_n270_), .A3(new_n330_), .A4(KEYINPUT27), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n273_), .A2(new_n284_), .A3(new_n329_), .A4(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G71gat), .B(G99gat), .ZN(new_n334_));
  XOR2_X1   g133(.A(new_n334_), .B(G43gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(new_n232_), .B(new_n335_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(new_n310_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(G227gat), .A2(G233gat), .ZN(new_n338_));
  INV_X1    g137(.A(G15gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT30), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT31), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n337_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n307_), .A2(KEYINPUT29), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(KEYINPUT89), .A3(new_n247_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G228gat), .A2(G233gat), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n346_), .B(KEYINPUT88), .Z(new_n347_));
  INV_X1    g146(.A(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n345_), .A2(new_n348_), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n344_), .A2(KEYINPUT89), .A3(new_n247_), .A4(new_n347_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(G78gat), .B(G106gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n349_), .A2(new_n350_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT92), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT92), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n349_), .A2(new_n354_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n349_), .A2(new_n350_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n351_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n353_), .A2(new_n355_), .A3(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n302_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT28), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G22gat), .B(G50gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n362_), .B(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT93), .B1(new_n359_), .B2(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n359_), .A2(new_n365_), .A3(KEYINPUT93), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n365_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(new_n352_), .A3(new_n358_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n343_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n368_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n343_), .B(new_n371_), .C1(new_n373_), .C2(new_n366_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n333_), .B1(new_n372_), .B2(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n371_), .B1(new_n373_), .B2(new_n366_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n343_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n281_), .A2(KEYINPUT32), .A3(new_n267_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n267_), .A2(KEYINPUT32), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n260_), .B(new_n381_), .C1(new_n262_), .C2(new_n204_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n328_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT33), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n327_), .A2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n318_), .B1(new_n315_), .B2(KEYINPUT98), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n386_), .B1(KEYINPUT98), .B2(new_n315_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n312_), .ZN(new_n388_));
  OAI211_X1 g187(.A(new_n387_), .B(new_n325_), .C1(new_n388_), .C2(new_n316_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n327_), .A2(new_n384_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n385_), .A2(new_n389_), .A3(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n383_), .B1(new_n391_), .B2(new_n271_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n378_), .A2(new_n379_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n376_), .A2(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G15gat), .B(G22gat), .ZN(new_n395_));
  INV_X1    g194(.A(G1gat), .ZN(new_n396_));
  INV_X1    g195(.A(G8gat), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT14), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n395_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G1gat), .B(G8gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G29gat), .B(G36gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G43gat), .B(G50gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n402_), .B(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n401_), .B(new_n404_), .Z(new_n405_));
  NAND2_X1  g204(.A1(G229gat), .A2(G233gat), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT81), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n404_), .B(KEYINPUT15), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n401_), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n411_), .B(KEYINPUT82), .Z(new_n412_));
  INV_X1    g211(.A(new_n401_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n404_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(new_n407_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n409_), .B1(new_n412_), .B2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G113gat), .B(G141gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G169gat), .B(G197gat), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n418_), .B(new_n419_), .Z(new_n420_));
  XNOR2_X1  g219(.A(new_n417_), .B(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n394_), .A2(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G183gat), .B(G211gat), .Z(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT80), .ZN(new_n424_));
  XOR2_X1   g223(.A(G127gat), .B(G155gat), .Z(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XOR2_X1   g225(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n427_));
  XNOR2_X1  g226(.A(new_n426_), .B(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT17), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n429_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G231gat), .A2(G233gat), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n401_), .B(new_n433_), .Z(new_n434_));
  INV_X1    g233(.A(G64gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(G57gat), .ZN(new_n436_));
  INV_X1    g235(.A(G57gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(G64gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT69), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n439_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT11), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n437_), .A2(G64gat), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n435_), .A2(G57gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT69), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT11), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n436_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G71gat), .B(G78gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n442_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  OAI211_X1 g250(.A(KEYINPUT11), .B(new_n449_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n434_), .B(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n431_), .A2(new_n432_), .A3(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT70), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n453_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n451_), .A2(KEYINPUT70), .A3(new_n452_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(new_n434_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n461_), .A2(new_n434_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n430_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n456_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT67), .ZN(new_n466_));
  INV_X1    g265(.A(G99gat), .ZN(new_n467_));
  INV_X1    g266(.A(G106gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT7), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n467_), .B(new_n468_), .C1(new_n469_), .C2(KEYINPUT66), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT66), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n471_), .A2(KEYINPUT7), .ZN(new_n472_));
  OAI21_X1  g271(.A(new_n466_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n469_), .A2(KEYINPUT66), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n471_), .A2(KEYINPUT7), .ZN(new_n475_));
  NOR2_X1   g274(.A1(G99gat), .A2(G106gat), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n474_), .A2(new_n475_), .A3(KEYINPUT67), .A4(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n473_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G99gat), .A2(G106gat), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n481_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n478_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(G85gat), .ZN(new_n487_));
  INV_X1    g286(.A(G92gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(G85gat), .A2(G92gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n492_), .B1(KEYINPUT68), .B2(KEYINPUT8), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n486_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT8), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT68), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n481_), .A2(new_n497_), .A3(new_n482_), .A4(new_n483_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n498_), .B1(new_n473_), .B2(new_n477_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n496_), .B1(new_n499_), .B2(new_n491_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT10), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n467_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n502_), .A2(new_n468_), .A3(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT64), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT65), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n506_), .A2(KEYINPUT9), .A3(G85gat), .A4(G92gat), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n507_), .A2(new_n481_), .A3(new_n483_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n491_), .A2(KEYINPUT9), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT9), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n506_), .B1(new_n490_), .B2(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n508_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n505_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n495_), .A2(new_n500_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(new_n410_), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n515_), .A2(KEYINPUT75), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(KEYINPUT75), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n498_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n478_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(KEYINPUT8), .B1(new_n520_), .B2(new_n492_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT64), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n504_), .B(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n481_), .A2(new_n483_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n510_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n511_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n524_), .B(new_n507_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n484_), .B1(new_n473_), .B2(new_n477_), .ZN(new_n528_));
  OAI22_X1  g327(.A1(new_n523_), .A2(new_n527_), .B1(new_n528_), .B2(new_n493_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n521_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(new_n404_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n518_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT76), .B1(new_n516_), .B2(new_n517_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G232gat), .A2(G233gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(KEYINPUT35), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n532_), .B1(new_n533_), .B2(new_n537_), .ZN(new_n538_));
  XOR2_X1   g337(.A(G134gat), .B(G162gat), .Z(new_n539_));
  XNOR2_X1  g338(.A(G190gat), .B(G218gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT36), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n536_), .A2(KEYINPUT35), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT76), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n518_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n537_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n543_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n538_), .B(new_n542_), .C1(new_n547_), .C2(new_n532_), .ZN(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(KEYINPUT77), .B(KEYINPUT36), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n541_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT78), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n532_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n533_), .A2(new_n537_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n554_), .B1(new_n555_), .B2(new_n543_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n553_), .B1(new_n556_), .B2(new_n538_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT37), .B1(new_n549_), .B2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n538_), .B1(new_n547_), .B2(new_n532_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n552_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n548_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n465_), .B1(new_n558_), .B2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT12), .B1(new_n521_), .B2(new_n529_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT71), .B1(new_n460_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n486_), .A2(new_n494_), .B1(new_n505_), .B2(new_n512_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n566_), .B1(new_n567_), .B2(new_n500_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT71), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n458_), .A4(new_n459_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n514_), .A2(new_n454_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n571_), .A2(new_n566_), .ZN(new_n572_));
  AND2_X1   g371(.A1(G230gat), .A2(G233gat), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n573_), .B1(new_n530_), .B2(new_n453_), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n565_), .A2(new_n570_), .A3(new_n572_), .A4(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT72), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n530_), .A2(new_n453_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n571_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(new_n573_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n458_), .A2(new_n514_), .A3(KEYINPUT12), .A4(new_n459_), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n581_), .A2(KEYINPUT71), .B1(new_n566_), .B2(new_n571_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n582_), .A2(KEYINPUT72), .A3(new_n570_), .A4(new_n574_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n577_), .A2(new_n580_), .A3(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G120gat), .B(G148gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(G176gat), .B(G204gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n584_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n584_), .A2(new_n589_), .ZN(new_n591_));
  AND3_X1   g390(.A1(new_n590_), .A2(KEYINPUT13), .A3(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(KEYINPUT13), .B1(new_n590_), .B2(new_n591_), .ZN(new_n593_));
  NOR2_X1   g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n563_), .A2(new_n594_), .ZN(new_n595_));
  OR3_X1    g394(.A1(new_n422_), .A2(KEYINPUT100), .A3(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT100), .B1(new_n422_), .B2(new_n595_), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n598_), .A2(new_n396_), .A3(new_n328_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT38), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n377_), .A2(new_n379_), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n332_), .B1(new_n602_), .B2(new_n374_), .ZN(new_n603_));
  AND4_X1   g402(.A1(new_n379_), .A2(new_n392_), .A3(new_n369_), .A4(new_n371_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n560_), .A2(new_n548_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n465_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n594_), .A2(new_n421_), .A3(new_n611_), .ZN(new_n612_));
  OR2_X1    g411(.A1(new_n612_), .A2(KEYINPUT101), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(KEYINPUT101), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n610_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OAI21_X1  g415(.A(G1gat), .B1(new_n616_), .B2(new_n329_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n599_), .A2(new_n600_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n601_), .A2(new_n617_), .A3(new_n618_), .ZN(G1324gat));
  AND2_X1   g418(.A1(new_n273_), .A2(new_n284_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n620_), .A2(new_n331_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n596_), .A2(new_n397_), .A3(new_n597_), .A4(new_n621_), .ZN(new_n622_));
  NAND4_X1  g421(.A1(new_n610_), .A2(new_n621_), .A3(new_n613_), .A4(new_n614_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT39), .ZN(new_n624_));
  AND3_X1   g423(.A1(new_n623_), .A2(new_n624_), .A3(G8gat), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n623_), .B2(G8gat), .ZN(new_n626_));
  OAI21_X1  g425(.A(new_n622_), .B1(new_n625_), .B2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n627_), .A2(KEYINPUT40), .ZN(new_n628_));
  XNOR2_X1  g427(.A(KEYINPUT103), .B(KEYINPUT104), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT40), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n622_), .B(new_n630_), .C1(new_n625_), .C2(new_n626_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n628_), .A2(new_n629_), .A3(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n629_), .B1(new_n628_), .B2(new_n631_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1325gat));
  OAI21_X1  g433(.A(G15gat), .B1(new_n616_), .B2(new_n379_), .ZN(new_n635_));
  OR2_X1    g434(.A1(new_n635_), .A2(KEYINPUT105), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(KEYINPUT105), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT41), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n636_), .A2(KEYINPUT41), .A3(new_n637_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n598_), .A2(new_n339_), .A3(new_n343_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n640_), .A2(new_n641_), .A3(new_n642_), .ZN(G1326gat));
  INV_X1    g442(.A(G22gat), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n378_), .A2(KEYINPUT106), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n378_), .A2(KEYINPUT106), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n598_), .A2(new_n644_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n647_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G22gat), .B1(new_n616_), .B2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n650_), .A2(KEYINPUT42), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(KEYINPUT42), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n648_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT107), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT107), .B(new_n648_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1327gat));
  NAND2_X1  g456(.A1(new_n609_), .A2(new_n465_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n594_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n422_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G29gat), .B1(new_n660_), .B2(new_n328_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT108), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n558_), .A2(new_n562_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n663_), .B1(new_n376_), .B2(new_n393_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT43), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n662_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n666_));
  OAI211_X1 g465(.A(KEYINPUT108), .B(KEYINPUT43), .C1(new_n605_), .C2(new_n663_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n663_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n665_), .B(new_n668_), .C1(new_n603_), .C2(new_n604_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n666_), .A2(new_n667_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n421_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n659_), .A2(new_n671_), .A3(new_n611_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n670_), .A2(KEYINPUT44), .A3(new_n672_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n673_), .A2(G29gat), .A3(new_n328_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n670_), .A2(new_n672_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n661_), .B1(new_n674_), .B2(new_n678_), .ZN(G1328gat));
  INV_X1    g478(.A(new_n672_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n669_), .ZN(new_n681_));
  OAI21_X1  g480(.A(KEYINPUT43), .B1(new_n605_), .B2(new_n663_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(new_n662_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n680_), .B1(new_n683_), .B2(new_n667_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n673_), .B(new_n621_), .C1(new_n684_), .C2(new_n676_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n685_), .A2(G36gat), .ZN(new_n686_));
  INV_X1    g485(.A(G36gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n660_), .A2(new_n687_), .A3(new_n621_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT45), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT110), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n691_), .A2(KEYINPUT46), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n690_), .A2(new_n692_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n686_), .B(new_n689_), .C1(new_n691_), .C2(KEYINPUT46), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1329gat));
  AOI21_X1  g494(.A(G43gat), .B1(new_n660_), .B2(new_n343_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT111), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n678_), .A2(G43gat), .A3(new_n343_), .A4(new_n673_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(KEYINPUT47), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT47), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n697_), .A2(new_n698_), .A3(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n700_), .A2(new_n702_), .ZN(G1330gat));
  INV_X1    g502(.A(G50gat), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n678_), .A2(new_n377_), .A3(new_n673_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(KEYINPUT112), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n706_), .B1(KEYINPUT112), .B2(new_n705_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n660_), .A2(new_n704_), .A3(new_n647_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1331gat));
  NAND2_X1  g508(.A1(new_n394_), .A2(new_n671_), .ZN(new_n710_));
  NOR4_X1   g509(.A1(new_n710_), .A2(new_n594_), .A3(new_n465_), .A4(new_n668_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(new_n437_), .A3(new_n328_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n610_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n659_), .A2(new_n671_), .A3(new_n611_), .ZN(new_n714_));
  NOR3_X1   g513(.A1(new_n713_), .A2(new_n329_), .A3(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n712_), .B1(new_n715_), .B2(new_n437_), .ZN(G1332gat));
  NOR2_X1   g515(.A1(new_n713_), .A2(new_n714_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n435_), .B1(new_n717_), .B2(new_n621_), .ZN(new_n718_));
  XOR2_X1   g517(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n711_), .A2(new_n435_), .A3(new_n621_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1333gat));
  INV_X1    g521(.A(G71gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n717_), .B2(new_n343_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT49), .Z(new_n725_));
  NAND3_X1  g524(.A1(new_n711_), .A2(new_n723_), .A3(new_n343_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1334gat));
  INV_X1    g526(.A(G78gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n717_), .B2(new_n647_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT50), .Z(new_n730_));
  NAND3_X1  g529(.A1(new_n711_), .A2(new_n728_), .A3(new_n647_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1335gat));
  NOR3_X1   g531(.A1(new_n710_), .A2(new_n658_), .A3(new_n594_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(new_n328_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n659_), .A2(new_n671_), .A3(new_n465_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n670_), .A2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n328_), .A2(G85gat), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT114), .Z(new_n739_));
  OAI22_X1  g538(.A1(G85gat), .A2(new_n734_), .B1(new_n737_), .B2(new_n739_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT115), .Z(G1336gat));
  INV_X1    g540(.A(new_n621_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G92gat), .B1(new_n737_), .B2(new_n742_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n733_), .A2(new_n488_), .A3(new_n621_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1337gat));
  OAI21_X1  g544(.A(G99gat), .B1(new_n737_), .B2(new_n379_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT116), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  OAI211_X1 g547(.A(KEYINPUT116), .B(G99gat), .C1(new_n737_), .C2(new_n379_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT117), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n343_), .A2(new_n502_), .A3(new_n503_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n750_), .B1(new_n733_), .B2(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n749_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(KEYINPUT51), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n748_), .A2(new_n755_), .A3(new_n749_), .A4(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1338gat));
  NAND3_X1  g556(.A1(new_n733_), .A2(new_n468_), .A3(new_n377_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n670_), .A2(new_n377_), .A3(new_n736_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n759_), .A2(new_n760_), .A3(G106gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n759_), .B2(G106gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n758_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT53), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n758_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n764_), .A2(new_n766_), .ZN(G1339gat));
  NAND2_X1  g566(.A1(new_n421_), .A2(new_n590_), .ZN(new_n768_));
  AND4_X1   g567(.A1(new_n570_), .A2(new_n565_), .A3(new_n572_), .A4(new_n574_), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n565_), .A2(new_n570_), .A3(new_n578_), .A4(new_n572_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n769_), .A2(KEYINPUT55), .B1(new_n573_), .B2(new_n770_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n577_), .A2(new_n772_), .A3(new_n583_), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n771_), .A2(new_n773_), .A3(KEYINPUT119), .ZN(new_n774_));
  AOI21_X1  g573(.A(KEYINPUT119), .B1(new_n771_), .B2(new_n773_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n589_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT56), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(KEYINPUT56), .B(new_n589_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n768_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n417_), .A2(new_n420_), .ZN(new_n781_));
  AND2_X1   g580(.A1(new_n405_), .A2(new_n406_), .ZN(new_n782_));
  OR2_X1    g581(.A1(new_n782_), .A2(new_n420_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n415_), .A2(new_n406_), .ZN(new_n784_));
  AOI22_X1  g583(.A1(new_n783_), .A2(KEYINPUT120), .B1(new_n412_), .B2(new_n784_), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(KEYINPUT120), .B2(new_n783_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n781_), .A2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n591_), .B2(new_n590_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n608_), .B1(new_n780_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT57), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n590_), .A2(new_n781_), .A3(new_n786_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT119), .ZN(new_n793_));
  AND3_X1   g592(.A1(new_n577_), .A2(new_n772_), .A3(new_n583_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n770_), .A2(new_n573_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n772_), .B2(new_n575_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n793_), .B1(new_n794_), .B2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n771_), .A2(new_n773_), .A3(KEYINPUT119), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(KEYINPUT56), .B1(new_n799_), .B2(new_n589_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n589_), .ZN(new_n801_));
  AOI211_X1 g600(.A(new_n777_), .B(new_n801_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n792_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT58), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  OAI211_X1 g604(.A(KEYINPUT58), .B(new_n792_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n805_), .A2(new_n668_), .A3(new_n806_), .ZN(new_n807_));
  OAI211_X1 g606(.A(new_n608_), .B(KEYINPUT57), .C1(new_n780_), .C2(new_n788_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n791_), .A2(new_n807_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n465_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n663_), .A2(new_n594_), .A3(new_n671_), .A4(new_n611_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT118), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n563_), .A2(KEYINPUT118), .A3(new_n671_), .A4(new_n594_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(KEYINPUT54), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT54), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n811_), .A2(new_n812_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n810_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT122), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT59), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n621_), .A2(new_n329_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n824_), .A2(new_n374_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n820_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n822_), .A2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n820_), .B(new_n825_), .C1(new_n821_), .C2(KEYINPUT59), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(G113gat), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT123), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n830_), .B1(new_n421_), .B2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n831_), .B2(new_n830_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT121), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n826_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n820_), .A2(KEYINPUT121), .A3(new_n825_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(new_n421_), .A3(new_n836_), .ZN(new_n837_));
  AOI22_X1  g636(.A1(new_n829_), .A2(new_n833_), .B1(new_n837_), .B2(new_n830_), .ZN(G1340gat));
  AOI21_X1  g637(.A(new_n594_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n839_));
  INV_X1    g638(.A(G120gat), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n835_), .A2(new_n836_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n594_), .B2(KEYINPUT60), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(KEYINPUT60), .B2(new_n840_), .ZN(new_n843_));
  OAI22_X1  g642(.A1(new_n839_), .A2(new_n840_), .B1(new_n841_), .B2(new_n843_), .ZN(G1341gat));
  AOI21_X1  g643(.A(new_n465_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n845_));
  INV_X1    g644(.A(G127gat), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n611_), .A2(new_n846_), .ZN(new_n847_));
  OAI22_X1  g646(.A1(new_n845_), .A2(new_n846_), .B1(new_n841_), .B2(new_n847_), .ZN(G1342gat));
  AOI21_X1  g647(.A(new_n663_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n849_));
  INV_X1    g648(.A(G134gat), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n609_), .A2(new_n850_), .ZN(new_n851_));
  OAI22_X1  g650(.A1(new_n849_), .A2(new_n850_), .B1(new_n841_), .B2(new_n851_), .ZN(G1343gat));
  AOI21_X1  g651(.A(new_n818_), .B1(new_n809_), .B2(new_n465_), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n853_), .A2(new_n602_), .A3(new_n824_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n421_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g655(.A1(new_n854_), .A2(new_n659_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g657(.A1(new_n854_), .A2(new_n611_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT61), .B(G155gat), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1346gat));
  INV_X1    g660(.A(G162gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n854_), .A2(new_n862_), .A3(new_n609_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n854_), .A2(new_n668_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n864_), .B2(new_n862_), .ZN(G1347gat));
  NOR3_X1   g664(.A1(new_n742_), .A2(new_n379_), .A3(new_n328_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n421_), .ZN(new_n867_));
  XOR2_X1   g666(.A(new_n867_), .B(KEYINPUT124), .Z(new_n868_));
  NAND3_X1  g667(.A1(new_n820_), .A2(new_n868_), .A3(new_n649_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n869_), .A2(new_n870_), .A3(G169gat), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n869_), .B2(G169gat), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT125), .ZN(new_n874_));
  INV_X1    g673(.A(new_n866_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n875_), .A2(new_n647_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n820_), .A2(new_n874_), .A3(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n876_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT125), .B1(new_n853_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n877_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n421_), .A2(new_n229_), .ZN(new_n881_));
  OAI22_X1  g680(.A1(new_n872_), .A2(new_n873_), .B1(new_n880_), .B2(new_n881_), .ZN(G1348gat));
  NAND3_X1  g681(.A1(new_n877_), .A2(new_n879_), .A3(new_n659_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n853_), .A2(new_n377_), .ZN(new_n884_));
  NOR3_X1   g683(.A1(new_n875_), .A2(new_n215_), .A3(new_n594_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n883_), .A2(new_n215_), .B1(new_n884_), .B2(new_n885_), .ZN(G1349gat));
  NOR2_X1   g685(.A1(new_n465_), .A2(new_n220_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n877_), .A2(new_n879_), .A3(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT126), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n877_), .A2(new_n879_), .A3(KEYINPUT126), .A4(new_n887_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n884_), .A2(new_n611_), .A3(new_n866_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(new_n206_), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n890_), .A2(new_n891_), .A3(new_n893_), .ZN(G1350gat));
  OAI21_X1  g693(.A(G190gat), .B1(new_n880_), .B2(new_n663_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n609_), .A2(new_n221_), .ZN(new_n896_));
  OAI21_X1  g695(.A(new_n895_), .B1(new_n880_), .B2(new_n896_), .ZN(G1351gat));
  NOR2_X1   g696(.A1(new_n742_), .A2(new_n328_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n663_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n806_), .A2(new_n899_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n611_), .B1(new_n900_), .B2(new_n808_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n372_), .B(new_n898_), .C1(new_n901_), .C2(new_n818_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(KEYINPUT127), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT127), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n820_), .A2(new_n904_), .A3(new_n372_), .A4(new_n898_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n905_), .ZN(new_n906_));
  AOI21_X1  g705(.A(G197gat), .B1(new_n906_), .B2(new_n421_), .ZN(new_n907_));
  AOI211_X1 g706(.A(new_n236_), .B(new_n671_), .C1(new_n903_), .C2(new_n905_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1352gat));
  AOI21_X1  g708(.A(new_n602_), .B1(new_n810_), .B2(new_n819_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n904_), .B1(new_n910_), .B2(new_n898_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n898_), .ZN(new_n912_));
  NOR4_X1   g711(.A1(new_n853_), .A2(KEYINPUT127), .A3(new_n602_), .A4(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n659_), .B1(new_n911_), .B2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(G204gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n906_), .A2(new_n233_), .A3(new_n659_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1353gat));
  NOR2_X1   g716(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n465_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n906_), .B2(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n920_), .ZN(new_n922_));
  AOI211_X1 g721(.A(new_n918_), .B(new_n922_), .C1(new_n903_), .C2(new_n905_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1354gat));
  INV_X1    g723(.A(G218gat), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n906_), .A2(new_n925_), .A3(new_n609_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n663_), .B1(new_n903_), .B2(new_n905_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n925_), .B2(new_n927_), .ZN(G1355gat));
endmodule


