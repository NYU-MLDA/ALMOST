//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n710_, new_n711_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n752_, new_n753_, new_n755_,
    new_n756_, new_n757_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n870_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n926_, new_n927_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n956_, new_n957_, new_n958_,
    new_n959_;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G78gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G22gat), .B(G50gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT85), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n211_), .A2(KEYINPUT1), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n213_), .B1(new_n211_), .B2(KEYINPUT1), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n215_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n218_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n222_), .A2(KEYINPUT2), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n216_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n222_), .A2(KEYINPUT2), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n217_), .A2(KEYINPUT3), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n223_), .A2(new_n225_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT86), .ZN(new_n229_));
  INV_X1    g028(.A(new_n213_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n211_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n229_), .B1(new_n211_), .B2(new_n230_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n228_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n221_), .A2(new_n234_), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT28), .B1(new_n235_), .B2(KEYINPUT29), .ZN(new_n236_));
  AND4_X1   g035(.A1(new_n223_), .A2(new_n226_), .A3(new_n225_), .A4(new_n227_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n233_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n237_), .B1(new_n238_), .B2(new_n231_), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n219_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n240_));
  OAI21_X1  g039(.A(KEYINPUT29), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  XOR2_X1   g040(.A(G197gat), .B(G204gat), .Z(new_n242_));
  OR2_X1    g041(.A1(new_n242_), .A2(KEYINPUT21), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(KEYINPUT21), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G211gat), .B(G218gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n244_), .A2(new_n245_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n241_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT28), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT29), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n234_), .A2(new_n221_), .A3(new_n250_), .A4(new_n251_), .ZN(new_n252_));
  AND3_X1   g051(.A1(new_n236_), .A2(new_n249_), .A3(new_n252_), .ZN(new_n253_));
  AOI21_X1  g052(.A(new_n249_), .B1(new_n236_), .B2(new_n252_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n209_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n236_), .A2(new_n252_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n249_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n236_), .A2(new_n249_), .A3(new_n252_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(new_n259_), .A3(new_n208_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n255_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G227gat), .A2(G233gat), .ZN(new_n263_));
  INV_X1    g062(.A(G15gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT30), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT31), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G71gat), .B(G99gat), .ZN(new_n269_));
  INV_X1    g068(.A(G43gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(G169gat), .ZN(new_n272_));
  INV_X1    g071(.A(G176gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G169gat), .A2(G176gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(KEYINPUT24), .A3(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT80), .ZN(new_n277_));
  INV_X1    g076(.A(G183gat), .ZN(new_n278_));
  INV_X1    g077(.A(G190gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(KEYINPUT23), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT23), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n281_), .A2(G183gat), .A3(G190gat), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n280_), .A2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT25), .B(G183gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(G190gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n274_), .A2(KEYINPUT24), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n277_), .A2(new_n283_), .A3(new_n288_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n275_), .ZN(new_n290_));
  OR2_X1    g089(.A1(new_n272_), .A2(KEYINPUT81), .ZN(new_n291_));
  AOI21_X1  g090(.A(G176gat), .B1(new_n291_), .B2(KEYINPUT22), .ZN(new_n292_));
  OR3_X1    g091(.A1(new_n272_), .A2(KEYINPUT81), .A3(KEYINPUT22), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n290_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n280_), .A2(KEYINPUT82), .A3(new_n282_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n295_), .B1(KEYINPUT82), .B2(new_n282_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(G183gat), .A2(G190gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n294_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT83), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n289_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n299_), .B1(new_n289_), .B2(new_n298_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n271_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n289_), .A2(new_n298_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n303_), .A2(KEYINPUT83), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n289_), .A2(new_n298_), .A3(new_n299_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n271_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n304_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n302_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G127gat), .B(G134gat), .Z(new_n309_));
  INV_X1    g108(.A(KEYINPUT84), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G127gat), .B(G134gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(KEYINPUT84), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G113gat), .B(G120gat), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n308_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n308_), .A2(new_n318_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n268_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n321_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n323_), .A2(new_n267_), .A3(new_n319_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G1gat), .B(G29gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(G85gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT0), .B(G57gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n311_), .A2(new_n313_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n314_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(new_n315_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n334_), .B1(new_n221_), .B2(new_n234_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n330_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n318_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n221_), .A2(new_n334_), .A3(new_n234_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(new_n339_), .A3(KEYINPUT4), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n337_), .A2(KEYINPUT91), .A3(new_n340_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n338_), .A2(new_n339_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n330_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  AOI21_X1  g143(.A(KEYINPUT91), .B1(new_n337_), .B2(new_n340_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n329_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT91), .ZN(new_n347_));
  INV_X1    g146(.A(new_n340_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n330_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n349_), .B1(new_n338_), .B2(KEYINPUT4), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n347_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n329_), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(new_n343_), .A4(new_n341_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n346_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n325_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT27), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G8gat), .B(G36gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT18), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G64gat), .B(G92gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  OAI21_X1  g159(.A(new_n248_), .B1(new_n300_), .B2(new_n301_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT90), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OAI211_X1 g162(.A(KEYINPUT90), .B(new_n248_), .C1(new_n300_), .C2(new_n301_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G226gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT19), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n283_), .B1(G183gat), .B2(G190gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT22), .B(G169gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n273_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT88), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n275_), .B(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT89), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n371_), .A2(new_n373_), .A3(new_n374_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n369_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n296_), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n286_), .A2(new_n287_), .A3(new_n276_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT87), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n286_), .A2(new_n287_), .A3(new_n276_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT87), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n381_), .A2(new_n296_), .A3(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n377_), .B1(new_n380_), .B2(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(KEYINPUT20), .B(new_n368_), .C1(new_n384_), .C2(new_n248_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n365_), .A2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT20), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n384_), .B2(new_n248_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n248_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n304_), .A2(new_n305_), .A3(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n368_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n360_), .B1(new_n387_), .B2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n385_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n360_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n395_), .A2(new_n396_), .A3(new_n392_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n356_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n389_), .A2(new_n391_), .ZN(new_n399_));
  OAI21_X1  g198(.A(KEYINPUT95), .B1(new_n399_), .B2(new_n367_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT95), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n389_), .A2(new_n391_), .A3(new_n401_), .A4(new_n368_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n400_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT93), .B(KEYINPUT20), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n377_), .B1(new_n296_), .B2(new_n381_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n405_), .A2(KEYINPUT94), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n248_), .B1(new_n405_), .B2(KEYINPUT94), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n404_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n368_), .B1(new_n365_), .B2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n396_), .B1(new_n403_), .B2(new_n409_), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n392_), .B1(new_n365_), .B2(new_n386_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n356_), .B1(new_n411_), .B2(new_n360_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  AND4_X1   g212(.A1(new_n262_), .A2(new_n355_), .A3(new_n398_), .A4(new_n413_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n352_), .A2(KEYINPUT33), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n351_), .A2(new_n343_), .A3(new_n341_), .A4(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n352_), .B1(new_n342_), .B2(new_n349_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n330_), .B1(new_n338_), .B2(KEYINPUT4), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n417_), .B1(new_n348_), .B2(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(new_n397_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n396_), .B1(new_n395_), .B2(new_n392_), .ZN(new_n422_));
  XOR2_X1   g221(.A(KEYINPUT92), .B(KEYINPUT33), .Z(new_n423_));
  NAND2_X1  g222(.A1(new_n353_), .A2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n420_), .A2(new_n421_), .A3(new_n422_), .A4(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n360_), .A2(KEYINPUT32), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n427_), .B1(new_n403_), .B2(new_n409_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n411_), .A2(new_n426_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(new_n354_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n262_), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n261_), .A2(new_n346_), .A3(new_n353_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n413_), .A2(new_n398_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n432_), .A2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n414_), .B1(new_n435_), .B2(new_n325_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G113gat), .B(G141gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G169gat), .B(G197gat), .ZN(new_n438_));
  XOR2_X1   g237(.A(new_n437_), .B(new_n438_), .Z(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G43gat), .B(G50gat), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(G36gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(G29gat), .ZN(new_n444_));
  INV_X1    g243(.A(G29gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n445_), .A2(G36gat), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n444_), .A2(new_n446_), .A3(KEYINPUT71), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT71), .B1(new_n444_), .B2(new_n446_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n442_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n444_), .A2(new_n446_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT71), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(new_n447_), .A3(new_n441_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n450_), .A2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n450_), .A2(new_n454_), .A3(new_n456_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G15gat), .B(G22gat), .ZN(new_n461_));
  INV_X1    g260(.A(G1gat), .ZN(new_n462_));
  INV_X1    g261(.A(G8gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G1gat), .B(G8gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n460_), .A2(new_n467_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n455_), .A2(new_n467_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G229gat), .A2(G233gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n468_), .A2(new_n469_), .A3(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(new_n467_), .B(new_n455_), .Z(new_n473_));
  NOR2_X1   g272(.A1(new_n473_), .A2(new_n470_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n440_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  OAI211_X1 g274(.A(new_n471_), .B(new_n439_), .C1(new_n473_), .C2(new_n470_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n475_), .A2(KEYINPUT79), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT79), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n478_), .B(new_n440_), .C1(new_n472_), .C2(new_n474_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(G85gat), .A2(G92gat), .ZN(new_n481_));
  NOR2_X1   g280(.A1(G85gat), .A2(G92gat), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G99gat), .A2(G106gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(KEYINPUT6), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(G99gat), .A3(G106gat), .ZN(new_n487_));
  AOI22_X1  g286(.A1(new_n483_), .A2(KEYINPUT9), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT65), .B1(new_n491_), .B2(G106gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT66), .B(G92gat), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT9), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n493_), .A2(new_n494_), .A3(G85gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT65), .ZN(new_n496_));
  NAND4_X1  g295(.A1(new_n489_), .A2(new_n496_), .A3(new_n205_), .A4(new_n490_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n488_), .A2(new_n492_), .A3(new_n495_), .A4(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G85gat), .B(G92gat), .ZN(new_n499_));
  OAI21_X1  g298(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n485_), .A2(new_n487_), .ZN(new_n504_));
  AOI211_X1 g303(.A(KEYINPUT8), .B(new_n499_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT8), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n507_));
  INV_X1    g306(.A(G99gat), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n508_), .A3(new_n205_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n486_), .B1(G99gat), .B2(G106gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n484_), .A2(KEYINPUT6), .ZN(new_n511_));
  OAI211_X1 g310(.A(new_n500_), .B(new_n509_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n506_), .B1(new_n512_), .B2(new_n483_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n498_), .B1(new_n505_), .B2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n514_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n510_), .A2(new_n511_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n509_), .A2(new_n500_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n483_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(KEYINPUT8), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n512_), .A2(new_n506_), .A3(new_n483_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n521_), .A2(new_n498_), .A3(new_n455_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n515_), .A2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT73), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT35), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n515_), .A2(new_n525_), .A3(new_n522_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G232gat), .A2(G233gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n526_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT73), .ZN(new_n531_));
  AOI211_X1 g330(.A(new_n531_), .B(new_n529_), .C1(new_n515_), .C2(new_n522_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n530_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G190gat), .B(G218gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT74), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G134gat), .B(G162gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n534_), .A2(KEYINPUT36), .A3(new_n538_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(KEYINPUT36), .ZN(new_n540_));
  INV_X1    g339(.A(new_n529_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n523_), .B2(KEYINPUT73), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n532_), .B1(new_n542_), .B2(new_n526_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n540_), .B1(new_n543_), .B2(KEYINPUT75), .ZN(new_n544_));
  AND4_X1   g343(.A1(KEYINPUT75), .A2(new_n530_), .A3(new_n533_), .A4(new_n540_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n539_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT37), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n548_), .B(new_n539_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G231gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n467_), .B(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(G71gat), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(G78gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n203_), .A2(G71gat), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(KEYINPUT11), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT67), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n559_), .B1(new_n557_), .B2(KEYINPUT11), .ZN(new_n560_));
  INV_X1    g359(.A(G64gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(G57gat), .ZN(new_n562_));
  INV_X1    g361(.A(G57gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(G64gat), .ZN(new_n564_));
  AND4_X1   g363(.A1(new_n559_), .A2(new_n562_), .A3(new_n564_), .A4(KEYINPUT11), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n558_), .B1(new_n560_), .B2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n562_), .A2(new_n564_), .A3(KEYINPUT11), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT67), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n562_), .A2(new_n564_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT11), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n562_), .A2(new_n564_), .A3(new_n559_), .A4(KEYINPUT11), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n568_), .A2(new_n571_), .A3(new_n556_), .A4(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n566_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n552_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G127gat), .B(G155gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT16), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G183gat), .B(G211gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  XNOR2_X1  g378(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n575_), .A2(new_n581_), .ZN(new_n582_));
  XOR2_X1   g381(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n584_), .B(KEYINPUT77), .Z(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n575_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n550_), .A2(new_n587_), .ZN(new_n588_));
  AND2_X1   g387(.A1(new_n566_), .A2(new_n573_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n521_), .A3(new_n498_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n514_), .A2(new_n574_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n590_), .A2(new_n591_), .A3(KEYINPUT12), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n514_), .A2(new_n593_), .A3(new_n574_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G230gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT64), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT68), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n590_), .A2(new_n591_), .A3(new_n598_), .ZN(new_n599_));
  AOI22_X1  g398(.A1(new_n521_), .A2(new_n498_), .B1(new_n573_), .B2(new_n566_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n597_), .B1(new_n600_), .B2(KEYINPUT68), .ZN(new_n601_));
  AOI22_X1  g400(.A1(new_n595_), .A2(new_n597_), .B1(new_n599_), .B2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G176gat), .B(G204gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT70), .ZN(new_n604_));
  XOR2_X1   g403(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(G120gat), .B(G148gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n606_), .B(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n602_), .B(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(KEYINPUT13), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n609_), .A2(KEYINPUT13), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n588_), .A2(new_n614_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n436_), .A2(new_n480_), .A3(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n462_), .A3(new_n354_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT38), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT97), .ZN(new_n619_));
  OAI21_X1  g418(.A(new_n619_), .B1(new_n436_), .B2(new_n546_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n261_), .B1(new_n425_), .B2(new_n430_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n413_), .A2(new_n398_), .A3(new_n433_), .ZN(new_n622_));
  OAI21_X1  g421(.A(new_n325_), .B1(new_n621_), .B2(new_n622_), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n413_), .A2(new_n398_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n624_), .A2(new_n262_), .A3(new_n355_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n546_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(KEYINPUT97), .A3(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n620_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n480_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n587_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n614_), .A2(new_n630_), .A3(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT96), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n629_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n354_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G1gat), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n618_), .A2(new_n636_), .ZN(G1324gat));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638_));
  INV_X1    g437(.A(new_n624_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n629_), .A2(KEYINPUT99), .A3(new_n639_), .A4(new_n633_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(G8gat), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n628_), .ZN(new_n643_));
  AOI21_X1  g442(.A(KEYINPUT97), .B1(new_n626_), .B2(new_n627_), .ZN(new_n644_));
  OAI211_X1 g443(.A(new_n639_), .B(new_n633_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT99), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT39), .B1(new_n642_), .B2(new_n647_), .ZN(new_n648_));
  NAND4_X1  g447(.A1(new_n647_), .A2(new_n640_), .A3(KEYINPUT39), .A4(G8gat), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n616_), .A2(new_n463_), .A3(new_n639_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT98), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n638_), .B1(new_n648_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT39), .ZN(new_n654_));
  INV_X1    g453(.A(new_n647_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(new_n655_), .B2(new_n641_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n656_), .A2(KEYINPUT40), .A3(new_n649_), .A4(new_n651_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n653_), .A2(new_n657_), .ZN(G1325gat));
  OAI21_X1  g457(.A(G15gat), .B1(new_n634_), .B2(new_n325_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT100), .B(KEYINPUT41), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(new_n660_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n325_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n616_), .A2(new_n264_), .A3(new_n663_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n661_), .A2(new_n662_), .A3(new_n664_), .ZN(G1326gat));
  INV_X1    g464(.A(G22gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n616_), .A2(new_n666_), .A3(new_n261_), .ZN(new_n667_));
  OAI21_X1  g466(.A(G22gat), .B1(new_n634_), .B2(new_n262_), .ZN(new_n668_));
  XNOR2_X1  g467(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n668_), .A2(new_n669_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n667_), .B1(new_n670_), .B2(new_n671_), .ZN(G1327gat));
  NOR3_X1   g471(.A1(new_n613_), .A2(new_n627_), .A3(new_n631_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n626_), .A2(new_n630_), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT104), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n626_), .A2(KEYINPUT104), .A3(new_n630_), .A4(new_n673_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(G29gat), .B1(new_n678_), .B2(new_n354_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n613_), .A2(new_n480_), .A3(new_n631_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT102), .B(KEYINPUT43), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n626_), .B2(new_n550_), .ZN(new_n683_));
  INV_X1    g482(.A(new_n550_), .ZN(new_n684_));
  AOI211_X1 g483(.A(KEYINPUT43), .B(new_n684_), .C1(new_n623_), .C2(new_n625_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n680_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT103), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n686_), .A2(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n688_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n635_), .A2(new_n445_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n679_), .B1(new_n691_), .B2(new_n692_), .ZN(G1328gat));
  NAND4_X1  g492(.A1(new_n676_), .A2(new_n443_), .A3(new_n639_), .A4(new_n677_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n694_), .B(KEYINPUT45), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n624_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(new_n443_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  OAI211_X1 g498(.A(KEYINPUT46), .B(new_n695_), .C1(new_n696_), .C2(new_n443_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(G1329gat));
  NAND3_X1  g500(.A1(new_n678_), .A2(new_n270_), .A3(new_n663_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n325_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(new_n270_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n704_), .A2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n702_), .B(new_n705_), .C1(new_n703_), .C2(new_n270_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1330gat));
  AOI21_X1  g508(.A(G50gat), .B1(new_n678_), .B2(new_n261_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n261_), .A2(G50gat), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n710_), .B1(new_n691_), .B2(new_n711_), .ZN(G1331gat));
  AOI211_X1 g511(.A(new_n614_), .B(new_n630_), .C1(new_n623_), .C2(new_n625_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n588_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n714_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n563_), .A3(new_n354_), .ZN(new_n716_));
  AND4_X1   g515(.A1(new_n629_), .A2(new_n613_), .A3(new_n480_), .A4(new_n631_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n717_), .A2(new_n354_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n716_), .B1(new_n718_), .B2(new_n563_), .ZN(G1332gat));
  NAND3_X1  g518(.A1(new_n715_), .A2(new_n561_), .A3(new_n639_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT48), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n717_), .A2(new_n639_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(G64gat), .ZN(new_n723_));
  AOI211_X1 g522(.A(KEYINPUT48), .B(new_n561_), .C1(new_n717_), .C2(new_n639_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n720_), .B1(new_n723_), .B2(new_n724_), .ZN(G1333gat));
  INV_X1    g524(.A(KEYINPUT49), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n717_), .A2(new_n663_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(G71gat), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT49), .B(new_n553_), .C1(new_n717_), .C2(new_n663_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n325_), .A2(G71gat), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT106), .ZN(new_n731_));
  OAI22_X1  g530(.A1(new_n728_), .A2(new_n729_), .B1(new_n714_), .B2(new_n731_), .ZN(G1334gat));
  NAND3_X1  g531(.A1(new_n715_), .A2(new_n203_), .A3(new_n261_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n717_), .A2(new_n261_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n734_), .B1(new_n735_), .B2(G78gat), .ZN(new_n736_));
  AOI211_X1 g535(.A(KEYINPUT50), .B(new_n203_), .C1(new_n717_), .C2(new_n261_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n733_), .B1(new_n736_), .B2(new_n737_), .ZN(G1335gat));
  NOR2_X1   g537(.A1(new_n627_), .A2(new_n631_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n713_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(G85gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(new_n354_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n613_), .A2(new_n480_), .A3(new_n587_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n683_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n663_), .B1(new_n432_), .B2(new_n434_), .ZN(new_n747_));
  OAI211_X1 g546(.A(new_n746_), .B(new_n550_), .C1(new_n747_), .C2(new_n414_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n744_), .B1(new_n745_), .B2(new_n748_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n749_), .A2(new_n354_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n743_), .B1(new_n750_), .B2(new_n742_), .ZN(G1336gat));
  AOI21_X1  g550(.A(G92gat), .B1(new_n741_), .B2(new_n639_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n639_), .A2(new_n493_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n749_), .B2(new_n753_), .ZN(G1337gat));
  NOR3_X1   g553(.A1(new_n740_), .A2(new_n325_), .A3(new_n491_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n749_), .A2(new_n663_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n756_), .B2(G99gat), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g557(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n759_));
  INV_X1    g558(.A(new_n744_), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n261_), .B(new_n760_), .C1(new_n683_), .C2(new_n685_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT108), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n684_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n748_), .B1(new_n764_), .B2(new_n682_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n765_), .A2(KEYINPUT108), .A3(new_n261_), .A4(new_n760_), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n763_), .A2(KEYINPUT52), .A3(G106gat), .A4(new_n766_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n713_), .A2(new_n205_), .A3(new_n261_), .A4(new_n739_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n768_), .B(new_n769_), .ZN(new_n770_));
  AND2_X1   g569(.A1(new_n767_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n763_), .A2(G106gat), .A3(new_n766_), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n759_), .B1(new_n771_), .B2(new_n774_), .ZN(new_n775_));
  AND4_X1   g574(.A1(new_n774_), .A2(new_n767_), .A3(new_n770_), .A4(new_n759_), .ZN(new_n776_));
  NOR2_X1   g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1339gat));
  INV_X1    g576(.A(G113gat), .ZN(new_n778_));
  INV_X1    g577(.A(new_n470_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n440_), .B1(new_n473_), .B2(new_n779_), .ZN(new_n780_));
  OR2_X1    g579(.A1(new_n780_), .A2(KEYINPUT111), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n468_), .A2(new_n469_), .A3(new_n779_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n780_), .A2(KEYINPUT111), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n781_), .A2(new_n782_), .A3(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n602_), .A2(new_n608_), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(new_n785_), .A3(new_n476_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT112), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n597_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n592_), .A2(new_n790_), .A3(new_n594_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT55), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n595_), .A2(new_n597_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT12), .B1(new_n514_), .B2(new_n574_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n795_), .A2(new_n600_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n594_), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT55), .B(new_n597_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n595_), .A2(KEYINPUT110), .A3(KEYINPUT55), .A4(new_n597_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n794_), .A2(new_n800_), .A3(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n608_), .ZN(new_n803_));
  AND3_X1   g602(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(KEYINPUT56), .B1(new_n802_), .B2(new_n803_), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n786_), .B(new_n789_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n550_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n802_), .A2(new_n803_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT56), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n802_), .A2(KEYINPUT56), .A3(new_n803_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n789_), .B1(new_n812_), .B2(new_n786_), .ZN(new_n813_));
  OAI21_X1  g612(.A(KEYINPUT113), .B1(new_n807_), .B2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n786_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n815_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT113), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n816_), .A2(new_n817_), .A3(new_n550_), .A4(new_n806_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n814_), .A2(new_n818_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n477_), .A2(new_n785_), .A3(new_n479_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n609_), .A2(new_n476_), .A3(new_n784_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT57), .B1(new_n823_), .B2(new_n627_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  AOI211_X1 g624(.A(new_n825_), .B(new_n546_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n824_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n819_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n819_), .A2(new_n827_), .A3(KEYINPUT114), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n830_), .A2(new_n587_), .A3(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(KEYINPUT54), .B1(new_n615_), .B2(new_n630_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n588_), .A2(new_n834_), .A3(new_n614_), .A4(new_n480_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n832_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n639_), .A2(new_n261_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n838_), .A2(new_n354_), .A3(new_n663_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n837_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n778_), .B1(new_n841_), .B2(new_n480_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(KEYINPUT115), .B(new_n778_), .C1(new_n841_), .C2(new_n480_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n836_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n816_), .A2(new_n550_), .A3(new_n806_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n631_), .B1(new_n827_), .B2(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n846_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n840_), .A2(new_n850_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n849_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n841_), .B2(KEYINPUT59), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n480_), .A2(new_n778_), .ZN(new_n855_));
  AOI22_X1  g654(.A1(new_n844_), .A2(new_n845_), .B1(new_n854_), .B2(new_n855_), .ZN(G1340gat));
  AOI21_X1  g655(.A(new_n839_), .B1(new_n832_), .B2(new_n836_), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT116), .B(G120gat), .Z(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n613_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n858_), .A2(KEYINPUT60), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(KEYINPUT117), .B2(new_n863_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n857_), .B(new_n864_), .C1(KEYINPUT117), .C2(new_n862_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n613_), .B(new_n852_), .C1(new_n857_), .C2(new_n850_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n865_), .B1(new_n867_), .B2(new_n858_), .ZN(G1341gat));
  AOI21_X1  g667(.A(G127gat), .B1(new_n857_), .B2(new_n631_), .ZN(new_n869_));
  INV_X1    g668(.A(G127gat), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n631_), .B2(KEYINPUT118), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(KEYINPUT118), .B2(new_n870_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n869_), .B1(new_n854_), .B2(new_n872_), .ZN(G1342gat));
  INV_X1    g672(.A(G134gat), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n684_), .A2(new_n874_), .ZN(new_n875_));
  OAI211_X1 g674(.A(new_n852_), .B(new_n875_), .C1(new_n857_), .C2(new_n850_), .ZN(new_n876_));
  AND3_X1   g675(.A1(new_n819_), .A2(new_n827_), .A3(KEYINPUT114), .ZN(new_n877_));
  AOI21_X1  g676(.A(KEYINPUT114), .B1(new_n819_), .B2(new_n827_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n877_), .A2(new_n878_), .A3(new_n631_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n546_), .B(new_n840_), .C1(new_n879_), .C2(new_n846_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(new_n874_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n876_), .A2(new_n881_), .ZN(new_n882_));
  INV_X1    g681(.A(KEYINPUT119), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n876_), .A2(new_n881_), .A3(KEYINPUT119), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(G1343gat));
  NAND4_X1  g685(.A1(new_n624_), .A2(new_n354_), .A3(new_n261_), .A4(new_n325_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(KEYINPUT120), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n837_), .A2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n630_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n613_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g692(.A1(new_n837_), .A2(new_n888_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n587_), .ZN(new_n895_));
  XOR2_X1   g694(.A(KEYINPUT61), .B(G155gat), .Z(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1346gat));
  OR3_X1    g696(.A1(new_n894_), .A2(G162gat), .A3(new_n627_), .ZN(new_n898_));
  OAI21_X1  g697(.A(G162gat), .B1(new_n894_), .B2(new_n684_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1347gat));
  NOR3_X1   g699(.A1(new_n624_), .A2(new_n354_), .A3(new_n325_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n262_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n630_), .B(new_n903_), .C1(new_n846_), .C2(new_n848_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n905_), .A2(KEYINPUT121), .A3(new_n272_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT62), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT121), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n904_), .B2(G169gat), .ZN(new_n909_));
  OR3_X1    g708(.A1(new_n906_), .A2(new_n907_), .A3(new_n909_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n905_), .A2(new_n370_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n907_), .B1(new_n906_), .B2(new_n909_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n910_), .A2(new_n911_), .A3(new_n912_), .ZN(G1348gat));
  AOI21_X1  g712(.A(new_n631_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n846_), .B1(new_n914_), .B2(new_n831_), .ZN(new_n915_));
  OR3_X1    g714(.A1(new_n915_), .A2(KEYINPUT122), .A3(new_n261_), .ZN(new_n916_));
  OAI21_X1  g715(.A(KEYINPUT122), .B1(new_n915_), .B2(new_n261_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n614_), .A2(new_n273_), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n916_), .A2(new_n917_), .A3(new_n901_), .A4(new_n918_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n903_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n273_), .B1(new_n920_), .B2(new_n614_), .ZN(new_n921_));
  AND2_X1   g720(.A1(new_n919_), .A2(new_n921_), .ZN(G1349gat));
  NOR3_X1   g721(.A1(new_n920_), .A2(new_n284_), .A3(new_n587_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n916_), .A2(new_n917_), .A3(new_n631_), .A4(new_n901_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n923_), .B1(new_n924_), .B2(new_n278_), .ZN(G1350gat));
  OAI21_X1  g724(.A(G190gat), .B1(new_n920_), .B2(new_n684_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n546_), .A2(new_n285_), .ZN(new_n927_));
  OAI21_X1  g726(.A(new_n926_), .B1(new_n920_), .B2(new_n927_), .ZN(G1351gat));
  NAND2_X1  g727(.A1(new_n433_), .A2(new_n325_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  OR2_X1    g729(.A1(new_n930_), .A2(KEYINPUT123), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(KEYINPUT123), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n931_), .A2(new_n639_), .A3(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(KEYINPUT124), .B1(new_n915_), .B2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT124), .ZN(new_n935_));
  INV_X1    g734(.A(new_n933_), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n935_), .B(new_n936_), .C1(new_n879_), .C2(new_n846_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n934_), .A2(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(G197gat), .B1(new_n938_), .B2(new_n630_), .ZN(new_n939_));
  INV_X1    g738(.A(G197gat), .ZN(new_n940_));
  AOI211_X1 g739(.A(new_n940_), .B(new_n480_), .C1(new_n934_), .C2(new_n937_), .ZN(new_n941_));
  NOR2_X1   g740(.A1(new_n939_), .A2(new_n941_), .ZN(G1352gat));
  NAND2_X1  g741(.A1(new_n938_), .A2(new_n613_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(G204gat), .ZN(new_n944_));
  INV_X1    g743(.A(G204gat), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n938_), .A2(new_n945_), .A3(new_n613_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n944_), .A2(new_n946_), .ZN(G1353gat));
  AOI21_X1  g746(.A(new_n587_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n938_), .A2(new_n948_), .ZN(new_n949_));
  NOR2_X1   g748(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n950_));
  XNOR2_X1  g749(.A(new_n950_), .B(KEYINPUT125), .ZN(new_n951_));
  INV_X1    g750(.A(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n949_), .A2(new_n952_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n938_), .A2(new_n951_), .A3(new_n948_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(G1354gat));
  NAND2_X1  g754(.A1(new_n938_), .A2(new_n546_), .ZN(new_n956_));
  INV_X1    g755(.A(G218gat), .ZN(new_n957_));
  NAND2_X1  g756(.A1(new_n550_), .A2(G218gat), .ZN(new_n958_));
  XOR2_X1   g757(.A(new_n958_), .B(KEYINPUT126), .Z(new_n959_));
  AOI22_X1  g758(.A1(new_n956_), .A2(new_n957_), .B1(new_n938_), .B2(new_n959_), .ZN(G1355gat));
endmodule


