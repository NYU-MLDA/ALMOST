//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n602_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n876_;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n203_));
  XOR2_X1   g002(.A(G71gat), .B(G78gat), .Z(new_n204_));
  NOR2_X1   g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  AND2_X1   g004(.A1(new_n203_), .A2(new_n204_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n202_), .A2(KEYINPUT11), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(new_n205_), .B1(new_n206_), .B2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G85gat), .ZN(new_n210_));
  INV_X1    g009(.A(G92gat), .ZN(new_n211_));
  NOR3_X1   g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT9), .ZN(new_n212_));
  XOR2_X1   g011(.A(G85gat), .B(G92gat), .Z(new_n213_));
  AOI21_X1  g012(.A(new_n212_), .B1(new_n213_), .B2(KEYINPUT9), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT10), .B(G99gat), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n215_), .A2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n219_));
  NOR2_X1   g018(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n218_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(KEYINPUT64), .A2(KEYINPUT6), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n217_), .A3(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n214_), .A2(new_n216_), .A3(new_n221_), .A4(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT65), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n221_), .A2(new_n226_), .ZN(new_n229_));
  OR3_X1    g028(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  OAI211_X1 g031(.A(new_n228_), .B(new_n213_), .C1(new_n229_), .C2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT8), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n221_), .A2(new_n226_), .A3(new_n231_), .A4(new_n230_), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n228_), .B1(new_n235_), .B2(new_n213_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n227_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  AOI211_X1 g036(.A(new_n228_), .B(KEYINPUT8), .C1(new_n235_), .C2(new_n213_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n209_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(KEYINPUT66), .A2(KEYINPUT12), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G230gat), .A2(G233gat), .ZN(new_n245_));
  OR3_X1    g044(.A1(new_n237_), .A2(new_n238_), .A3(new_n209_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n239_), .A2(new_n240_), .A3(new_n242_), .ZN(new_n247_));
  NAND4_X1  g046(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .A4(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n239_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n245_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n248_), .A2(new_n251_), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G120gat), .B(G148gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT5), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G176gat), .B(G204gat), .ZN(new_n255_));
  XOR2_X1   g054(.A(new_n254_), .B(new_n255_), .Z(new_n256_));
  NAND2_X1  g055(.A1(new_n252_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n256_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n248_), .A2(new_n251_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n257_), .A2(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT13), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT13), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n257_), .A2(new_n262_), .A3(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G127gat), .B(G134gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G113gat), .B(G120gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G71gat), .B(G99gat), .ZN(new_n269_));
  INV_X1    g068(.A(G43gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G227gat), .A2(G233gat), .ZN(new_n272_));
  INV_X1    g071(.A(G15gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n271_), .B(new_n274_), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT23), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n277_), .A2(G183gat), .A3(G190gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(KEYINPUT82), .ZN(new_n279_));
  INV_X1    g078(.A(G183gat), .ZN(new_n280_));
  INV_X1    g079(.A(G190gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT23), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  OR2_X1    g082(.A1(G169gat), .A2(G176gat), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n283_), .B1(KEYINPUT24), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT83), .ZN(new_n286_));
  OR2_X1    g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n285_), .A2(new_n286_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT25), .B(G183gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OR2_X1    g090(.A1(new_n291_), .A2(KEYINPUT80), .ZN(new_n292_));
  NAND2_X1  g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n293_), .B(KEYINPUT81), .Z(new_n294_));
  NAND2_X1  g093(.A1(new_n284_), .A2(KEYINPUT24), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n294_), .A2(new_n296_), .B1(new_n291_), .B2(KEYINPUT80), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n287_), .A2(new_n288_), .A3(new_n292_), .A4(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n282_), .B(KEYINPUT84), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n278_), .B(KEYINPUT85), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  OAI21_X1  g100(.A(new_n301_), .B1(G183gat), .B2(G190gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(KEYINPUT22), .B(G169gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n294_), .B1(G176gat), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n302_), .A2(new_n306_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n298_), .A2(KEYINPUT30), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(KEYINPUT30), .B1(new_n298_), .B2(new_n307_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n276_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n298_), .A2(new_n307_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT30), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n298_), .A2(KEYINPUT30), .A3(new_n307_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n313_), .A2(new_n275_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT31), .ZN(new_n316_));
  AND3_X1   g115(.A1(new_n310_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n316_), .B1(new_n310_), .B2(new_n315_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n268_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n310_), .A2(new_n315_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(KEYINPUT31), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n310_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n322_), .A2(new_n267_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n320_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G141gat), .A2(G148gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT2), .ZN(new_n329_));
  OAI22_X1  g128(.A1(KEYINPUT86), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n330_));
  NAND2_X1  g129(.A1(KEYINPUT86), .A2(KEYINPUT3), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OR2_X1    g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(KEYINPUT86), .A3(KEYINPUT3), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n329_), .A2(new_n332_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(G155gat), .ZN(new_n336_));
  INV_X1    g135(.A(G162gat), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n336_), .A2(new_n337_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n335_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n339_), .A2(KEYINPUT1), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT1), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n338_), .B1(new_n343_), .B2(new_n340_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n328_), .B(new_n333_), .C1(new_n342_), .C2(new_n344_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n341_), .A2(new_n345_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(new_n346_), .A2(KEYINPUT4), .A3(new_n267_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n347_), .B(KEYINPUT97), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n346_), .B(new_n268_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT4), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n348_), .A2(G225gat), .A3(G233gat), .A4(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G1gat), .B(G29gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT0), .ZN(new_n355_));
  INV_X1    g154(.A(G57gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n355_), .B(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(new_n210_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n351_), .A2(new_n353_), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n359_), .B1(new_n351_), .B2(new_n353_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(G226gat), .A2(G233gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(KEYINPUT19), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G211gat), .B(G218gat), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT90), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT88), .B(G197gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(G204gat), .ZN(new_n368_));
  INV_X1    g167(.A(G197gat), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n368_), .B1(new_n369_), .B2(G204gat), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n366_), .A2(KEYINPUT21), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT91), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT89), .B1(new_n367_), .B2(G204gat), .ZN(new_n374_));
  INV_X1    g173(.A(G204gat), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n374_), .B1(G197gat), .B2(new_n375_), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n367_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT21), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n378_), .B(new_n364_), .C1(KEYINPUT21), .C2(new_n370_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n373_), .A2(new_n379_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n311_), .A2(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n373_), .A2(new_n379_), .ZN(new_n382_));
  AOI22_X1  g181(.A1(new_n279_), .A2(new_n282_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n383_));
  OR2_X1    g182(.A1(new_n383_), .A2(KEYINPUT95), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n305_), .B1(new_n383_), .B2(KEYINPUT95), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT94), .B(KEYINPUT24), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n386_), .A2(new_n293_), .A3(new_n284_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n387_), .B1(new_n284_), .B2(new_n386_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n388_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n290_), .B(KEYINPUT93), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n289_), .ZN(new_n391_));
  AOI22_X1  g190(.A1(new_n384_), .A2(new_n385_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT20), .B1(new_n382_), .B2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n363_), .B1(new_n381_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT20), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n395_), .B1(new_n311_), .B2(new_n380_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n363_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n382_), .A2(new_n392_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n396_), .A2(new_n397_), .A3(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n394_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G8gat), .B(G36gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n401_), .B(KEYINPUT18), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(KEYINPUT96), .ZN(new_n403_));
  XOR2_X1   g202(.A(G64gat), .B(G92gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(KEYINPUT32), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  OAI22_X1  g206(.A1(new_n360_), .A2(new_n361_), .B1(new_n400_), .B2(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n397_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n409_), .A2(KEYINPUT99), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n381_), .A2(new_n393_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n409_), .A2(KEYINPUT99), .B1(new_n412_), .B2(new_n397_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n406_), .B1(new_n411_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n360_), .A2(KEYINPUT33), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n351_), .A2(new_n353_), .A3(new_n359_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n416_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n348_), .A2(new_n352_), .A3(new_n350_), .ZN(new_n419_));
  XOR2_X1   g218(.A(new_n349_), .B(KEYINPUT98), .Z(new_n420_));
  OAI211_X1 g219(.A(new_n358_), .B(new_n419_), .C1(new_n420_), .C2(new_n352_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n415_), .A2(new_n418_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n405_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n400_), .A2(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n394_), .A2(new_n399_), .A3(new_n405_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  OAI22_X1  g225(.A1(new_n408_), .A2(new_n414_), .B1(new_n422_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT29), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n346_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT28), .ZN(new_n430_));
  XOR2_X1   g229(.A(G22gat), .B(G50gat), .Z(new_n431_));
  OR2_X1    g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n430_), .A2(new_n431_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT87), .ZN(new_n434_));
  AND3_X1   g233(.A1(new_n432_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n434_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n346_), .A2(new_n428_), .ZN(new_n437_));
  OAI211_X1 g236(.A(G228gat), .B(G233gat), .C1(new_n382_), .C2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G228gat), .A2(G233gat), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n380_), .B(new_n439_), .C1(new_n428_), .C2(new_n346_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G78gat), .B(G106gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n442_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n444_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n445_));
  OAI22_X1  g244(.A1(new_n435_), .A2(new_n436_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT92), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n445_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n432_), .A2(new_n433_), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n438_), .A2(new_n440_), .A3(KEYINPUT92), .A4(new_n444_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .A4(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n446_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n327_), .A2(new_n427_), .A3(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n412_), .A2(new_n397_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n311_), .A2(new_n380_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(new_n398_), .A3(KEYINPUT20), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(new_n363_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT99), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n456_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n423_), .B1(new_n461_), .B2(new_n410_), .ZN(new_n462_));
  AND2_X1   g261(.A1(new_n425_), .A2(KEYINPUT27), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT27), .ZN(new_n464_));
  AOI22_X1  g263(.A1(new_n462_), .A2(new_n463_), .B1(new_n426_), .B2(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n360_), .A2(new_n361_), .ZN(new_n466_));
  AND4_X1   g265(.A1(new_n324_), .A2(new_n319_), .A3(new_n452_), .A4(new_n446_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n324_), .A2(new_n319_), .B1(new_n446_), .B2(new_n452_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n465_), .B(new_n466_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n455_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT75), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G15gat), .B(G22gat), .ZN(new_n472_));
  INV_X1    g271(.A(G1gat), .ZN(new_n473_));
  INV_X1    g272(.A(G8gat), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT14), .B1(new_n473_), .B2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G1gat), .B(G8gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G29gat), .B(G36gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G43gat), .B(G50gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n471_), .B1(new_n478_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT76), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n485_), .B1(new_n478_), .B2(new_n482_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n478_), .A2(new_n482_), .A3(new_n485_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n484_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n488_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n483_), .B1(new_n490_), .B2(new_n486_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n489_), .A2(new_n491_), .A3(G229gat), .A4(G233gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n478_), .A2(new_n482_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n481_), .B(KEYINPUT15), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n494_), .B2(new_n478_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G229gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT77), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n495_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G113gat), .B(G141gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G169gat), .B(G197gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n499_), .B(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n492_), .A2(new_n498_), .A3(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT78), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n502_), .B1(new_n492_), .B2(new_n498_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n504_), .A2(new_n505_), .ZN(new_n508_));
  OAI21_X1  g307(.A(KEYINPUT79), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n505_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(KEYINPUT78), .A3(new_n503_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT79), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n506_), .ZN(new_n513_));
  AND4_X1   g312(.A1(new_n264_), .A2(new_n470_), .A3(new_n509_), .A4(new_n513_), .ZN(new_n514_));
  XOR2_X1   g313(.A(G190gat), .B(G218gat), .Z(new_n515_));
  XNOR2_X1  g314(.A(G134gat), .B(G162gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT36), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n518_), .B(KEYINPUT71), .Z(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT67), .B(KEYINPUT34), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G232gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT35), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  OR2_X1    g324(.A1(new_n234_), .A2(new_n236_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n238_), .ZN(new_n527_));
  NAND4_X1  g326(.A1(new_n526_), .A2(new_n481_), .A3(new_n527_), .A4(new_n227_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n523_), .A2(new_n524_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT69), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n525_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n494_), .B1(new_n237_), .B2(new_n238_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT68), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n528_), .A2(new_n529_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n532_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n532_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n537_));
  OAI211_X1 g336(.A(KEYINPUT72), .B(new_n520_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(new_n535_), .ZN(new_n539_));
  AOI211_X1 g338(.A(new_n524_), .B(new_n523_), .C1(new_n528_), .C2(KEYINPUT69), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n532_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n517_), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT70), .B(KEYINPUT36), .Z(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n542_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n538_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n519_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n548_), .A2(KEYINPUT72), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT37), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT73), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n518_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT37), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n552_), .A2(new_n553_), .A3(new_n546_), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n550_), .A2(new_n551_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n551_), .B1(new_n550_), .B2(new_n554_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G231gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n478_), .B(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(new_n209_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G127gat), .B(G155gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(G183gat), .B(G211gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(KEYINPUT17), .A3(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(new_n565_), .B(KEYINPUT17), .Z(new_n568_));
  OAI21_X1  g367(.A(new_n567_), .B1(new_n560_), .B2(new_n568_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n557_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n514_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n466_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n572_), .A2(new_n473_), .A3(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT38), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n552_), .A2(new_n546_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n577_), .B1(new_n455_), .B2(new_n469_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n569_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n507_), .A2(new_n508_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n264_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT100), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(G1gat), .B1(new_n584_), .B2(new_n466_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n575_), .A2(new_n585_), .ZN(G1324gat));
  INV_X1    g385(.A(new_n465_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n572_), .A2(new_n474_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT39), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n580_), .A2(new_n583_), .A3(new_n587_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n589_), .B1(new_n590_), .B2(G8gat), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT101), .ZN(new_n592_));
  AND2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n590_), .A2(new_n589_), .A3(G8gat), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n594_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n588_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g396(.A(G15gat), .B1(new_n584_), .B2(new_n327_), .ZN(new_n598_));
  XOR2_X1   g397(.A(KEYINPUT102), .B(KEYINPUT41), .Z(new_n599_));
  OR2_X1    g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n598_), .A2(new_n599_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n572_), .A2(new_n273_), .A3(new_n326_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n600_), .A2(new_n601_), .A3(new_n602_), .ZN(G1326gat));
  OAI21_X1  g402(.A(G22gat), .B1(new_n584_), .B2(new_n454_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT42), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n454_), .A2(G22gat), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n605_), .B1(new_n571_), .B2(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT103), .ZN(G1327gat));
  NOR2_X1   g407(.A1(new_n576_), .A2(new_n579_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n514_), .A2(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(G29gat), .B1(new_n610_), .B2(new_n573_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT106), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n583_), .A2(new_n569_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT104), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n557_), .A2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n536_), .A2(new_n537_), .ZN(new_n616_));
  AOI22_X1  g415(.A1(new_n548_), .A2(KEYINPUT72), .B1(new_n616_), .B2(new_n545_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n548_), .A2(KEYINPUT72), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n553_), .B1(new_n617_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n554_), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT73), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n550_), .A2(new_n551_), .A3(new_n554_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT104), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n615_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n470_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT43), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT43), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n557_), .A2(new_n470_), .A3(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT105), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n613_), .B1(new_n628_), .B2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n612_), .B1(new_n632_), .B2(KEYINPUT44), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n630_), .A2(KEYINPUT105), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n630_), .A2(KEYINPUT105), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n627_), .B1(new_n615_), .B2(new_n624_), .ZN(new_n636_));
  OAI22_X1  g435(.A1(new_n634_), .A2(new_n635_), .B1(new_n636_), .B2(new_n629_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n613_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT44), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n639_), .A2(KEYINPUT106), .A3(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n633_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n637_), .A2(KEYINPUT44), .A3(new_n638_), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n643_), .A2(G29gat), .A3(new_n573_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n611_), .B1(new_n642_), .B2(new_n644_), .ZN(G1328gat));
  INV_X1    g444(.A(G36gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n610_), .A2(new_n646_), .A3(new_n587_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT45), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n643_), .A2(new_n587_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n649_), .B1(new_n633_), .B2(new_n641_), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n648_), .B1(new_n650_), .B2(new_n646_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT46), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT46), .B(new_n648_), .C1(new_n650_), .C2(new_n646_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1329gat));
  NAND2_X1  g454(.A1(new_n610_), .A2(new_n326_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(KEYINPUT107), .B(G43gat), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n327_), .A2(new_n270_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n643_), .A2(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n659_), .B1(new_n642_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(G1330gat));
  AOI21_X1  g463(.A(G50gat), .B1(new_n610_), .B2(new_n453_), .ZN(new_n665_));
  AND3_X1   g464(.A1(new_n643_), .A2(G50gat), .A3(new_n453_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n665_), .B1(new_n642_), .B2(new_n666_), .ZN(G1331gat));
  INV_X1    g466(.A(new_n264_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n569_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n578_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G57gat), .B1(new_n670_), .B2(new_n466_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n264_), .A2(new_n581_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n627_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n570_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n573_), .A2(new_n356_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n671_), .B1(new_n675_), .B2(new_n676_), .ZN(G1332gat));
  OAI21_X1  g476(.A(G64gat), .B1(new_n670_), .B2(new_n465_), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n678_), .B(KEYINPUT48), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n465_), .A2(G64gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n675_), .B2(new_n680_), .ZN(G1333gat));
  OAI21_X1  g480(.A(G71gat), .B1(new_n670_), .B2(new_n327_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT49), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n327_), .A2(G71gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n675_), .B2(new_n684_), .ZN(G1334gat));
  OAI21_X1  g484(.A(G78gat), .B1(new_n670_), .B2(new_n454_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n686_), .B(KEYINPUT50), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n454_), .A2(G78gat), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT109), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n687_), .B1(new_n675_), .B2(new_n689_), .ZN(G1335gat));
  NOR2_X1   g489(.A1(new_n673_), .A2(new_n579_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n637_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(G85gat), .B1(new_n692_), .B2(new_n466_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n674_), .A2(new_n609_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n573_), .A2(new_n210_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n693_), .B1(new_n694_), .B2(new_n695_), .ZN(G1336gat));
  NOR3_X1   g495(.A1(new_n692_), .A2(new_n211_), .A3(new_n465_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n211_), .B1(new_n694_), .B2(new_n465_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n698_), .B(KEYINPUT110), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n697_), .A2(new_n699_), .ZN(G1337gat));
  NOR3_X1   g499(.A1(new_n694_), .A2(new_n215_), .A3(new_n327_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n637_), .A2(new_n326_), .A3(new_n691_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n701_), .B1(new_n702_), .B2(G99gat), .ZN(new_n703_));
  XOR2_X1   g502(.A(KEYINPUT111), .B(KEYINPUT51), .Z(new_n704_));
  XNOR2_X1  g503(.A(new_n703_), .B(new_n704_), .ZN(G1338gat));
  OR3_X1    g504(.A1(new_n694_), .A2(G106gat), .A3(new_n454_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n637_), .A2(new_n453_), .A3(new_n691_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(G106gat), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n708_), .A2(KEYINPUT52), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n708_), .A2(KEYINPUT52), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT112), .B(KEYINPUT53), .Z(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(G1339gat));
  NOR2_X1   g512(.A1(new_n587_), .A2(new_n466_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n467_), .ZN(new_n715_));
  INV_X1    g514(.A(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT58), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT114), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT55), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n248_), .A2(new_n718_), .A3(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n244_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(new_n250_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n719_), .B1(new_n248_), .B2(new_n718_), .ZN(new_n724_));
  OAI211_X1 g523(.A(KEYINPUT56), .B(new_n256_), .C1(new_n723_), .C2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT116), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n248_), .A2(new_n718_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT55), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(new_n720_), .A3(new_n722_), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n730_), .A2(KEYINPUT116), .A3(KEYINPUT56), .A4(new_n256_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n727_), .A2(new_n731_), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n256_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT117), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT56), .ZN(new_n735_));
  AND3_X1   g534(.A1(new_n733_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n733_), .B2(new_n735_), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n732_), .A2(new_n736_), .A3(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n503_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n489_), .A2(new_n491_), .A3(new_n497_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n497_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n502_), .B1(new_n495_), .B2(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n739_), .B1(new_n740_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n259_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n717_), .B1(new_n738_), .B2(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n733_), .A2(new_n735_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(KEYINPUT117), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n733_), .A2(new_n734_), .A3(new_n735_), .ZN(new_n748_));
  NAND4_X1  g547(.A1(new_n747_), .A2(new_n748_), .A3(new_n727_), .A4(new_n731_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n749_), .A2(KEYINPUT58), .A3(new_n259_), .A4(new_n743_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n745_), .A2(new_n557_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n260_), .A2(new_n743_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n581_), .A2(new_n259_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n746_), .B2(new_n725_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n752_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  AOI211_X1 g555(.A(KEYINPUT115), .B(new_n753_), .C1(new_n746_), .C2(new_n725_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n576_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT57), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  OAI211_X1 g559(.A(KEYINPUT57), .B(new_n576_), .C1(new_n756_), .C2(new_n757_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n751_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(new_n569_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n669_), .A2(new_n264_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n669_), .A2(new_n264_), .A3(KEYINPUT113), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n764_), .B1(new_n557_), .B2(new_n769_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n623_), .A2(KEYINPUT54), .A3(new_n767_), .A4(new_n768_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT118), .B1(new_n763_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n775_), .B(new_n772_), .C1(new_n762_), .C2(new_n569_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n716_), .B1(new_n774_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(G113gat), .B1(new_n778_), .B2(new_n581_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT120), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(KEYINPUT59), .ZN(new_n781_));
  XOR2_X1   g580(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n782_));
  NAND2_X1  g581(.A1(new_n716_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n783_), .B1(new_n763_), .B2(new_n773_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n780_), .B1(new_n781_), .B2(new_n785_), .ZN(new_n786_));
  AOI211_X1 g585(.A(KEYINPUT120), .B(new_n784_), .C1(new_n777_), .C2(KEYINPUT59), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n509_), .A2(G113gat), .A3(new_n513_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n779_), .B1(new_n788_), .B2(new_n789_), .ZN(G1340gat));
  NAND3_X1  g589(.A1(new_n781_), .A2(new_n668_), .A3(new_n785_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(G120gat), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n264_), .A2(KEYINPUT60), .A3(G120gat), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n793_), .B1(KEYINPUT60), .B2(G120gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n792_), .B1(new_n777_), .B2(new_n794_), .ZN(G1341gat));
  AOI21_X1  g594(.A(G127gat), .B1(new_n778_), .B2(new_n579_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n579_), .A2(KEYINPUT121), .A3(G127gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(KEYINPUT121), .B2(G127gat), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n796_), .B1(new_n788_), .B2(new_n798_), .ZN(G1342gat));
  AOI21_X1  g598(.A(G134gat), .B1(new_n778_), .B2(new_n577_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n557_), .A2(G134gat), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n788_), .B2(new_n801_), .ZN(G1343gat));
  OAI211_X1 g601(.A(new_n468_), .B(new_n714_), .C1(new_n774_), .C2(new_n776_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n581_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  XOR2_X1   g604(.A(KEYINPUT122), .B(G141gat), .Z(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(G1344gat));
  INV_X1    g606(.A(new_n803_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n668_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g609(.A(new_n468_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n762_), .A2(new_n569_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n775_), .B1(new_n812_), .B2(new_n772_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n763_), .A2(KEYINPUT118), .A3(new_n773_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n811_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT123), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n579_), .A4(new_n714_), .ZN(new_n817_));
  OAI21_X1  g616(.A(KEYINPUT123), .B1(new_n803_), .B2(new_n569_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(KEYINPUT61), .B(G155gat), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n820_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n817_), .A2(new_n818_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1346gat));
  NOR3_X1   g623(.A1(new_n803_), .A2(new_n337_), .A3(new_n626_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n808_), .A2(new_n577_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n826_), .B2(new_n337_), .ZN(G1347gat));
  NOR2_X1   g626(.A1(new_n812_), .A2(new_n772_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n465_), .A2(new_n573_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n326_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(new_n454_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n828_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  OAI21_X1  g633(.A(G169gat), .B1(new_n834_), .B2(new_n804_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT62), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n835_), .A2(new_n836_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n833_), .A2(new_n581_), .A3(new_n303_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(G1348gat));
  INV_X1    g639(.A(G176gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n841_), .B1(new_n834_), .B2(new_n264_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n453_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n843_), .A2(G176gat), .A3(new_n668_), .A4(new_n831_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT124), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n842_), .A2(new_n844_), .A3(KEYINPUT124), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(G1349gat));
  NOR3_X1   g648(.A1(new_n834_), .A2(new_n569_), .A3(new_n289_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n843_), .A2(new_n579_), .A3(new_n831_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n280_), .ZN(G1350gat));
  OAI21_X1  g651(.A(G190gat), .B1(new_n834_), .B2(new_n623_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n833_), .A2(new_n577_), .A3(new_n390_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(G1351gat));
  NAND2_X1  g654(.A1(new_n815_), .A2(new_n829_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(G197gat), .B1(new_n857_), .B2(new_n581_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n856_), .A2(new_n369_), .A3(new_n804_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(G1352gat));
  NAND3_X1  g659(.A1(new_n857_), .A2(new_n375_), .A3(new_n668_), .ZN(new_n861_));
  OAI21_X1  g660(.A(G204gat), .B1(new_n856_), .B2(new_n264_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1353gat));
  AOI21_X1  g662(.A(new_n569_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n815_), .A2(new_n829_), .A3(new_n864_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(KEYINPUT125), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n866_));
  XOR2_X1   g665(.A(new_n866_), .B(KEYINPUT126), .Z(new_n867_));
  OAI21_X1  g666(.A(KEYINPUT125), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n865_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n867_), .B1(new_n865_), .B2(new_n868_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1354gat));
  NAND2_X1  g671(.A1(new_n857_), .A2(new_n577_), .ZN(new_n873_));
  INV_X1    g672(.A(G218gat), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n623_), .A2(new_n874_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT127), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n873_), .A2(new_n874_), .B1(new_n857_), .B2(new_n876_), .ZN(G1355gat));
endmodule


