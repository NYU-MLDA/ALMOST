//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n765_, new_n766_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n914_, new_n915_, new_n917_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n924_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n202_));
  XOR2_X1   g001(.A(G8gat), .B(G36gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT23), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT72), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT72), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n208_), .A2(new_n211_), .A3(KEYINPUT23), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT73), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n208_), .A2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(KEYINPUT73), .A2(G183gat), .A3(G190gat), .ZN(new_n216_));
  AOI21_X1  g015(.A(KEYINPUT23), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G169gat), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  OAI22_X1  g019(.A1(new_n213_), .A2(new_n217_), .B1(KEYINPUT24), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT74), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OAI221_X1 g022(.A(KEYINPUT74), .B1(KEYINPUT24), .B2(new_n220_), .C1(new_n213_), .C2(new_n217_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(G190gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT26), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT26), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G190gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(G183gat), .ZN(new_n232_));
  OR2_X1    g031(.A1(new_n232_), .A2(KEYINPUT25), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n231_), .B1(KEYINPUT71), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT25), .B(G183gat), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n235_), .A2(KEYINPUT71), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n226_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n223_), .A2(new_n224_), .A3(new_n237_), .ZN(new_n238_));
  XNOR2_X1  g037(.A(KEYINPUT77), .B(G176gat), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT75), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(new_n218_), .A3(KEYINPUT22), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT22), .ZN(new_n242_));
  OAI21_X1  g041(.A(KEYINPUT75), .B1(new_n242_), .B2(G169gat), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n241_), .A3(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT76), .B1(new_n218_), .B2(KEYINPUT22), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT76), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(new_n242_), .A3(G169gat), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n245_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n225_), .B1(new_n244_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT78), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n232_), .A2(new_n227_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT23), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n208_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n216_), .ZN(new_n255_));
  AOI21_X1  g054(.A(KEYINPUT73), .B1(G183gat), .B2(G190gat), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n252_), .B(new_n254_), .C1(new_n257_), .C2(new_n253_), .ZN(new_n258_));
  OAI211_X1 g057(.A(KEYINPUT78), .B(new_n225_), .C1(new_n244_), .C2(new_n248_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n251_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n238_), .A2(new_n260_), .ZN(new_n261_));
  XOR2_X1   g060(.A(G211gat), .B(G218gat), .Z(new_n262_));
  INV_X1    g061(.A(G197gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT83), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT83), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(G197gat), .ZN(new_n266_));
  INV_X1    g065(.A(G204gat), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n264_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT21), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n269_), .B1(G197gat), .B2(G204gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n262_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(KEYINPUT84), .B(KEYINPUT21), .Z(new_n272_));
  AOI21_X1  g071(.A(new_n267_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(G197gat), .A2(G204gat), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n272_), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n273_), .A2(new_n274_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G211gat), .B(G218gat), .ZN(new_n278_));
  NOR2_X1   g077(.A1(new_n278_), .A2(new_n269_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n276_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n261_), .A2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G226gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT19), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT20), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n208_), .A2(new_n211_), .A3(KEYINPUT23), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n211_), .B1(new_n208_), .B2(KEYINPUT23), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n253_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n289_), .A2(new_n290_), .B1(new_n232_), .B2(new_n227_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT22), .B(G169gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n239_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(new_n225_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT24), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n295_), .A2(KEYINPUT88), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(KEYINPUT88), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n225_), .B(new_n220_), .C1(new_n296_), .C2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n235_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n300_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n298_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n302_));
  OAI21_X1  g101(.A(new_n254_), .B1(new_n257_), .B2(new_n253_), .ZN(new_n303_));
  OAI22_X1  g102(.A1(new_n291_), .A2(new_n294_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n282_), .B(new_n286_), .C1(new_n281_), .C2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT89), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n271_), .A2(new_n275_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n238_), .A2(new_n260_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n285_), .B1(new_n304_), .B2(new_n281_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n306_), .B1(new_n310_), .B2(new_n284_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n284_), .ZN(new_n312_));
  AOI211_X1 g111(.A(KEYINPUT89), .B(new_n312_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n313_));
  OAI211_X1 g112(.A(new_n207_), .B(new_n305_), .C1(new_n311_), .C2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  AND3_X1   g114(.A1(new_n308_), .A2(new_n312_), .A3(new_n309_), .ZN(new_n316_));
  XOR2_X1   g115(.A(KEYINPUT96), .B(KEYINPUT20), .Z(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n318_), .B1(new_n304_), .B2(new_n281_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT97), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT97), .ZN(new_n321_));
  OAI211_X1 g120(.A(new_n321_), .B(new_n318_), .C1(new_n304_), .C2(new_n281_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n282_), .A2(new_n320_), .A3(new_n322_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n316_), .B1(new_n323_), .B2(new_n284_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT27), .B1(new_n324_), .B2(new_n207_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n202_), .B1(new_n315_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n207_), .ZN(new_n327_));
  AND2_X1   g126(.A1(new_n323_), .A2(new_n284_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n327_), .B1(new_n328_), .B2(new_n316_), .ZN(new_n329_));
  NAND4_X1  g128(.A1(new_n329_), .A2(KEYINPUT99), .A3(KEYINPUT27), .A4(new_n314_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n305_), .B1(new_n311_), .B2(new_n313_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n327_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT91), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(new_n314_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT27), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n332_), .A2(KEYINPUT91), .A3(new_n327_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n335_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n331_), .A2(new_n338_), .ZN(new_n339_));
  AND3_X1   g138(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  OAI22_X1  g141(.A1(KEYINPUT80), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI211_X1 g144(.A(KEYINPUT80), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n342_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348_));
  NOR2_X1   g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n347_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT1), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n349_), .A2(KEYINPUT1), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n353_), .B1(new_n354_), .B2(new_n348_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(G141gat), .A2(G148gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(KEYINPUT79), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT79), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(G141gat), .B2(G148gat), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n357_), .A2(new_n359_), .B1(G141gat), .B2(G148gat), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n351_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n363_), .A3(KEYINPUT29), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n347_), .A2(new_n350_), .B1(new_n355_), .B2(new_n360_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT81), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G228gat), .ZN(new_n369_));
  INV_X1    g168(.A(G233gat), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n370_), .A2(KEYINPUT82), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(KEYINPUT82), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n369_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(new_n307_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT86), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT85), .B(KEYINPUT29), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n281_), .B1(new_n365_), .B2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n376_), .B1(new_n378_), .B2(new_n373_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n377_), .B1(new_n351_), .B2(new_n361_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n376_), .B(new_n373_), .C1(new_n380_), .C2(new_n307_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n375_), .B1(new_n379_), .B2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G22gat), .B(G50gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT28), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n365_), .A2(new_n386_), .A3(new_n366_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n386_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n385_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n351_), .A2(new_n366_), .A3(new_n361_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT28), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n392_), .A2(new_n387_), .A3(new_n384_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n390_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n383_), .A2(KEYINPUT87), .A3(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n373_), .B1(new_n380_), .B2(new_n307_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT86), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n397_), .A2(new_n381_), .B1(new_n368_), .B2(new_n374_), .ZN(new_n398_));
  AND3_X1   g197(.A1(new_n392_), .A2(new_n387_), .A3(new_n384_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n384_), .B1(new_n392_), .B2(new_n387_), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT87), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT87), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n390_), .A2(new_n402_), .A3(new_n393_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n398_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  XOR2_X1   g203(.A(G78gat), .B(G106gat), .Z(new_n405_));
  AND3_X1   g204(.A1(new_n395_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(new_n395_), .B2(new_n404_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n339_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G71gat), .B(G99gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n411_), .B(G43gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n261_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(G127gat), .B(G134gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G113gat), .B(G120gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n414_), .B(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n413_), .B(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G227gat), .A2(G233gat), .ZN(new_n419_));
  INV_X1    g218(.A(G15gat), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n419_), .B(new_n420_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n421_), .B(KEYINPUT30), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT31), .ZN(new_n423_));
  XOR2_X1   g222(.A(new_n418_), .B(new_n423_), .Z(new_n424_));
  NAND2_X1  g223(.A1(new_n362_), .A2(new_n417_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n365_), .A2(new_n416_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(KEYINPUT4), .A3(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT4), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n362_), .A2(new_n417_), .A3(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT92), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n362_), .A2(new_n417_), .A3(KEYINPUT92), .A4(new_n428_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n427_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G225gat), .A2(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n433_), .A2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G1gat), .B(G29gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G57gat), .B(G85gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n444_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n436_), .A2(new_n446_), .A3(new_n438_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n445_), .A2(KEYINPUT98), .A3(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT98), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n446_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n450_));
  AOI211_X1 g249(.A(new_n444_), .B(new_n437_), .C1(new_n433_), .C2(new_n435_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n449_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n448_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n410_), .A2(new_n424_), .A3(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n408_), .A2(new_n453_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n331_), .A2(new_n457_), .A3(new_n338_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT100), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n331_), .A2(new_n457_), .A3(new_n338_), .A4(KEYINPUT100), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n433_), .A2(new_n435_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n425_), .A2(new_n426_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n465_), .A2(new_n435_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n446_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n464_), .A2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n445_), .B1(new_n463_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n450_), .A2(KEYINPUT33), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n471_), .B1(new_n335_), .B2(new_n337_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT94), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n207_), .A2(KEYINPUT32), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n324_), .A2(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n305_), .B(new_n475_), .C1(new_n311_), .C2(new_n313_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT95), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n478_), .A2(new_n479_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n477_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n482_), .B1(new_n472_), .B2(KEYINPUT94), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n408_), .B1(new_n474_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n462_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n424_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n456_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT70), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT68), .B(G15gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(G22gat), .ZN(new_n490_));
  INV_X1    g289(.A(G1gat), .ZN(new_n491_));
  INV_X1    g290(.A(G8gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(KEYINPUT14), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n490_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT69), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(G1gat), .B(G8gat), .Z(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n494_), .B(KEYINPUT69), .ZN(new_n499_));
  INV_X1    g298(.A(new_n497_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n498_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(G29gat), .B(G36gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT65), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G43gat), .B(G50gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n502_), .A2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(KEYINPUT15), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n512_), .A2(new_n498_), .A3(new_n501_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G229gat), .A2(G233gat), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n508_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n498_), .A2(new_n501_), .A3(new_n506_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n514_), .B1(new_n508_), .B2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n488_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(G113gat), .B(G141gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G169gat), .B(G197gat), .ZN(new_n520_));
  XOR2_X1   g319(.A(new_n519_), .B(new_n520_), .Z(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n518_), .A2(new_n522_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n488_), .B(new_n521_), .C1(new_n515_), .C2(new_n517_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(G230gat), .A2(G233gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G99gat), .A2(G106gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT6), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(G106gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT10), .B(G99gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n530_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(G85gat), .ZN(new_n535_));
  INV_X1    g334(.A(G92gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT9), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G85gat), .A2(G92gat), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT64), .ZN(new_n540_));
  AND3_X1   g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n538_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n540_), .B1(new_n539_), .B2(new_n538_), .ZN(new_n542_));
  OAI221_X1 g341(.A(new_n537_), .B1(new_n538_), .B2(new_n539_), .C1(new_n541_), .C2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n534_), .A2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n537_), .A2(new_n539_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT7), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n545_), .B1(new_n530_), .B2(new_n550_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n551_), .A2(KEYINPUT8), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n551_), .A2(KEYINPUT8), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n544_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n557_));
  XOR2_X1   g356(.A(G71gat), .B(G78gat), .Z(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n557_), .A2(new_n558_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n554_), .A2(new_n562_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n561_), .B(new_n544_), .C1(new_n552_), .C2(new_n553_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n563_), .A2(new_n564_), .A3(KEYINPUT12), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n554_), .A2(new_n562_), .A3(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n527_), .B1(new_n565_), .B2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n526_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G120gat), .B(G148gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT5), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G176gat), .B(G204gat), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n572_), .B(new_n573_), .Z(new_n574_));
  NOR2_X1   g373(.A1(new_n570_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n570_), .A2(new_n574_), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n576_), .A2(KEYINPUT13), .A3(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT13), .B1(new_n576_), .B2(new_n577_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(G231gat), .A2(G233gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n561_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n502_), .B(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(G127gat), .B(G155gat), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT16), .ZN(new_n585_));
  XOR2_X1   g384(.A(G183gat), .B(G211gat), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT17), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n583_), .A2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT17), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n587_), .A2(new_n591_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n590_), .B1(new_n592_), .B2(new_n583_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G134gat), .B(G162gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT36), .Z(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n554_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n600_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G232gat), .A2(G233gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT34), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n603_), .A2(KEYINPUT35), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n554_), .A2(new_n506_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n601_), .A2(new_n604_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(KEYINPUT35), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  OAI211_X1 g407(.A(KEYINPUT35), .B(new_n603_), .C1(new_n601_), .C2(new_n605_), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n599_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(KEYINPUT67), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT67), .ZN(new_n612_));
  AOI211_X1 g411(.A(new_n612_), .B(new_n599_), .C1(new_n608_), .C2(new_n609_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n597_), .A2(KEYINPUT36), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n608_), .A2(new_n615_), .A3(new_n609_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT66), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n594_), .B1(new_n614_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n616_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(new_n610_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n621_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(KEYINPUT37), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n580_), .B(new_n593_), .C1(new_n619_), .C2(new_n623_), .ZN(new_n624_));
  NOR3_X1   g423(.A1(new_n487_), .A2(new_n525_), .A3(new_n624_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n625_), .A2(new_n491_), .A3(new_n453_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  XOR2_X1   g426(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n628_));
  OR2_X1    g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n487_), .A2(new_n621_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n580_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n593_), .ZN(new_n632_));
  NOR3_X1   g431(.A1(new_n631_), .A2(new_n525_), .A3(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n630_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(G1gat), .B1(new_n635_), .B2(new_n454_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n627_), .A2(new_n628_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n629_), .A2(new_n636_), .A3(new_n637_), .ZN(G1324gat));
  INV_X1    g437(.A(new_n339_), .ZN(new_n639_));
  OR3_X1    g438(.A1(new_n635_), .A2(KEYINPUT103), .A3(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(KEYINPUT103), .B1(new_n635_), .B2(new_n639_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(G8gat), .A3(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(KEYINPUT104), .B(KEYINPUT39), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n643_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n640_), .A2(G8gat), .A3(new_n645_), .A4(new_n641_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n625_), .A2(new_n492_), .A3(new_n339_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(KEYINPUT102), .Z(new_n648_));
  NAND3_X1  g447(.A1(new_n644_), .A2(new_n646_), .A3(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND4_X1  g450(.A1(new_n644_), .A2(KEYINPUT40), .A3(new_n646_), .A4(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1325gat));
  AOI21_X1  g452(.A(new_n420_), .B1(new_n634_), .B2(new_n424_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT41), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n625_), .A2(new_n420_), .A3(new_n424_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1326gat));
  INV_X1    g456(.A(G22gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n658_), .B1(new_n634_), .B2(new_n409_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n625_), .A2(new_n658_), .A3(new_n409_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT106), .ZN(G1327gat));
  NAND2_X1  g463(.A1(new_n335_), .A2(new_n337_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n665_), .A2(new_n470_), .A3(new_n469_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT94), .ZN(new_n667_));
  OR2_X1    g466(.A1(new_n480_), .A2(new_n481_), .ZN(new_n668_));
  AOI22_X1  g467(.A1(new_n666_), .A2(new_n667_), .B1(new_n668_), .B2(new_n477_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n409_), .B1(new_n669_), .B2(new_n473_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n460_), .A2(new_n461_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n486_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n672_), .A2(new_n455_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n525_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n622_), .A2(new_n593_), .ZN(new_n675_));
  AND4_X1   g474(.A1(new_n673_), .A2(new_n674_), .A3(new_n580_), .A4(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(G29gat), .B1(new_n676_), .B2(new_n453_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT43), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n619_), .A2(new_n623_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n424_), .B1(new_n462_), .B2(new_n484_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n678_), .B(new_n679_), .C1(new_n680_), .C2(new_n456_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n673_), .A2(KEYINPUT107), .A3(new_n678_), .A4(new_n679_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n679_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT43), .B1(new_n487_), .B2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n683_), .A2(new_n684_), .A3(new_n686_), .ZN(new_n687_));
  NOR3_X1   g486(.A1(new_n631_), .A2(new_n525_), .A3(new_n593_), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT44), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n687_), .A2(KEYINPUT44), .A3(new_n688_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT108), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT108), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n687_), .A2(new_n692_), .A3(KEYINPUT44), .A4(new_n688_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n689_), .B1(new_n691_), .B2(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n453_), .A2(G29gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n677_), .B1(new_n694_), .B2(new_n695_), .ZN(G1328gat));
  XNOR2_X1  g495(.A(KEYINPUT109), .B(KEYINPUT46), .ZN(new_n697_));
  INV_X1    g496(.A(G36gat), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n691_), .A2(new_n693_), .ZN(new_n699_));
  NOR2_X1   g498(.A1(new_n689_), .A2(new_n639_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n698_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n676_), .A2(new_n698_), .A3(new_n339_), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT45), .Z(new_n703_));
  OAI21_X1  g502(.A(new_n697_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT110), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n701_), .A2(new_n703_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(KEYINPUT46), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n708_), .B(new_n697_), .C1(new_n701_), .C2(new_n703_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n705_), .A2(new_n707_), .A3(new_n709_), .ZN(G1329gat));
  NAND3_X1  g509(.A1(new_n694_), .A2(G43gat), .A3(new_n424_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n676_), .A2(new_n424_), .ZN(new_n713_));
  OR2_X1    g512(.A1(new_n713_), .A2(G43gat), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT111), .ZN(new_n715_));
  OAI21_X1  g514(.A(KEYINPUT47), .B1(new_n712_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n715_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT47), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n718_), .A3(new_n711_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n719_), .ZN(G1330gat));
  AOI21_X1  g519(.A(G50gat), .B1(new_n676_), .B2(new_n409_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n409_), .A2(G50gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n694_), .B2(new_n722_), .ZN(G1331gat));
  NOR2_X1   g522(.A1(new_n487_), .A2(new_n674_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(new_n724_), .B(KEYINPUT112), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n618_), .A2(new_n614_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT37), .ZN(new_n727_));
  INV_X1    g526(.A(new_n623_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n632_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  AND3_X1   g528(.A1(new_n725_), .A2(new_n631_), .A3(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(G57gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n731_), .A3(new_n453_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n580_), .A2(new_n674_), .A3(new_n632_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n630_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(G57gat), .B1(new_n735_), .B2(new_n454_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n732_), .A2(new_n736_), .ZN(G1332gat));
  INV_X1    g536(.A(G64gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n734_), .B2(new_n339_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT48), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n730_), .A2(new_n738_), .A3(new_n339_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT113), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n742_), .B(new_n743_), .ZN(G1333gat));
  NOR2_X1   g543(.A1(new_n486_), .A2(G71gat), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT114), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n730_), .A2(new_n746_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G71gat), .B1(new_n735_), .B2(new_n486_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(KEYINPUT49), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(KEYINPUT49), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n747_), .B1(new_n749_), .B2(new_n750_), .ZN(G1334gat));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n734_), .B2(new_n409_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT50), .Z(new_n754_));
  NAND3_X1  g553(.A1(new_n730_), .A2(new_n752_), .A3(new_n409_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1335gat));
  AND3_X1   g555(.A1(new_n725_), .A2(new_n631_), .A3(new_n675_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G85gat), .B1(new_n757_), .B2(new_n453_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT115), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n580_), .A2(new_n674_), .A3(new_n593_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n687_), .A2(new_n760_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT116), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n454_), .A2(new_n535_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n759_), .B1(new_n762_), .B2(new_n763_), .ZN(G1336gat));
  NAND3_X1  g563(.A1(new_n757_), .A2(new_n536_), .A3(new_n339_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n762_), .A2(new_n339_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(new_n536_), .ZN(G1337gat));
  NAND3_X1  g566(.A1(new_n757_), .A2(new_n424_), .A3(new_n533_), .ZN(new_n768_));
  OAI21_X1  g567(.A(G99gat), .B1(new_n761_), .B2(new_n486_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g570(.A1(new_n757_), .A2(new_n531_), .A3(new_n409_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n687_), .A2(new_n409_), .A3(new_n760_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT117), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(G106gat), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n774_), .B1(new_n773_), .B2(G106gat), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n776_), .A2(new_n777_), .A3(KEYINPUT52), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n773_), .A2(G106gat), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(KEYINPUT117), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n779_), .B1(new_n781_), .B2(new_n775_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n772_), .B1(new_n778_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n772_), .C1(new_n778_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  INV_X1    g586(.A(KEYINPUT120), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n523_), .A2(new_n524_), .A3(new_n576_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n565_), .A2(new_n527_), .A3(new_n567_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(KEYINPUT55), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n791_), .A2(new_n568_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT118), .ZN(new_n793_));
  AOI211_X1 g592(.A(KEYINPUT55), .B(new_n527_), .C1(new_n565_), .C2(new_n567_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n568_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(KEYINPUT55), .A3(new_n790_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n794_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT118), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n574_), .B1(new_n795_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT56), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n793_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n797_), .A2(KEYINPUT118), .A3(new_n798_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n803_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(KEYINPUT56), .A3(new_n574_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n789_), .B1(new_n802_), .B2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n516_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n506_), .B1(new_n498_), .B2(new_n501_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n514_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n514_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n508_), .A2(new_n513_), .A3(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n522_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n521_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT119), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n814_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n521_), .B1(new_n810_), .B2(new_n812_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n811_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n508_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n522_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT119), .B1(new_n818_), .B2(new_n821_), .ZN(new_n822_));
  AOI22_X1  g621(.A1(new_n817_), .A2(new_n822_), .B1(new_n577_), .B2(new_n576_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n622_), .B1(new_n807_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT57), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n575_), .B1(new_n817_), .B2(new_n822_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT56), .B1(new_n805_), .B2(new_n574_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n574_), .ZN(new_n829_));
  AOI211_X1 g628(.A(new_n801_), .B(new_n829_), .C1(new_n803_), .C2(new_n804_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n827_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT58), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n827_), .B(KEYINPUT58), .C1(new_n828_), .C2(new_n830_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n679_), .A3(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(KEYINPUT57), .B(new_n622_), .C1(new_n807_), .C2(new_n823_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n826_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n729_), .A2(new_n838_), .A3(new_n525_), .A4(new_n580_), .ZN(new_n839_));
  OAI21_X1  g638(.A(KEYINPUT54), .B1(new_n624_), .B2(new_n674_), .ZN(new_n840_));
  AOI22_X1  g639(.A1(new_n837_), .A2(new_n632_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n410_), .A2(new_n424_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n841_), .A2(new_n454_), .A3(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n788_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n837_), .A2(new_n632_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n839_), .A2(new_n840_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n842_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n453_), .A3(new_n849_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n850_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n848_), .A2(new_n844_), .A3(new_n453_), .A4(new_n849_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT121), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n841_), .A2(new_n454_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n844_), .A4(new_n849_), .ZN(new_n856_));
  AOI22_X1  g655(.A1(new_n845_), .A2(new_n851_), .B1(new_n853_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  OAI21_X1  g657(.A(G113gat), .B1(new_n858_), .B2(new_n525_), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n525_), .A2(G113gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n850_), .B2(new_n860_), .ZN(G1340gat));
  NAND2_X1  g660(.A1(new_n845_), .A2(new_n851_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n853_), .A2(new_n856_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n862_), .A2(new_n631_), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT122), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n580_), .A2(G120gat), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n843_), .B1(KEYINPUT60), .B2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n857_), .A2(KEYINPUT122), .A3(new_n631_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n866_), .A2(new_n868_), .A3(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G120gat), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n868_), .A2(KEYINPUT60), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1341gat));
  OAI21_X1  g672(.A(G127gat), .B1(new_n858_), .B2(new_n632_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n632_), .A2(G127gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n850_), .B2(new_n875_), .ZN(G1342gat));
  INV_X1    g675(.A(G134gat), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n857_), .B2(new_n679_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n850_), .A2(G134gat), .A3(new_n622_), .ZN(new_n879_));
  OR3_X1    g678(.A1(new_n878_), .A2(KEYINPUT123), .A3(new_n879_), .ZN(new_n880_));
  OAI21_X1  g679(.A(KEYINPUT123), .B1(new_n878_), .B2(new_n879_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1343gat));
  NOR3_X1   g681(.A1(new_n339_), .A2(new_n424_), .A3(new_n408_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n854_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n674_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n631_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g688(.A1(new_n884_), .A2(new_n632_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT61), .B(G155gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  OAI21_X1  g691(.A(G162gat), .B1(new_n884_), .B2(new_n685_), .ZN(new_n893_));
  OR2_X1    g692(.A1(new_n622_), .A2(G162gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n884_), .B2(new_n894_), .ZN(G1347gat));
  NAND3_X1  g694(.A1(new_n424_), .A2(new_n408_), .A3(new_n454_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n841_), .A2(new_n639_), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n674_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n898_), .A2(KEYINPUT124), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n218_), .B1(new_n898_), .B2(KEYINPUT124), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT62), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n897_), .A2(new_n292_), .A3(new_n674_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n899_), .A2(KEYINPUT62), .A3(new_n900_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n903_), .A2(new_n904_), .A3(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(KEYINPUT125), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n903_), .A2(new_n908_), .A3(new_n904_), .A4(new_n905_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1348gat));
  NAND2_X1  g709(.A1(new_n897_), .A2(new_n631_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n219_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n912_), .B1(new_n239_), .B2(new_n911_), .ZN(G1349gat));
  NAND2_X1  g712(.A1(new_n897_), .A2(new_n593_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n914_), .A2(new_n235_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n915_), .B1(new_n232_), .B2(new_n914_), .ZN(G1350gat));
  AOI21_X1  g715(.A(new_n227_), .B1(new_n897_), .B2(new_n679_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n622_), .A2(new_n231_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n897_), .B2(new_n918_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(KEYINPUT126), .ZN(G1351gat));
  AND4_X1   g719(.A1(new_n486_), .A2(new_n848_), .A3(new_n457_), .A4(new_n339_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n674_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n631_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G204gat), .ZN(G1353gat));
  AND2_X1   g724(.A1(new_n921_), .A2(new_n593_), .ZN(new_n926_));
  XOR2_X1   g725(.A(KEYINPUT63), .B(G211gat), .Z(new_n927_));
  AOI21_X1  g726(.A(KEYINPUT127), .B1(new_n926_), .B2(new_n927_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n929_));
  MUX2_X1   g728(.A(new_n929_), .B(new_n927_), .S(new_n926_), .Z(new_n930_));
  AOI21_X1  g729(.A(new_n928_), .B1(new_n930_), .B2(KEYINPUT127), .ZN(G1354gat));
  INV_X1    g730(.A(G218gat), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n921_), .A2(new_n932_), .A3(new_n621_), .ZN(new_n933_));
  AND2_X1   g732(.A1(new_n921_), .A2(new_n679_), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n934_), .B2(new_n932_), .ZN(G1355gat));
endmodule


