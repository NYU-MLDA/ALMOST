//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n804_, new_n805_, new_n806_, new_n807_, new_n809_,
    new_n810_, new_n811_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n834_,
    new_n835_, new_n836_, new_n837_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n910_, new_n911_,
    new_n913_, new_n915_, new_n916_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n937_, new_n939_, new_n940_, new_n942_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n963_, new_n964_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G197gat), .B(G204gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT21), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT91), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT91), .ZN(new_n208_));
  INV_X1    g007(.A(G204gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(new_n209_), .A2(G197gat), .ZN(new_n210_));
  INV_X1    g009(.A(G197gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(G204gat), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n208_), .B(KEYINPUT21), .C1(new_n210_), .C2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(KEYINPUT92), .B1(new_n209_), .B2(G197gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT92), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(new_n211_), .A3(G204gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n209_), .A2(G197gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n214_), .A2(new_n216_), .A3(new_n205_), .A4(new_n217_), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n206_), .A2(new_n207_), .A3(new_n213_), .A4(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT93), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n207_), .A2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G211gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n222_), .A2(G218gat), .ZN(new_n223_));
  INV_X1    g022(.A(G218gat), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n224_), .A2(G211gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT93), .B1(new_n223_), .B2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n214_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n227_));
  NAND4_X1  g026(.A1(new_n221_), .A2(new_n226_), .A3(new_n227_), .A4(KEYINPUT21), .ZN(new_n228_));
  AND2_X1   g027(.A1(new_n219_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT97), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT96), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT22), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(G169gat), .ZN(new_n233_));
  INV_X1    g032(.A(G169gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(KEYINPUT22), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n231_), .B1(new_n233_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n234_), .A2(KEYINPUT22), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n232_), .A2(G169gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(new_n238_), .A3(KEYINPUT96), .ZN(new_n239_));
  AOI21_X1  g038(.A(G176gat), .B1(new_n236_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G183gat), .A2(G190gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT23), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(G183gat), .A2(G190gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n243_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(G169gat), .A2(G176gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n230_), .B1(new_n240_), .B2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G176gat), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n237_), .A2(new_n238_), .A3(KEYINPUT96), .ZN(new_n251_));
  AOI21_X1  g050(.A(KEYINPUT96), .B1(new_n237_), .B2(new_n238_), .ZN(new_n252_));
  OAI21_X1  g051(.A(new_n250_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n248_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(new_n254_), .A3(KEYINPUT97), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n249_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT81), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n257_), .A2(new_n234_), .A3(new_n250_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT81), .B1(G169gat), .B2(G176gat), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT95), .B(KEYINPUT24), .ZN(new_n261_));
  INV_X1    g060(.A(new_n247_), .ZN(new_n262_));
  OR3_X1    g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n261_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n243_), .A2(new_n245_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT25), .B(G183gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(G190gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .A4(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n229_), .B1(new_n256_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(G183gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT25), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT80), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(new_n271_), .B2(KEYINPUT25), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT25), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(KEYINPUT80), .A3(G183gat), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n267_), .A2(new_n272_), .A3(new_n274_), .A4(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT24), .ZN(new_n278_));
  INV_X1    g077(.A(new_n259_), .ZN(new_n279_));
  NOR3_X1   g078(.A1(KEYINPUT81), .A2(G169gat), .A3(G176gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n258_), .A2(KEYINPUT24), .A3(new_n247_), .A4(new_n259_), .ZN(new_n282_));
  NAND4_X1  g081(.A1(new_n277_), .A2(new_n281_), .A3(new_n265_), .A4(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n232_), .A2(new_n234_), .A3(new_n250_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n246_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n219_), .A2(new_n283_), .A3(new_n228_), .A4(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT20), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n203_), .B1(new_n270_), .B2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n256_), .A2(new_n229_), .A3(new_n269_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n203_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT20), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n219_), .A2(new_n228_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n283_), .A2(new_n286_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n292_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n290_), .A2(new_n291_), .A3(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  XNOR2_X1  g098(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(KEYINPUT32), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n289_), .A2(new_n296_), .A3(new_n303_), .ZN(new_n304_));
  NOR3_X1   g103(.A1(new_n270_), .A2(new_n203_), .A3(new_n288_), .ZN(new_n305_));
  OAI211_X1 g104(.A(new_n229_), .B(new_n269_), .C1(new_n240_), .C2(new_n248_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n291_), .B1(new_n306_), .B2(new_n295_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n305_), .A2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n304_), .B1(new_n308_), .B2(new_n303_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n310_), .B1(KEYINPUT1), .B2(new_n311_), .ZN(new_n312_));
  OR2_X1    g111(.A1(new_n311_), .A2(KEYINPUT1), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(G141gat), .A2(G148gat), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n314_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(G127gat), .B(G134gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(G113gat), .B(G120gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT3), .ZN(new_n323_));
  INV_X1    g122(.A(G141gat), .ZN(new_n324_));
  INV_X1    g123(.A(G148gat), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n323_), .A2(new_n324_), .A3(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT2), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n315_), .A2(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n326_), .A2(new_n328_), .A3(new_n329_), .A4(new_n330_), .ZN(new_n331_));
  XOR2_X1   g130(.A(G155gat), .B(G162gat), .Z(new_n332_));
  AND3_X1   g131(.A1(new_n331_), .A2(KEYINPUT86), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT86), .B1(new_n331_), .B2(new_n332_), .ZN(new_n334_));
  OAI211_X1 g133(.A(new_n319_), .B(new_n322_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n335_));
  AOI211_X1 g134(.A(new_n316_), .B(new_n317_), .C1(new_n312_), .C2(new_n313_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n331_), .A2(new_n332_), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT86), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n331_), .A2(KEYINPUT86), .A3(new_n332_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n336_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n320_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n321_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(new_n343_), .A3(KEYINPUT84), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT84), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n320_), .A2(new_n321_), .A3(KEYINPUT83), .ZN(new_n347_));
  AOI21_X1  g146(.A(KEYINPUT83), .B1(new_n320_), .B2(new_n321_), .ZN(new_n348_));
  OAI211_X1 g147(.A(new_n344_), .B(new_n346_), .C1(new_n347_), .C2(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n335_), .B(KEYINPUT4), .C1(new_n341_), .C2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT100), .ZN(new_n351_));
  INV_X1    g150(.A(new_n349_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n319_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT100), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n354_), .A2(new_n355_), .A3(KEYINPUT4), .A4(new_n335_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n351_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G225gat), .A2(G233gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n359_), .B1(new_n354_), .B2(KEYINPUT4), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n357_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n354_), .A2(new_n335_), .A3(new_n358_), .ZN(new_n363_));
  XOR2_X1   g162(.A(G1gat), .B(G29gat), .Z(new_n364_));
  XNOR2_X1  g163(.A(G57gat), .B(G85gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT101), .B(KEYINPUT0), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n362_), .A2(new_n363_), .A3(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n360_), .B1(new_n351_), .B2(new_n356_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n363_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n368_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n309_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT99), .ZN(new_n375_));
  AND3_X1   g174(.A1(new_n289_), .A2(new_n302_), .A3(new_n296_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n302_), .B1(new_n289_), .B2(new_n296_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n375_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n240_), .A2(new_n248_), .A3(new_n230_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT97), .B1(new_n253_), .B2(new_n254_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n269_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n293_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n288_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n291_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n290_), .A2(new_n291_), .A3(new_n295_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n301_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n288_), .B1(new_n293_), .B2(new_n381_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n302_), .B(new_n296_), .C1(new_n387_), .C2(new_n291_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(KEYINPUT99), .A3(new_n388_), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n371_), .A2(new_n372_), .A3(new_n368_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n378_), .A2(new_n389_), .B1(KEYINPUT33), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n354_), .A2(new_n335_), .A3(new_n359_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n368_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n354_), .A2(KEYINPUT4), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n394_), .A2(new_n359_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n393_), .B1(new_n357_), .B2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT33), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n396_), .B1(new_n370_), .B2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n374_), .B1(new_n391_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400_));
  OAI211_X1 g199(.A(new_n400_), .B(new_n319_), .C1(new_n333_), .C2(new_n334_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT28), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n339_), .A2(new_n340_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT28), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n403_), .A2(new_n404_), .A3(new_n400_), .A4(new_n319_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT87), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n402_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n406_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT89), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n411_), .A2(G228gat), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(G228gat), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n410_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT90), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n353_), .A2(KEYINPUT29), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT88), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n229_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n353_), .A2(KEYINPUT88), .A3(KEYINPUT29), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n415_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n416_), .A2(KEYINPUT94), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT94), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n353_), .A2(new_n422_), .A3(KEYINPUT29), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n293_), .A2(new_n415_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AND3_X1   g224(.A1(new_n421_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n409_), .B1(new_n420_), .B2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n404_), .B1(new_n341_), .B2(new_n400_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n401_), .A2(KEYINPUT28), .ZN(new_n429_));
  OAI21_X1  g228(.A(KEYINPUT87), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n402_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n417_), .B1(new_n341_), .B2(new_n400_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n433_), .A2(new_n293_), .A3(new_n419_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n415_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n421_), .A2(new_n423_), .A3(new_n425_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n432_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n427_), .A2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G22gat), .B(G50gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G78gat), .B(G106gat), .ZN(new_n441_));
  XOR2_X1   g240(.A(new_n440_), .B(new_n441_), .Z(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n427_), .A2(new_n438_), .A3(new_n442_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n370_), .A2(new_n373_), .ZN(new_n447_));
  AND3_X1   g246(.A1(new_n427_), .A2(new_n442_), .A3(new_n438_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n442_), .B1(new_n427_), .B2(new_n438_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n447_), .B1(new_n448_), .B2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n388_), .A2(KEYINPUT27), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n387_), .A2(new_n291_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n306_), .A2(new_n295_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n203_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n302_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT102), .B1(new_n451_), .B2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT27), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n457_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n301_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT102), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(KEYINPUT27), .A4(new_n388_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n456_), .A2(new_n458_), .A3(new_n461_), .ZN(new_n462_));
  OAI22_X1  g261(.A1(new_n399_), .A2(new_n446_), .B1(new_n450_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G227gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(G71gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT30), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n294_), .B(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n469_), .A2(G99gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n294_), .B(KEYINPUT30), .ZN(new_n471_));
  INV_X1    g270(.A(G99gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G15gat), .B(G43gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT82), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n470_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n476_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n467_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n471_), .A2(new_n472_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n469_), .A2(G99gat), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n475_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n470_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(new_n466_), .A3(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT85), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n479_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n349_), .B(KEYINPUT31), .Z(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n479_), .A2(new_n484_), .A3(new_n485_), .A4(new_n487_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT103), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n492_), .B1(new_n446_), .B2(new_n462_), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n448_), .A2(new_n449_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n458_), .A2(new_n461_), .ZN(new_n495_));
  NAND4_X1  g294(.A1(new_n494_), .A2(new_n495_), .A3(KEYINPUT103), .A4(new_n456_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n370_), .A2(new_n373_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n491_), .A2(new_n498_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n463_), .A2(new_n491_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT13), .ZN(new_n501_));
  NAND2_X1  g300(.A1(G230gat), .A2(G233gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT6), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT6), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n506_), .A2(G99gat), .A3(G106gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(G106gat), .ZN(new_n510_));
  XOR2_X1   g309(.A(KEYINPUT10), .B(G99gat), .Z(new_n511_));
  AOI21_X1  g310(.A(new_n509_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G85gat), .B(G92gat), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n514_), .B(new_n515_), .C1(KEYINPUT9), .C2(G92gat), .ZN(new_n516_));
  INV_X1    g315(.A(new_n515_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(KEYINPUT9), .A2(G92gat), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n513_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n512_), .A2(new_n516_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT8), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT66), .ZN(new_n522_));
  OAI21_X1  g321(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NOR3_X1   g323(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n522_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT7), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(new_n472_), .A3(new_n510_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n528_), .A2(KEYINPUT66), .A3(new_n523_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n526_), .A2(new_n529_), .A3(new_n508_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n521_), .B1(new_n530_), .B2(new_n517_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n528_), .A2(new_n523_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n509_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n521_), .A2(KEYINPUT65), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n521_), .A2(KEYINPUT65), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n517_), .A2(new_n534_), .A3(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(new_n533_), .A2(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n520_), .B1(new_n531_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT67), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G57gat), .B(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT68), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G71gat), .B(G78gat), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n542_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT68), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n541_), .B(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n543_), .A2(new_n544_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT67), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n520_), .B(new_n551_), .C1(new_n531_), .C2(new_n537_), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n539_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n550_), .B1(new_n539_), .B2(new_n552_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n503_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n539_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n556_));
  AND2_X1   g355(.A1(new_n545_), .A2(new_n549_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n557_), .A2(KEYINPUT12), .A3(new_n538_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(KEYINPUT69), .B(KEYINPUT12), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n556_), .B(new_n558_), .C1(new_n554_), .C2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n555_), .B1(new_n561_), .B2(new_n503_), .ZN(new_n562_));
  XOR2_X1   g361(.A(G120gat), .B(G148gat), .Z(new_n563_));
  XNOR2_X1  g362(.A(G176gat), .B(G204gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  XNOR2_X1  g364(.A(KEYINPUT70), .B(KEYINPUT5), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n565_), .B(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n562_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n567_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n555_), .B(new_n569_), .C1(new_n561_), .C2(new_n503_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n568_), .A2(KEYINPUT71), .A3(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT71), .B1(new_n568_), .B2(new_n570_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n501_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT71), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n539_), .A2(new_n552_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n575_), .A2(new_n557_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(new_n559_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n558_), .A2(new_n556_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n577_), .A2(new_n578_), .A3(new_n502_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n569_), .B1(new_n579_), .B2(new_n555_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n570_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n574_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n568_), .A2(KEYINPUT71), .A3(new_n570_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(KEYINPUT13), .A3(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n573_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G15gat), .B(G22gat), .ZN(new_n586_));
  INV_X1    g385(.A(G1gat), .ZN(new_n587_));
  INV_X1    g386(.A(G8gat), .ZN(new_n588_));
  OAI21_X1  g387(.A(KEYINPUT14), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n586_), .A2(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G1gat), .B(G8gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(G29gat), .B(G36gat), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G43gat), .B(G50gat), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(new_n596_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n593_), .A2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n592_), .A2(new_n599_), .A3(new_n598_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G229gat), .A2(G233gat), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n603_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT78), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n600_), .B(KEYINPUT15), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(new_n592_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n609_), .A2(new_n601_), .A3(new_n604_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n610_), .ZN(new_n611_));
  XOR2_X1   g410(.A(G113gat), .B(G141gat), .Z(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT79), .ZN(new_n613_));
  XOR2_X1   g412(.A(G169gat), .B(G197gat), .Z(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n611_), .B(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n585_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n500_), .A2(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(G127gat), .B(G155gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT16), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n620_), .B(new_n621_), .Z(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n550_), .A2(new_n593_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n550_), .A2(new_n593_), .ZN(new_n626_));
  NAND4_X1  g425(.A1(new_n625_), .A2(G231gat), .A3(G233gat), .A4(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628_));
  INV_X1    g427(.A(new_n626_), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n628_), .B1(new_n629_), .B2(new_n624_), .ZN(new_n630_));
  AND2_X1   g429(.A1(new_n627_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT76), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n623_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT17), .B1(new_n631_), .B2(new_n623_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT17), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n635_), .B1(new_n636_), .B2(new_n633_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G190gat), .B(G218gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G134gat), .B(G162gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n638_), .B(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT36), .Z(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT74), .Z(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n538_), .A2(new_n608_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT73), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G232gat), .A2(G233gat), .ZN(new_n646_));
  XOR2_X1   g445(.A(new_n646_), .B(KEYINPUT34), .Z(new_n647_));
  INV_X1    g446(.A(KEYINPUT35), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n645_), .A2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n539_), .A2(new_n600_), .A3(new_n552_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n647_), .A2(new_n648_), .ZN(new_n652_));
  XOR2_X1   g451(.A(new_n652_), .B(KEYINPUT72), .Z(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n608_), .B2(new_n538_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n650_), .B1(new_n651_), .B2(new_n654_), .ZN(new_n655_));
  AOI211_X1 g454(.A(new_n648_), .B(new_n647_), .C1(new_n644_), .C2(KEYINPUT73), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n651_), .A2(new_n654_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n643_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n656_), .A2(new_n657_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n650_), .A2(new_n651_), .A3(new_n654_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n640_), .A2(KEYINPUT36), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n659_), .A2(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(KEYINPUT75), .B(KEYINPUT37), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n659_), .A2(new_n663_), .A3(new_n665_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n637_), .A2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT77), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n618_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(new_n587_), .A3(new_n498_), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT38), .ZN(new_n675_));
  OR2_X1    g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n664_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n500_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n637_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n617_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G1gat), .B1(new_n681_), .B2(new_n447_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n674_), .A2(new_n675_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n676_), .A2(new_n682_), .A3(new_n683_), .ZN(G1324gat));
  NAND3_X1  g483(.A1(new_n673_), .A2(new_n588_), .A3(new_n462_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT39), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n678_), .A2(new_n680_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n462_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n686_), .B1(new_n688_), .B2(G8gat), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT39), .B(new_n588_), .C1(new_n687_), .C2(new_n462_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n685_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n691_), .B(new_n692_), .Z(G1325gat));
  OAI21_X1  g492(.A(G15gat), .B1(new_n681_), .B2(new_n491_), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n694_), .A2(KEYINPUT105), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(KEYINPUT105), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n695_), .A2(KEYINPUT41), .A3(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT41), .B1(new_n695_), .B2(new_n696_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n672_), .A2(G15gat), .A3(new_n491_), .ZN(new_n699_));
  OR3_X1    g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(G1326gat));
  OAI21_X1  g499(.A(G22gat), .B1(new_n681_), .B2(new_n494_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT42), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n494_), .A2(G22gat), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n702_), .B1(new_n672_), .B2(new_n703_), .ZN(G1327gat));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n659_), .A2(new_n663_), .A3(new_n665_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n665_), .B1(new_n659_), .B2(new_n663_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n705_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n667_), .A2(new_n668_), .A3(KEYINPUT107), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n497_), .A2(new_n499_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n378_), .A2(new_n389_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n390_), .A2(KEYINPUT33), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n712_), .A2(new_n398_), .A3(new_n713_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n498_), .B(new_n304_), .C1(new_n303_), .C2(new_n308_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n446_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n450_), .A2(new_n462_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n491_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n710_), .B1(new_n711_), .B2(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n720_));
  OR2_X1    g519(.A1(new_n669_), .A2(KEYINPUT43), .ZN(new_n721_));
  OAI22_X1  g520(.A1(new_n719_), .A2(new_n720_), .B1(new_n500_), .B2(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n617_), .A2(new_n637_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n722_), .A2(KEYINPUT44), .A3(new_n723_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n498_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(G29gat), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n637_), .A2(new_n664_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n618_), .A2(new_n730_), .ZN(new_n731_));
  OR3_X1    g530(.A1(new_n731_), .A2(G29gat), .A3(new_n447_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n729_), .A2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT108), .ZN(G1328gat));
  OR2_X1    g533(.A1(new_n462_), .A2(KEYINPUT109), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n462_), .A2(KEYINPUT109), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n731_), .A2(G36gat), .A3(new_n738_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT45), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n726_), .A2(new_n462_), .A3(new_n727_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G36gat), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n740_), .A2(new_n742_), .A3(KEYINPUT46), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1329gat));
  INV_X1    g546(.A(G43gat), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n491_), .A2(new_n748_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n726_), .A2(new_n727_), .A3(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT110), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n726_), .A2(new_n752_), .A3(new_n727_), .A4(new_n749_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n748_), .B1(new_n731_), .B2(new_n491_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n751_), .A2(new_n753_), .A3(new_n754_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n755_), .B(new_n757_), .ZN(G1330gat));
  NOR2_X1   g557(.A1(new_n731_), .A2(new_n494_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(G50gat), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n726_), .A2(new_n727_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n446_), .A2(G50gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(G1331gat));
  INV_X1    g562(.A(new_n616_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n573_), .A2(new_n764_), .A3(new_n584_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n500_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(new_n671_), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n447_), .B1(new_n767_), .B2(KEYINPUT112), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(KEYINPUT112), .B2(new_n767_), .ZN(new_n769_));
  INV_X1    g568(.A(G57gat), .ZN(new_n770_));
  NOR4_X1   g569(.A1(new_n500_), .A2(new_n679_), .A3(new_n765_), .A4(new_n677_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n447_), .A2(new_n770_), .ZN(new_n772_));
  AOI22_X1  g571(.A1(new_n769_), .A2(new_n770_), .B1(new_n771_), .B2(new_n772_), .ZN(G1332gat));
  INV_X1    g572(.A(G64gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n771_), .B2(new_n737_), .ZN(new_n775_));
  XNOR2_X1  g574(.A(KEYINPUT113), .B(KEYINPUT48), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n775_), .B(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n767_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n774_), .A3(new_n737_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1333gat));
  INV_X1    g579(.A(new_n491_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n465_), .B1(new_n771_), .B2(new_n781_), .ZN(new_n782_));
  XOR2_X1   g581(.A(new_n782_), .B(KEYINPUT49), .Z(new_n783_));
  NAND3_X1  g582(.A1(new_n778_), .A2(new_n465_), .A3(new_n781_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(G1334gat));
  INV_X1    g584(.A(G78gat), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n771_), .B2(new_n446_), .ZN(new_n787_));
  XOR2_X1   g586(.A(new_n787_), .B(KEYINPUT50), .Z(new_n788_));
  NAND3_X1  g587(.A1(new_n778_), .A2(new_n786_), .A3(new_n446_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(G1335gat));
  NOR3_X1   g589(.A1(new_n571_), .A2(new_n572_), .A3(new_n501_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT13), .B1(new_n582_), .B2(new_n583_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n793_), .A2(KEYINPUT114), .A3(new_n764_), .A4(new_n679_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT114), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n795_), .B1(new_n765_), .B2(new_n637_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n722_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n498_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n766_), .A2(new_n730_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n447_), .A2(G85gat), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n799_), .A2(G85gat), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n802_), .B(KEYINPUT115), .Z(G1336gat));
  INV_X1    g602(.A(G92gat), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n800_), .A2(new_n804_), .A3(new_n462_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n798_), .A2(new_n737_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(new_n806_), .B2(new_n804_), .ZN(new_n807_));
  XOR2_X1   g606(.A(new_n807_), .B(KEYINPUT116), .Z(G1337gat));
  NAND3_X1  g607(.A1(new_n722_), .A2(new_n781_), .A3(new_n797_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(G99gat), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT117), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n781_), .A2(new_n511_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n766_), .A2(new_n811_), .A3(new_n730_), .A4(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n711_), .A2(new_n718_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n765_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n730_), .A4(new_n812_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT117), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n813_), .A2(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n810_), .A2(KEYINPUT119), .A3(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT118), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT51), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n810_), .A2(KEYINPUT118), .A3(new_n818_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT51), .ZN(new_n824_));
  AOI22_X1  g623(.A1(new_n809_), .A2(G99gat), .B1(new_n817_), .B2(new_n813_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT118), .B1(new_n825_), .B2(KEYINPUT119), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n822_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT120), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n822_), .B(new_n829_), .C1(new_n824_), .C2(new_n826_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(G1338gat));
  NAND3_X1  g630(.A1(new_n800_), .A2(new_n510_), .A3(new_n446_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n722_), .A2(new_n446_), .A3(new_n797_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT52), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n833_), .A2(new_n834_), .A3(G106gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n834_), .B1(new_n833_), .B2(G106gat), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n832_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g637(.A1(new_n616_), .A2(new_n570_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n561_), .B2(new_n503_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n561_), .A2(new_n503_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n567_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT56), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n843_), .A2(KEYINPUT56), .A3(new_n567_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n839_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  OR2_X1    g647(.A1(new_n611_), .A2(new_n615_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n609_), .A2(new_n601_), .A3(new_n605_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n603_), .A2(new_n604_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n850_), .A2(new_n615_), .A3(new_n851_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n849_), .A2(new_n852_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n853_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n664_), .B1(new_n848_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n853_), .A2(new_n570_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n847_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT56), .B1(new_n843_), .B2(new_n567_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n858_), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT58), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n669_), .ZN(new_n864_));
  OAI211_X1 g663(.A(KEYINPUT58), .B(new_n858_), .C1(new_n859_), .C2(new_n860_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n863_), .A2(new_n864_), .A3(new_n865_), .ZN(new_n866_));
  OAI211_X1 g665(.A(KEYINPUT57), .B(new_n664_), .C1(new_n848_), .C2(new_n854_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n857_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n670_), .A2(new_n616_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n585_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT121), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n869_), .B(new_n585_), .C1(KEYINPUT121), .C2(KEYINPUT54), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(KEYINPUT121), .A2(KEYINPUT54), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n868_), .A2(new_n679_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n497_), .A2(new_n498_), .A3(new_n781_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(G113gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(new_n880_), .A3(new_n616_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n868_), .A2(new_n679_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n875_), .A2(new_n876_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n878_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(KEYINPUT59), .A3(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT59), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n887_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n764_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n881_), .B1(new_n889_), .B2(new_n880_), .ZN(G1340gat));
  AOI21_X1  g689(.A(new_n585_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n891_));
  INV_X1    g690(.A(G120gat), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n585_), .A2(KEYINPUT60), .ZN(new_n894_));
  MUX2_X1   g693(.A(KEYINPUT60), .B(new_n894_), .S(new_n892_), .Z(new_n895_));
  AND3_X1   g694(.A1(new_n879_), .A2(new_n893_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n893_), .B1(new_n879_), .B2(new_n895_), .ZN(new_n897_));
  OAI22_X1  g696(.A1(new_n891_), .A2(new_n892_), .B1(new_n896_), .B2(new_n897_), .ZN(G1341gat));
  INV_X1    g697(.A(G127gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n879_), .A2(new_n899_), .A3(new_n637_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n679_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n899_), .ZN(G1342gat));
  INV_X1    g701(.A(G134gat), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n879_), .A2(new_n903_), .A3(new_n677_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n669_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n904_), .B1(new_n905_), .B2(new_n903_), .ZN(G1343gat));
  NOR2_X1   g705(.A1(new_n877_), .A2(new_n781_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n494_), .A2(new_n447_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n738_), .A2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n907_), .A2(new_n616_), .A3(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g711(.A1(new_n907_), .A2(new_n793_), .A3(new_n910_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g713(.A1(new_n907_), .A2(new_n637_), .A3(new_n910_), .ZN(new_n915_));
  XNOR2_X1  g714(.A(KEYINPUT61), .B(G155gat), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n915_), .B(new_n916_), .ZN(G1346gat));
  INV_X1    g716(.A(G162gat), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n710_), .A2(new_n918_), .ZN(new_n919_));
  AND3_X1   g718(.A1(new_n907_), .A2(new_n910_), .A3(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT123), .ZN(new_n921_));
  NOR4_X1   g720(.A1(new_n877_), .A2(new_n781_), .A3(new_n664_), .A4(new_n909_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n921_), .B1(new_n922_), .B2(G162gat), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n884_), .A2(new_n491_), .A3(new_n677_), .A4(new_n910_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n924_), .A2(KEYINPUT123), .A3(new_n918_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n920_), .B1(new_n923_), .B2(new_n925_), .ZN(G1347gat));
  AND3_X1   g725(.A1(new_n737_), .A2(new_n494_), .A3(new_n499_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n884_), .A2(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(G169gat), .B1(new_n928_), .B2(new_n764_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n928_), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n932_), .B(new_n616_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n930_), .ZN(new_n934_));
  OAI211_X1 g733(.A(G169gat), .B(new_n934_), .C1(new_n928_), .C2(new_n764_), .ZN(new_n935_));
  NAND3_X1  g734(.A1(new_n931_), .A2(new_n933_), .A3(new_n935_), .ZN(G1348gat));
  NOR2_X1   g735(.A1(new_n928_), .A2(new_n585_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(new_n250_), .ZN(G1349gat));
  NOR3_X1   g737(.A1(new_n928_), .A2(new_n266_), .A3(new_n679_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n932_), .A2(new_n637_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n939_), .B1(new_n271_), .B2(new_n940_), .ZN(G1350gat));
  OAI21_X1  g740(.A(G190gat), .B1(new_n928_), .B2(new_n669_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n677_), .A2(new_n267_), .ZN(new_n943_));
  XOR2_X1   g742(.A(new_n943_), .B(KEYINPUT125), .Z(new_n944_));
  OAI21_X1  g743(.A(new_n942_), .B1(new_n928_), .B2(new_n944_), .ZN(G1351gat));
  NOR2_X1   g744(.A1(new_n738_), .A2(new_n450_), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n907_), .A2(new_n616_), .A3(new_n946_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(G197gat), .ZN(G1352gat));
  NOR4_X1   g747(.A1(new_n877_), .A2(new_n450_), .A3(new_n781_), .A4(new_n738_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(KEYINPUT126), .A2(G204gat), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n949_), .A2(new_n793_), .A3(new_n950_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n907_), .A2(new_n946_), .ZN(new_n952_));
  NOR2_X1   g751(.A1(new_n952_), .A2(new_n585_), .ZN(new_n953_));
  XOR2_X1   g752(.A(KEYINPUT126), .B(G204gat), .Z(new_n954_));
  OAI21_X1  g753(.A(new_n951_), .B1(new_n953_), .B2(new_n954_), .ZN(G1353gat));
  INV_X1    g754(.A(KEYINPUT63), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(new_n222_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n637_), .B1(new_n956_), .B2(new_n222_), .ZN(new_n958_));
  XNOR2_X1  g757(.A(new_n958_), .B(KEYINPUT127), .ZN(new_n959_));
  AOI21_X1  g758(.A(new_n957_), .B1(new_n949_), .B2(new_n959_), .ZN(new_n960_));
  AND4_X1   g759(.A1(new_n907_), .A2(new_n946_), .A3(new_n957_), .A4(new_n959_), .ZN(new_n961_));
  NOR2_X1   g760(.A1(new_n960_), .A2(new_n961_), .ZN(G1354gat));
  OAI21_X1  g761(.A(G218gat), .B1(new_n952_), .B2(new_n669_), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n949_), .A2(new_n224_), .A3(new_n677_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n963_), .A2(new_n964_), .ZN(G1355gat));
endmodule


