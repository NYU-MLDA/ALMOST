//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 1 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:03 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n911_,
    new_n912_, new_n913_, new_n914_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_;
  NAND2_X1  g000(.A1(G141gat), .A2(G148gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND3_X1  g003(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n205_));
  OR2_X1    g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  OAI211_X1 g005(.A(new_n204_), .B(new_n205_), .C1(new_n206_), .C2(KEYINPUT3), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT87), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  NOR2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT85), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n211_), .A2(new_n214_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n215_), .B(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n214_), .A2(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n206_), .A2(new_n202_), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n219_), .A2(KEYINPUT86), .A3(new_n220_), .ZN(new_n221_));
  AOI21_X1  g020(.A(KEYINPUT86), .B1(new_n219_), .B2(new_n220_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n216_), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT28), .B1(new_n223_), .B2(KEYINPUT29), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n214_), .A2(new_n215_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n225_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n219_), .A2(new_n220_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT86), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n219_), .A2(KEYINPUT86), .A3(new_n220_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n226_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT28), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT29), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G22gat), .B(G50gat), .ZN(new_n235_));
  AND3_X1   g034(.A1(new_n224_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n235_), .B1(new_n224_), .B2(new_n234_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G78gat), .B(G106gat), .ZN(new_n240_));
  INV_X1    g039(.A(G233gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT88), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n242_), .A2(G228gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(G228gat), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n241_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n223_), .A2(KEYINPUT29), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G197gat), .B(G204gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G211gat), .B(G218gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n250_), .A2(new_n252_), .A3(KEYINPUT21), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n251_), .B1(new_n250_), .B2(KEYINPUT21), .ZN(new_n254_));
  INV_X1    g053(.A(G197gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT89), .A3(G204gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT21), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT89), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n257_), .B1(new_n258_), .B2(new_n249_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n253_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n247_), .B1(new_n248_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n260_), .ZN(new_n262_));
  AOI211_X1 g061(.A(new_n262_), .B(new_n246_), .C1(new_n223_), .C2(KEYINPUT29), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n240_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT91), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n260_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n246_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n248_), .A2(new_n260_), .A3(new_n247_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n240_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n268_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(KEYINPUT90), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT91), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n272_), .B(new_n240_), .C1(new_n261_), .C2(new_n263_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT90), .ZN(new_n274_));
  NAND4_X1  g073(.A1(new_n267_), .A2(new_n268_), .A3(new_n274_), .A4(new_n269_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n265_), .A2(new_n271_), .A3(new_n273_), .A4(new_n275_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n267_), .A2(new_n268_), .A3(KEYINPUT92), .A4(new_n269_), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n238_), .A2(new_n264_), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT92), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n270_), .A2(new_n279_), .ZN(new_n280_));
  AOI22_X1  g079(.A1(new_n239_), .A2(new_n276_), .B1(new_n278_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT27), .ZN(new_n282_));
  NAND2_X1  g081(.A1(G226gat), .A2(G233gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT19), .ZN(new_n284_));
  XOR2_X1   g083(.A(KEYINPUT77), .B(G183gat), .Z(new_n285_));
  OR2_X1    g084(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n285_), .A2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT80), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT80), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n293_), .A2(G183gat), .A3(G190gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n290_), .B1(new_n295_), .B2(KEYINPUT23), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT81), .ZN(new_n297_));
  AOI21_X1  g096(.A(G176gat), .B1(new_n297_), .B2(KEYINPUT22), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n298_), .A2(G169gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(G169gat), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n289_), .A2(new_n296_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(KEYINPUT23), .B1(new_n292_), .B2(new_n294_), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n291_), .A2(KEYINPUT23), .ZN(new_n303_));
  INV_X1    g102(.A(G169gat), .ZN(new_n304_));
  INV_X1    g103(.A(G176gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OAI22_X1  g105(.A1(new_n302_), .A2(new_n303_), .B1(KEYINPUT24), .B2(new_n306_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n286_), .A2(KEYINPUT26), .A3(new_n287_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT25), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT26), .ZN(new_n310_));
  AOI22_X1  g109(.A1(new_n309_), .A2(G183gat), .B1(new_n310_), .B2(G190gat), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n308_), .B(new_n311_), .C1(new_n285_), .C2(new_n309_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G169gat), .A2(G176gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n306_), .A2(KEYINPUT24), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT79), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n307_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(KEYINPUT79), .A3(new_n314_), .ZN(new_n318_));
  AOI211_X1 g117(.A(new_n260_), .B(new_n301_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n319_));
  OAI22_X1  g118(.A1(new_n302_), .A2(new_n303_), .B1(G183gat), .B2(G190gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT22), .B(G169gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(new_n305_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n320_), .A2(new_n313_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n306_), .A2(new_n313_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT93), .B(KEYINPUT24), .ZN(new_n325_));
  OR2_X1    g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT25), .B(G183gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT26), .B(G190gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n325_), .A2(new_n304_), .A3(new_n305_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n326_), .A2(new_n296_), .A3(new_n329_), .A4(new_n330_), .ZN(new_n331_));
  AND2_X1   g130(.A1(new_n323_), .A2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT20), .B1(new_n332_), .B2(new_n262_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n284_), .B1(new_n319_), .B2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT20), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n335_), .B1(new_n332_), .B2(new_n262_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n284_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n301_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n336_), .B(new_n337_), .C1(new_n262_), .C2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(G8gat), .B(G36gat), .Z(new_n340_));
  XNOR2_X1  g139(.A(G64gat), .B(G92gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n342_), .B(new_n343_), .Z(new_n344_));
  AND3_X1   g143(.A1(new_n334_), .A2(new_n339_), .A3(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n344_), .B1(new_n334_), .B2(new_n339_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n282_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(new_n344_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n315_), .A2(new_n316_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n307_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n318_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n301_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n260_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n337_), .B1(new_n354_), .B2(new_n336_), .ZN(new_n355_));
  NOR3_X1   g154(.A1(new_n319_), .A2(new_n333_), .A3(new_n284_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n348_), .B1(new_n355_), .B2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n334_), .A2(new_n339_), .A3(new_n344_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(KEYINPUT27), .A3(new_n358_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n347_), .A2(new_n359_), .A3(KEYINPUT99), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT99), .B1(new_n347_), .B2(new_n359_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n281_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(KEYINPUT100), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT100), .ZN(new_n364_));
  OAI211_X1 g163(.A(new_n281_), .B(new_n364_), .C1(new_n360_), .C2(new_n361_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n363_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G227gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G71gat), .ZN(new_n368_));
  INV_X1    g167(.A(G99gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n368_), .B(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n353_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G15gat), .B(G43gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT82), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT30), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n338_), .B(new_n370_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n374_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  XOR2_X1   g177(.A(G127gat), .B(G134gat), .Z(new_n379_));
  XOR2_X1   g178(.A(G113gat), .B(G120gat), .Z(new_n380_));
  XOR2_X1   g179(.A(new_n379_), .B(new_n380_), .Z(new_n381_));
  XOR2_X1   g180(.A(new_n381_), .B(KEYINPUT31), .Z(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT83), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n375_), .A2(new_n378_), .A3(new_n383_), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n384_), .A2(KEYINPUT84), .ZN(new_n385_));
  AND2_X1   g184(.A1(new_n375_), .A2(new_n378_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n386_), .A2(new_n382_), .ZN(new_n387_));
  AND2_X1   g186(.A1(new_n384_), .A2(KEYINPUT84), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n385_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n223_), .A2(new_n381_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n381_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n391_), .B(new_n216_), .C1(new_n222_), .C2(new_n221_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(KEYINPUT4), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G225gat), .A2(G233gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT4), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n223_), .A2(new_n396_), .A3(new_n381_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n393_), .A2(new_n395_), .A3(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n390_), .A2(new_n394_), .A3(new_n392_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT95), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT95), .ZN(new_n401_));
  NAND4_X1  g200(.A1(new_n390_), .A2(new_n392_), .A3(new_n401_), .A4(new_n394_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n398_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G1gat), .B(G29gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n404_), .B(G85gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(KEYINPUT0), .B(G57gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n403_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n407_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n398_), .A2(new_n400_), .A3(new_n409_), .A4(new_n402_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n408_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n389_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n366_), .A2(new_n414_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n400_), .A2(new_n402_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT96), .ZN(new_n417_));
  NOR2_X1   g216(.A1(new_n417_), .A2(KEYINPUT33), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n416_), .A2(new_n409_), .A3(new_n398_), .A4(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n410_), .A2(new_n418_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n393_), .A2(new_n394_), .A3(new_n397_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n390_), .A2(new_n395_), .A3(new_n392_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n407_), .ZN(new_n425_));
  OAI21_X1  g224(.A(KEYINPUT97), .B1(new_n423_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n346_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n393_), .A2(new_n394_), .A3(new_n397_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT97), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n428_), .A2(new_n429_), .A3(new_n407_), .A4(new_n424_), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n426_), .A2(new_n427_), .A3(new_n358_), .A4(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n422_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n344_), .A2(KEYINPUT32), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n355_), .A2(new_n356_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n334_), .A2(new_n339_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n434_), .B1(KEYINPUT98), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT98), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n433_), .B1(new_n435_), .B2(new_n437_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n436_), .A2(new_n438_), .B1(new_n410_), .B2(new_n408_), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n281_), .B1(new_n432_), .B2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n276_), .A2(new_n239_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n278_), .A2(new_n280_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n347_), .A2(new_n359_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(new_n412_), .A3(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n389_), .B1(new_n440_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n415_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(G36gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(G29gat), .ZN(new_n450_));
  INV_X1    g249(.A(G29gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G36gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(KEYINPUT69), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n450_), .A2(new_n452_), .A3(KEYINPUT69), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G43gat), .B(G50gat), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n456_), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n450_), .A2(new_n452_), .A3(KEYINPUT69), .ZN(new_n459_));
  OAI21_X1  g258(.A(new_n458_), .B1(new_n459_), .B2(new_n453_), .ZN(new_n460_));
  XOR2_X1   g259(.A(KEYINPUT70), .B(KEYINPUT15), .Z(new_n461_));
  AND3_X1   g260(.A1(new_n457_), .A2(new_n460_), .A3(new_n461_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n461_), .B1(new_n457_), .B2(new_n460_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G15gat), .B(G22gat), .ZN(new_n465_));
  INV_X1    g264(.A(G8gat), .ZN(new_n466_));
  OR2_X1    g265(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n467_));
  NAND2_X1  g266(.A1(KEYINPUT74), .A2(G1gat), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n466_), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT14), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n465_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G1gat), .B(G8gat), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n471_), .A2(new_n473_), .ZN(new_n474_));
  OAI211_X1 g273(.A(new_n465_), .B(new_n472_), .C1(new_n469_), .C2(new_n470_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n464_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G229gat), .A2(G233gat), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n457_), .A2(new_n460_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(new_n476_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n479_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT76), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n457_), .A2(new_n460_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(new_n475_), .A3(new_n474_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n481_), .A2(new_n483_), .A3(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n479_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n477_), .A2(KEYINPUT76), .A3(new_n484_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n486_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n482_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G113gat), .B(G141gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G169gat), .B(G197gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n482_), .A2(new_n489_), .A3(new_n493_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n448_), .A2(KEYINPUT101), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT101), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n446_), .B1(new_n366_), .B2(new_n414_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n497_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n499_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n498_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT37), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G190gat), .B(G218gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G134gat), .B(G162gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(new_n507_), .B(KEYINPUT36), .Z(new_n508_));
  NAND2_X1  g307(.A1(G232gat), .A2(G233gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(KEYINPUT34), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT35), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT6), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  OR2_X1    g318(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n520_));
  INV_X1    g319(.A(G106gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(G85gat), .ZN(new_n524_));
  INV_X1    g323(.A(G92gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G85gat), .A2(G92gat), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n526_), .A2(KEYINPUT9), .A3(new_n527_), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n527_), .A2(KEYINPUT9), .ZN(new_n529_));
  NAND4_X1  g328(.A1(new_n519_), .A2(new_n523_), .A3(new_n528_), .A4(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n526_), .A2(new_n527_), .ZN(new_n531_));
  OAI21_X1  g330(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  AOI211_X1 g334(.A(KEYINPUT8), .B(new_n531_), .C1(new_n535_), .C2(new_n519_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT8), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT7), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(new_n369_), .A3(new_n521_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n517_), .B1(G99gat), .B2(G106gat), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n515_), .A2(KEYINPUT6), .ZN(new_n541_));
  OAI211_X1 g340(.A(new_n532_), .B(new_n539_), .C1(new_n540_), .C2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n531_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n537_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n530_), .B1(new_n536_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT66), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(KEYINPUT66), .B(new_n530_), .C1(new_n536_), .C2(new_n544_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n464_), .A3(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT71), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT71), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n547_), .A2(new_n464_), .A3(new_n551_), .A4(new_n548_), .ZN(new_n552_));
  OAI22_X1  g351(.A1(new_n545_), .A2(new_n484_), .B1(KEYINPUT35), .B2(new_n510_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AND4_X1   g353(.A1(new_n514_), .A2(new_n550_), .A3(new_n552_), .A4(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n553_), .B1(new_n549_), .B2(KEYINPUT71), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n514_), .B1(new_n556_), .B2(new_n552_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n508_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n550_), .A2(new_n552_), .A3(new_n554_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n513_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n507_), .A2(KEYINPUT36), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n556_), .A2(new_n514_), .A3(new_n552_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n504_), .B1(new_n558_), .B2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT72), .B1(new_n555_), .B2(new_n557_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT72), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n560_), .A2(new_n566_), .A3(new_n562_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n565_), .A2(new_n567_), .A3(new_n508_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(new_n504_), .A3(new_n563_), .ZN(new_n569_));
  INV_X1    g368(.A(KEYINPUT73), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n568_), .A2(KEYINPUT73), .A3(new_n504_), .A4(new_n563_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n564_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G231gat), .A2(G233gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT75), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n476_), .B(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G57gat), .B(G64gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT11), .ZN(new_n578_));
  XOR2_X1   g377(.A(G71gat), .B(G78gat), .Z(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n579_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n577_), .A2(KEYINPUT11), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n581_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n576_), .B(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G127gat), .B(G155gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT16), .ZN(new_n587_));
  XOR2_X1   g386(.A(G183gat), .B(G211gat), .Z(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT17), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n585_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT17), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n589_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n591_), .B1(new_n594_), .B2(new_n585_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n573_), .A2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT67), .ZN(new_n597_));
  INV_X1    g396(.A(new_n530_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n542_), .A2(new_n543_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT8), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n542_), .A2(new_n537_), .A3(new_n543_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n598_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT65), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n602_), .A2(new_n603_), .A3(new_n584_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n582_), .A2(new_n583_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(new_n580_), .ZN(new_n606_));
  OAI21_X1  g405(.A(KEYINPUT65), .B1(new_n545_), .B2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n545_), .A2(new_n606_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n604_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(G230gat), .A2(G233gat), .ZN(new_n610_));
  XOR2_X1   g409(.A(new_n610_), .B(KEYINPUT64), .Z(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n581_), .B(KEYINPUT12), .C1(new_n583_), .C2(new_n582_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n547_), .A2(new_n548_), .A3(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT12), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n602_), .B2(new_n584_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n611_), .B1(new_n602_), .B2(new_n584_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G120gat), .B(G148gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT5), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G176gat), .B(G204gat), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n621_), .B(new_n622_), .Z(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n612_), .A2(new_n619_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n624_), .B1(new_n612_), .B2(new_n619_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n597_), .B1(new_n626_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR3_X1   g428(.A1(new_n626_), .A2(new_n597_), .A3(new_n627_), .ZN(new_n630_));
  OAI22_X1  g429(.A1(new_n629_), .A2(new_n630_), .B1(KEYINPUT68), .B2(KEYINPUT13), .ZN(new_n631_));
  OR3_X1    g430(.A1(new_n626_), .A2(new_n597_), .A3(new_n627_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n632_), .A2(new_n628_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n631_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n596_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n503_), .A2(KEYINPUT102), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(KEYINPUT102), .B1(new_n503_), .B2(new_n637_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n411_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n642_));
  XOR2_X1   g441(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n643_));
  NAND3_X1  g442(.A1(new_n641_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n635_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n645_), .A2(new_n501_), .A3(new_n595_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n568_), .A2(new_n563_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n448_), .A2(new_n646_), .A3(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(G1gat), .B1(new_n649_), .B2(new_n412_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n644_), .A2(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n643_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1324gat));
  NOR2_X1   g452(.A1(new_n360_), .A2(new_n361_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n641_), .A2(new_n466_), .A3(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n500_), .A2(new_n647_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n657_), .A2(new_n654_), .A3(new_n646_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n656_), .B1(new_n658_), .B2(G8gat), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  AOI211_X1 g460(.A(KEYINPUT104), .B(new_n656_), .C1(new_n658_), .C2(G8gat), .ZN(new_n662_));
  OR2_X1    g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n658_), .A2(new_n656_), .A3(G8gat), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT105), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n658_), .A2(KEYINPUT105), .A3(new_n656_), .A4(G8gat), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n655_), .B(KEYINPUT40), .C1(new_n663_), .C2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n668_), .A2(new_n662_), .A3(new_n661_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n654_), .ZN(new_n672_));
  NOR4_X1   g471(.A1(new_n639_), .A2(new_n640_), .A3(G8gat), .A4(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n669_), .A2(new_n674_), .ZN(G1325gat));
  INV_X1    g474(.A(new_n389_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G15gat), .B1(new_n649_), .B2(new_n676_), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT41), .Z(new_n678_));
  INV_X1    g477(.A(new_n641_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n676_), .A2(G15gat), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(G1326gat));
  OAI21_X1  g480(.A(G22gat), .B1(new_n649_), .B2(new_n281_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT42), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n281_), .A2(G22gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n679_), .B2(new_n684_), .ZN(G1327gat));
  INV_X1    g484(.A(new_n595_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n648_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n635_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n498_), .B2(new_n502_), .ZN(new_n689_));
  AOI21_X1  g488(.A(G29gat), .B1(new_n689_), .B2(new_n411_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n635_), .A2(new_n497_), .A3(new_n595_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n573_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT43), .B1(new_n500_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n413_), .B1(new_n363_), .B2(new_n365_), .ZN(new_n695_));
  OAI211_X1 g494(.A(new_n694_), .B(new_n573_), .C1(new_n695_), .C2(new_n446_), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n691_), .B1(new_n693_), .B2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT44), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n693_), .A2(new_n696_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n691_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT107), .ZN(new_n703_));
  XOR2_X1   g502(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n702_), .A2(new_n703_), .A3(new_n705_), .ZN(new_n706_));
  OAI21_X1  g505(.A(KEYINPUT107), .B1(new_n697_), .B2(new_n704_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n699_), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n412_), .A2(new_n451_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n690_), .B1(new_n708_), .B2(new_n709_), .ZN(G1328gat));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n672_), .A2(G36gat), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n689_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n711_), .B1(new_n689_), .B2(new_n712_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n698_), .A2(new_n654_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n707_), .B2(new_n706_), .ZN(new_n716_));
  OAI221_X1 g515(.A(KEYINPUT46), .B1(new_n713_), .B2(new_n714_), .C1(new_n716_), .C2(new_n449_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT46), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n706_), .A2(new_n707_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n715_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n449_), .B1(new_n719_), .B2(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n713_), .A2(new_n714_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n717_), .A2(new_n723_), .ZN(G1329gat));
  NAND4_X1  g523(.A1(new_n719_), .A2(G43gat), .A3(new_n389_), .A4(new_n698_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n689_), .A2(new_n389_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n726_), .A2(G43gat), .ZN(new_n727_));
  XNOR2_X1  g526(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n725_), .A2(new_n727_), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n725_), .B2(new_n727_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1330gat));
  AOI21_X1  g530(.A(G50gat), .B1(new_n689_), .B2(new_n443_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n443_), .A2(G50gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n732_), .B1(new_n708_), .B2(new_n733_), .ZN(G1331gat));
  NAND4_X1  g533(.A1(new_n657_), .A2(new_n501_), .A3(new_n645_), .A4(new_n686_), .ZN(new_n735_));
  INV_X1    g534(.A(G57gat), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(new_n412_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n500_), .A2(new_n497_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n738_), .A2(new_n645_), .A3(new_n596_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  OR2_X1    g539(.A1(new_n740_), .A2(KEYINPUT109), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(KEYINPUT109), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n411_), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n737_), .B1(new_n743_), .B2(new_n736_), .ZN(G1332gat));
  OAI21_X1  g543(.A(G64gat), .B1(new_n735_), .B2(new_n672_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(KEYINPUT48), .ZN(new_n746_));
  OR2_X1    g545(.A1(new_n672_), .A2(G64gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n739_), .B2(new_n747_), .ZN(G1333gat));
  OAI21_X1  g547(.A(G71gat), .B1(new_n735_), .B2(new_n676_), .ZN(new_n749_));
  XOR2_X1   g548(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n750_));
  XNOR2_X1  g549(.A(new_n749_), .B(new_n750_), .ZN(new_n751_));
  OR2_X1    g550(.A1(new_n676_), .A2(G71gat), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n751_), .B1(new_n739_), .B2(new_n752_), .ZN(G1334gat));
  OAI21_X1  g552(.A(G78gat), .B1(new_n735_), .B2(new_n281_), .ZN(new_n754_));
  XOR2_X1   g553(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n755_));
  XNOR2_X1  g554(.A(new_n754_), .B(new_n755_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n281_), .A2(G78gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n739_), .B2(new_n757_), .ZN(G1335gat));
  NAND3_X1  g557(.A1(new_n645_), .A2(new_n501_), .A3(new_n595_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n759_), .B1(new_n693_), .B2(new_n696_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n760_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n412_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n738_), .A2(new_n645_), .A3(new_n687_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n524_), .A3(new_n411_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(G1336gat));
  OAI21_X1  g565(.A(G92gat), .B1(new_n761_), .B2(new_n672_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n525_), .A3(new_n654_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1337gat));
  OAI21_X1  g568(.A(G99gat), .B1(new_n761_), .B2(new_n676_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n389_), .A2(new_n520_), .A3(new_n522_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n763_), .B2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g572(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT112), .ZN(new_n775_));
  INV_X1    g574(.A(new_n759_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n700_), .A2(new_n775_), .A3(new_n443_), .A4(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(G106gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n775_), .B1(new_n760_), .B2(new_n443_), .ZN(new_n779_));
  OAI21_X1  g578(.A(KEYINPUT52), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n700_), .A2(new_n443_), .A3(new_n776_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT112), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT52), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n782_), .A2(new_n783_), .A3(G106gat), .A4(new_n777_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n780_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n443_), .A2(new_n521_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n763_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n774_), .B1(new_n785_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n774_), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n787_), .B(new_n790_), .C1(new_n780_), .C2(new_n784_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1339gat));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793_));
  INV_X1    g592(.A(new_n496_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n493_), .B1(new_n482_), .B2(new_n489_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n625_), .B(new_n793_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n793_), .B1(new_n497_), .B2(new_n625_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n615_), .A2(new_n607_), .A3(new_n604_), .A4(new_n617_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n611_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT116), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(KEYINPUT116), .A3(new_n611_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT55), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n619_), .A2(new_n805_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n615_), .A2(KEYINPUT55), .A3(new_n617_), .A4(new_n618_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n803_), .A2(new_n804_), .A3(new_n806_), .A4(new_n807_), .ZN(new_n808_));
  AND3_X1   g607(.A1(new_n808_), .A2(KEYINPUT56), .A3(new_n623_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT56), .B1(new_n808_), .B2(new_n623_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n799_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n478_), .A2(new_n487_), .A3(new_n481_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n486_), .A2(new_n479_), .A3(new_n488_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n813_), .A3(new_n494_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n496_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n632_), .B2(new_n628_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n647_), .B1(new_n811_), .B2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT57), .B1(new_n818_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  INV_X1    g621(.A(new_n804_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n806_), .A2(new_n807_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT116), .B1(new_n800_), .B2(new_n611_), .ZN(new_n825_));
  NOR3_X1   g624(.A1(new_n823_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n822_), .B1(new_n826_), .B2(new_n624_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n808_), .A2(KEYINPUT56), .A3(new_n623_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n816_), .B1(new_n829_), .B2(new_n799_), .ZN(new_n830_));
  OAI211_X1 g629(.A(KEYINPUT117), .B(new_n821_), .C1(new_n830_), .C2(new_n647_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n626_), .A2(new_n815_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n832_), .B1(new_n809_), .B2(new_n810_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT58), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n829_), .A2(KEYINPUT58), .A3(new_n832_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n573_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n820_), .A2(new_n831_), .A3(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n839_));
  AOI211_X1 g638(.A(new_n497_), .B(new_n595_), .C1(new_n839_), .C2(KEYINPUT54), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n635_), .A2(new_n840_), .ZN(new_n841_));
  OAI22_X1  g640(.A1(new_n573_), .A2(new_n841_), .B1(new_n839_), .B2(KEYINPUT54), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n839_), .A2(KEYINPUT54), .ZN(new_n843_));
  INV_X1    g642(.A(new_n841_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n692_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n838_), .A2(new_n595_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n366_), .A2(new_n389_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n412_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT118), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(KEYINPUT59), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n852_));
  NOR4_X1   g651(.A1(new_n846_), .A2(new_n847_), .A3(new_n412_), .A4(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(KEYINPUT119), .B1(new_n851_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n852_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n848_), .A2(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT119), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n856_), .B(new_n857_), .C1(new_n848_), .C2(new_n850_), .ZN(new_n858_));
  AND4_X1   g657(.A1(G113gat), .A2(new_n854_), .A3(new_n858_), .A4(new_n497_), .ZN(new_n859_));
  AOI21_X1  g658(.A(G113gat), .B1(new_n848_), .B2(new_n497_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1340gat));
  NOR3_X1   g660(.A1(new_n851_), .A2(new_n635_), .A3(new_n853_), .ZN(new_n862_));
  INV_X1    g661(.A(G120gat), .ZN(new_n863_));
  INV_X1    g662(.A(new_n848_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT120), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n863_), .B2(KEYINPUT60), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n863_), .B1(new_n635_), .B2(KEYINPUT60), .ZN(new_n867_));
  MUX2_X1   g666(.A(new_n865_), .B(new_n866_), .S(new_n867_), .Z(new_n868_));
  OAI22_X1  g667(.A1(new_n862_), .A2(new_n863_), .B1(new_n864_), .B2(new_n868_), .ZN(G1341gat));
  AND4_X1   g668(.A1(G127gat), .A2(new_n854_), .A3(new_n858_), .A4(new_n686_), .ZN(new_n870_));
  AOI21_X1  g669(.A(G127gat), .B1(new_n848_), .B2(new_n686_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1342gat));
  XOR2_X1   g671(.A(KEYINPUT121), .B(G134gat), .Z(new_n873_));
  AND4_X1   g672(.A1(new_n573_), .A2(new_n854_), .A3(new_n858_), .A4(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(G134gat), .B1(new_n848_), .B2(new_n647_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1343gat));
  NAND2_X1  g675(.A1(new_n838_), .A2(new_n595_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n845_), .A2(new_n842_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n412_), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n654_), .A2(new_n389_), .A3(new_n281_), .ZN(new_n880_));
  AOI21_X1  g679(.A(KEYINPUT122), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n882_));
  INV_X1    g681(.A(new_n880_), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n846_), .A2(new_n882_), .A3(new_n412_), .A4(new_n883_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n881_), .A2(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n497_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n645_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT123), .B(G148gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1345gat));
  OAI21_X1  g689(.A(new_n686_), .B1(new_n881_), .B2(new_n884_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT124), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n893_), .B(new_n686_), .C1(new_n881_), .C2(new_n884_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(KEYINPUT61), .B(G155gat), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n892_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n892_), .B2(new_n894_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1346gat));
  INV_X1    g697(.A(G162gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n885_), .A2(new_n899_), .A3(new_n647_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n885_), .A2(new_n573_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n900_), .B1(new_n901_), .B2(new_n899_), .ZN(G1347gat));
  NOR4_X1   g701(.A1(new_n846_), .A2(new_n443_), .A3(new_n672_), .A4(new_n413_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n304_), .B1(new_n903_), .B2(new_n497_), .ZN(new_n904_));
  OR2_X1    g703(.A1(new_n904_), .A2(KEYINPUT62), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n903_), .A2(new_n321_), .A3(new_n497_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n904_), .A2(KEYINPUT62), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n905_), .A2(new_n906_), .A3(new_n907_), .ZN(G1348gat));
  NAND2_X1  g707(.A1(new_n903_), .A2(new_n645_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g709(.A1(new_n903_), .A2(new_n686_), .ZN(new_n911_));
  OR3_X1    g710(.A1(new_n911_), .A2(KEYINPUT125), .A3(new_n327_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n285_), .B1(new_n903_), .B2(new_n686_), .ZN(new_n913_));
  OAI21_X1  g712(.A(KEYINPUT125), .B1(new_n911_), .B2(new_n327_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(G1350gat));
  NAND3_X1  g714(.A1(new_n903_), .A2(new_n328_), .A3(new_n647_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n903_), .A2(new_n573_), .ZN(new_n917_));
  INV_X1    g716(.A(G190gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n916_), .B1(new_n917_), .B2(new_n918_), .ZN(G1351gat));
  NAND2_X1  g718(.A1(new_n877_), .A2(new_n878_), .ZN(new_n920_));
  NOR4_X1   g719(.A1(new_n672_), .A2(new_n389_), .A3(new_n411_), .A4(new_n281_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n920_), .A2(new_n921_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n922_), .A2(new_n501_), .ZN(new_n923_));
  XNOR2_X1  g722(.A(new_n923_), .B(new_n255_), .ZN(G1352gat));
  INV_X1    g723(.A(new_n922_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n645_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(G204gat), .ZN(G1353gat));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n928_), .B1(new_n925_), .B2(new_n686_), .ZN(new_n929_));
  XOR2_X1   g728(.A(KEYINPUT63), .B(G211gat), .Z(new_n930_));
  NOR3_X1   g729(.A1(new_n922_), .A2(new_n595_), .A3(new_n930_), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n929_), .A2(new_n931_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(KEYINPUT126), .ZN(G1354gat));
  AND3_X1   g732(.A1(new_n925_), .A2(G218gat), .A3(new_n573_), .ZN(new_n934_));
  NOR3_X1   g733(.A1(new_n922_), .A2(KEYINPUT127), .A3(new_n648_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n935_), .A2(G218gat), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT127), .B1(new_n922_), .B2(new_n648_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n934_), .B1(new_n936_), .B2(new_n937_), .ZN(G1355gat));
endmodule


