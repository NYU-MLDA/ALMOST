//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n596_, new_n597_, new_n598_, new_n599_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n639_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n645_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n656_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n809_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_;
  XNOR2_X1  g000(.A(KEYINPUT82), .B(G183gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT25), .ZN(new_n203_));
  OAI21_X1  g002(.A(new_n203_), .B1(KEYINPUT25), .B2(G183gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT24), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(G169gat), .B2(G176gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n208_), .B1(G169gat), .B2(G176gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G183gat), .A2(G190gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT23), .ZN(new_n211_));
  OR3_X1    g010(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n209_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n206_), .A2(new_n213_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n211_), .B1(G190gat), .B2(new_n202_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT83), .B(G176gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT22), .B(G169gat), .ZN(new_n217_));
  AOI22_X1  g016(.A1(new_n216_), .A2(new_n217_), .B1(G169gat), .B2(G176gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G227gat), .A2(G233gat), .ZN(new_n221_));
  INV_X1    g020(.A(G15gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(KEYINPUT30), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n220_), .B(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G127gat), .B(G134gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G113gat), .B(G120gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT84), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT85), .B1(new_n226_), .B2(new_n227_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n226_), .A2(new_n227_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT85), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n230_), .A2(new_n231_), .A3(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(new_n225_), .B(new_n235_), .Z(new_n236_));
  XNOR2_X1  g035(.A(G71gat), .B(G99gat), .ZN(new_n237_));
  INV_X1    g036(.A(G43gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT31), .ZN(new_n240_));
  OR2_X1    g039(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n236_), .A2(new_n240_), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G1gat), .B(G29gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(G85gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT0), .B(G57gat), .ZN(new_n246_));
  XOR2_X1   g045(.A(new_n245_), .B(new_n246_), .Z(new_n247_));
  INV_X1    g046(.A(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT4), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G141gat), .A2(G148gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT86), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G141gat), .A2(G148gat), .ZN(new_n252_));
  NAND3_X1  g051(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n253_));
  AND3_X1   g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(G155gat), .B(G162gat), .Z(new_n255_));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT3), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n250_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT2), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n252_), .A2(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n259_), .A2(new_n261_), .A3(new_n262_), .A4(new_n263_), .ZN(new_n264_));
  AOI22_X1  g063(.A1(new_n254_), .A2(new_n257_), .B1(new_n255_), .B2(new_n264_), .ZN(new_n265_));
  OR2_X1    g064(.A1(new_n235_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n228_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n265_), .B1(new_n267_), .B2(new_n232_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n249_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n269_), .B1(new_n249_), .B2(new_n266_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G225gat), .A2(G233gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n266_), .A2(new_n268_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(new_n271_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n248_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n273_), .A2(new_n248_), .A3(new_n275_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(G204gat), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n281_), .A2(G197gat), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(G197gat), .ZN(new_n283_));
  OAI21_X1  g082(.A(KEYINPUT21), .B1(new_n282_), .B2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G211gat), .B(G218gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT88), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n283_), .B1(new_n282_), .B2(new_n286_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n287_), .B1(new_n286_), .B2(new_n282_), .ZN(new_n288_));
  OAI211_X1 g087(.A(new_n284_), .B(new_n285_), .C1(new_n288_), .C2(KEYINPUT21), .ZN(new_n289_));
  INV_X1    g088(.A(new_n285_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n288_), .A2(KEYINPUT21), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n289_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n220_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT20), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G226gat), .A2(G233gat), .ZN(new_n295_));
  XNOR2_X1  g094(.A(new_n295_), .B(KEYINPUT19), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n211_), .B1(G183gat), .B2(G190gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT93), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n218_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT25), .B(G183gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n205_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n213_), .A2(new_n303_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n304_), .A2(KEYINPUT92), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(KEYINPUT92), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n301_), .A2(new_n305_), .A3(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n297_), .B1(new_n292_), .B2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G8gat), .B(G36gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT18), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G64gat), .B(G92gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n296_), .B(KEYINPUT91), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT20), .B1(new_n220_), .B2(new_n292_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n314_), .B1(new_n307_), .B2(new_n292_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n308_), .B(new_n312_), .C1(new_n313_), .C2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT27), .ZN(new_n317_));
  INV_X1    g116(.A(new_n292_), .ZN(new_n318_));
  AND3_X1   g117(.A1(new_n318_), .A2(new_n301_), .A3(new_n304_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n296_), .B1(new_n319_), .B2(new_n294_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT97), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n315_), .A2(new_n313_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n312_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n317_), .B1(new_n325_), .B2(KEYINPUT98), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT98), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n323_), .A2(new_n327_), .A3(new_n324_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n308_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n324_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(KEYINPUT94), .A3(new_n316_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT94), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n330_), .A2(new_n333_), .A3(new_n324_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT27), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  OAI211_X1 g137(.A(G228gat), .B(G233gat), .C1(new_n318_), .C2(KEYINPUT89), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(G106gat), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT29), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n292_), .B1(new_n265_), .B2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G78gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n340_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT90), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n265_), .A2(new_n341_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n346_), .B(new_n347_), .ZN(new_n348_));
  XOR2_X1   g147(.A(G22gat), .B(G50gat), .Z(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n344_), .A2(new_n345_), .A3(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n345_), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n351_), .B1(new_n352_), .B2(new_n344_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  AND4_X1   g153(.A1(new_n280_), .A2(new_n329_), .A3(new_n338_), .A4(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT95), .ZN(new_n356_));
  OR3_X1    g155(.A1(new_n276_), .A2(new_n356_), .A3(KEYINPUT33), .ZN(new_n357_));
  OAI21_X1  g156(.A(KEYINPUT33), .B1(new_n276_), .B2(new_n356_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n266_), .A2(new_n268_), .A3(new_n272_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n248_), .B(new_n359_), .C1(new_n270_), .C2(new_n272_), .ZN(new_n360_));
  NAND4_X1  g159(.A1(new_n357_), .A2(new_n335_), .A3(new_n358_), .A4(new_n360_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n312_), .A2(KEYINPUT32), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n321_), .A2(new_n322_), .A3(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n330_), .A2(KEYINPUT96), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT96), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n330_), .A2(new_n365_), .ZN(new_n366_));
  OAI22_X1  g165(.A1(new_n363_), .A2(new_n364_), .B1(new_n366_), .B2(new_n362_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(new_n279_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n354_), .B1(new_n361_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n243_), .B1(new_n355_), .B2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(new_n243_), .A2(new_n279_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n329_), .A2(new_n338_), .A3(new_n353_), .A4(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT99), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  AOI22_X1  g173(.A1(new_n328_), .A2(new_n326_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n375_), .A2(KEYINPUT99), .A3(new_n353_), .A4(new_n371_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n370_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n379_));
  OR2_X1    g178(.A1(KEYINPUT69), .A2(KEYINPUT13), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G120gat), .B(G148gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT5), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G176gat), .B(G204gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n382_), .B(new_n383_), .Z(new_n384_));
  NAND2_X1  g183(.A1(G99gat), .A2(G106gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT6), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT6), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(G99gat), .A3(G106gat), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  OR2_X1    g188(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n390_));
  INV_X1    g189(.A(G106gat), .ZN(new_n391_));
  NAND2_X1  g190(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n389_), .B1(KEYINPUT64), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT64), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n390_), .A2(new_n395_), .A3(new_n391_), .A4(new_n392_), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT9), .ZN(new_n397_));
  AND2_X1   g196(.A1(G85gat), .A2(G92gat), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G85gat), .A2(G92gat), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n397_), .B1(new_n400_), .B2(KEYINPUT65), .ZN(new_n401_));
  INV_X1    g200(.A(G85gat), .ZN(new_n402_));
  INV_X1    g201(.A(G92gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G85gat), .A2(G92gat), .ZN(new_n405_));
  NAND4_X1  g204(.A1(new_n404_), .A2(KEYINPUT65), .A3(new_n397_), .A4(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n404_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n394_), .B(new_n396_), .C1(new_n401_), .C2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G57gat), .B(G64gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(KEYINPUT11), .ZN(new_n410_));
  XOR2_X1   g209(.A(G71gat), .B(G78gat), .Z(new_n411_));
  OR2_X1    g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n409_), .A2(KEYINPUT11), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n410_), .A2(new_n411_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n412_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT8), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n386_), .A2(new_n388_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT67), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT7), .ZN(new_n420_));
  INV_X1    g219(.A(G99gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n420_), .A2(new_n421_), .A3(new_n391_), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n386_), .A2(new_n388_), .A3(KEYINPUT67), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n419_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n416_), .B1(new_n427_), .B2(new_n400_), .ZN(new_n428_));
  XOR2_X1   g227(.A(KEYINPUT66), .B(KEYINPUT8), .Z(new_n429_));
  INV_X1    g228(.A(new_n400_), .ZN(new_n430_));
  AOI211_X1 g229(.A(new_n429_), .B(new_n430_), .C1(new_n417_), .C2(new_n425_), .ZN(new_n431_));
  OAI211_X1 g230(.A(new_n408_), .B(new_n415_), .C1(new_n428_), .C2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G230gat), .A2(G233gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n407_), .A2(new_n401_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n393_), .A2(KEYINPUT64), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n436_), .A2(new_n417_), .A3(new_n396_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  AND3_X1   g237(.A1(new_n386_), .A2(new_n388_), .A3(KEYINPUT67), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT67), .B1(new_n386_), .B2(new_n388_), .ZN(new_n440_));
  NOR3_X1   g239(.A1(new_n439_), .A2(new_n440_), .A3(new_n424_), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT8), .B1(new_n441_), .B2(new_n430_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n430_), .A2(new_n429_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n443_), .B1(new_n389_), .B2(new_n424_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n438_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT12), .B1(new_n445_), .B2(new_n415_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n408_), .B1(new_n428_), .B2(new_n431_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT12), .ZN(new_n448_));
  INV_X1    g247(.A(new_n415_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n434_), .B1(new_n446_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n447_), .A2(new_n449_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n433_), .B1(new_n452_), .B2(new_n432_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n384_), .B1(new_n451_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n433_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n455_), .B1(new_n445_), .B2(new_n415_), .ZN(new_n456_));
  AND3_X1   g255(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n448_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n456_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n452_), .A2(new_n432_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n460_), .A2(new_n455_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n384_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n459_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  AND3_X1   g262(.A1(new_n454_), .A2(KEYINPUT68), .A3(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(KEYINPUT68), .B1(new_n454_), .B2(new_n463_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n379_), .B(new_n380_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT68), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n451_), .A2(new_n453_), .A3(new_n384_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n462_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n467_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n454_), .A2(KEYINPUT68), .A3(new_n463_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n470_), .A2(KEYINPUT69), .A3(KEYINPUT13), .A4(new_n471_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n466_), .A2(KEYINPUT70), .A3(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(KEYINPUT70), .B1(new_n466_), .B2(new_n472_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G29gat), .B(G36gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G43gat), .B(G50gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT71), .B(KEYINPUT15), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n479_), .B(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(new_n447_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT74), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n477_), .B(new_n478_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n408_), .B(new_n484_), .C1(new_n428_), .C2(new_n431_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G232gat), .A2(G233gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT34), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n487_), .B(KEYINPUT35), .Z(new_n488_));
  NAND4_X1  g287(.A1(new_n482_), .A2(new_n483_), .A3(new_n485_), .A4(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n482_), .A2(new_n485_), .A3(new_n488_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT74), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n487_), .A2(KEYINPUT35), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n492_), .B1(new_n482_), .B2(new_n485_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n489_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G190gat), .B(G218gat), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT72), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G134gat), .B(G162gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n497_), .B(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(KEYINPUT73), .B(KEYINPUT36), .Z(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n494_), .A2(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n499_), .B(KEYINPUT36), .ZN(new_n504_));
  OAI211_X1 g303(.A(new_n489_), .B(new_n504_), .C1(new_n491_), .C2(new_n493_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(KEYINPUT76), .B(KEYINPUT37), .Z(new_n508_));
  XOR2_X1   g307(.A(new_n504_), .B(KEYINPUT75), .Z(new_n509_));
  OAI21_X1  g308(.A(new_n503_), .B1(new_n494_), .B2(new_n509_), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n507_), .A2(new_n508_), .B1(new_n510_), .B2(KEYINPUT37), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G1gat), .B(G8gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT77), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G15gat), .B(G22gat), .ZN(new_n514_));
  INV_X1    g313(.A(G1gat), .ZN(new_n515_));
  INV_X1    g314(.A(G8gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT14), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n514_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n513_), .A2(new_n518_), .ZN(new_n519_));
  OR2_X1    g318(.A1(new_n512_), .A2(KEYINPUT77), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n512_), .A2(KEYINPUT77), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n520_), .A2(new_n517_), .A3(new_n514_), .A4(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n519_), .A2(new_n522_), .ZN(new_n523_));
  OR2_X1    g322(.A1(new_n414_), .A2(new_n413_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G231gat), .A2(G233gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n412_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n524_), .B2(new_n412_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n523_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n528_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n519_), .A2(new_n522_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(new_n526_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(new_n532_), .A3(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(G127gat), .B(G155gat), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT16), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G183gat), .B(G211gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT78), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n529_), .A2(new_n532_), .A3(new_n540_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n538_), .A2(KEYINPUT17), .ZN(new_n542_));
  AND3_X1   g341(.A1(new_n539_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n541_), .B1(new_n539_), .B2(new_n542_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n511_), .A2(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n476_), .A2(new_n547_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n548_), .A2(KEYINPUT79), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(KEYINPUT79), .ZN(new_n550_));
  XOR2_X1   g349(.A(G113gat), .B(G141gat), .Z(new_n551_));
  XOR2_X1   g350(.A(G169gat), .B(G197gat), .Z(new_n552_));
  XOR2_X1   g351(.A(new_n551_), .B(new_n552_), .Z(new_n553_));
  XOR2_X1   g352(.A(new_n553_), .B(KEYINPUT80), .Z(new_n554_));
  XNOR2_X1  g353(.A(new_n484_), .B(new_n480_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n555_), .A2(new_n531_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n523_), .A2(new_n479_), .ZN(new_n559_));
  NOR3_X1   g358(.A1(new_n556_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n559_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n523_), .A2(new_n479_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n557_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n554_), .B1(new_n560_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT81), .ZN(new_n565_));
  INV_X1    g364(.A(new_n553_), .ZN(new_n566_));
  OR3_X1    g365(.A1(new_n560_), .A2(new_n563_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT81), .ZN(new_n568_));
  OAI211_X1 g367(.A(new_n568_), .B(new_n554_), .C1(new_n560_), .C2(new_n563_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n565_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n570_));
  NAND4_X1  g369(.A1(new_n378_), .A2(new_n549_), .A3(new_n550_), .A4(new_n570_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n571_), .A2(G1gat), .A3(new_n280_), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n573_));
  AND2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n572_), .A2(new_n573_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n476_), .A2(new_n570_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n378_), .A2(new_n577_), .ZN(new_n578_));
  NOR3_X1   g377(.A1(new_n578_), .A2(new_n546_), .A3(new_n507_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n515_), .B1(new_n579_), .B2(new_n279_), .ZN(new_n580_));
  OR3_X1    g379(.A1(new_n574_), .A2(new_n575_), .A3(new_n580_), .ZN(G1324gat));
  INV_X1    g380(.A(KEYINPUT39), .ZN(new_n582_));
  INV_X1    g381(.A(new_n375_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n579_), .A2(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n582_), .B1(new_n584_), .B2(G8gat), .ZN(new_n585_));
  AOI211_X1 g384(.A(KEYINPUT39), .B(new_n516_), .C1(new_n579_), .C2(new_n583_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n516_), .ZN(new_n587_));
  OAI22_X1  g386(.A1(new_n585_), .A2(new_n586_), .B1(new_n571_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT40), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(G1325gat));
  INV_X1    g389(.A(new_n243_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n222_), .B1(new_n579_), .B2(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT41), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n222_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n593_), .B1(new_n571_), .B2(new_n594_), .ZN(G1326gat));
  INV_X1    g394(.A(G22gat), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n596_), .B1(new_n579_), .B2(new_n354_), .ZN(new_n597_));
  XOR2_X1   g396(.A(new_n597_), .B(KEYINPUT42), .Z(new_n598_));
  NAND2_X1  g397(.A1(new_n354_), .A2(new_n596_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n598_), .B1(new_n571_), .B2(new_n599_), .ZN(G1327gat));
  NAND3_X1  g399(.A1(new_n375_), .A2(new_n280_), .A3(new_n354_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n361_), .A2(new_n368_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(new_n353_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n601_), .A2(new_n603_), .ZN(new_n604_));
  AOI22_X1  g403(.A1(new_n604_), .A2(new_n243_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(new_n576_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n545_), .A2(new_n506_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  OR3_X1    g407(.A1(new_n608_), .A2(G29gat), .A3(new_n280_), .ZN(new_n609_));
  OR2_X1    g408(.A1(KEYINPUT101), .A2(KEYINPUT43), .ZN(new_n610_));
  NAND2_X1  g409(.A1(KEYINPUT101), .A2(KEYINPUT43), .ZN(new_n611_));
  INV_X1    g410(.A(new_n511_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n610_), .B(new_n611_), .C1(new_n605_), .C2(new_n612_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n378_), .A2(KEYINPUT101), .A3(KEYINPUT43), .A4(new_n511_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n577_), .A2(new_n546_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n613_), .A2(new_n614_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT44), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n613_), .A2(KEYINPUT44), .A3(new_n614_), .A4(new_n616_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n619_), .A2(new_n279_), .A3(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT102), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G29gat), .B1(new_n621_), .B2(new_n622_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n609_), .B1(new_n623_), .B2(new_n624_), .ZN(G1328gat));
  INV_X1    g424(.A(KEYINPUT103), .ZN(new_n626_));
  XNOR2_X1  g425(.A(KEYINPUT104), .B(KEYINPUT46), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n619_), .A2(new_n583_), .A3(new_n620_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n628_), .A2(G36gat), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n375_), .A2(G36gat), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n606_), .A2(new_n607_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT45), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n626_), .B(new_n627_), .C1(new_n629_), .C2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n627_), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n633_), .B1(new_n628_), .B2(G36gat), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n635_), .B1(new_n636_), .B2(KEYINPUT103), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(G1329gat));
  NAND4_X1  g437(.A1(new_n619_), .A2(G43gat), .A3(new_n591_), .A4(new_n620_), .ZN(new_n639_));
  OAI21_X1  g438(.A(new_n238_), .B1(new_n608_), .B2(new_n243_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g441(.A1(new_n619_), .A2(G50gat), .A3(new_n354_), .A4(new_n620_), .ZN(new_n643_));
  INV_X1    g442(.A(G50gat), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n644_), .B1(new_n608_), .B2(new_n353_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n643_), .A2(new_n645_), .ZN(G1331gat));
  AOI211_X1 g445(.A(new_n476_), .B(new_n570_), .C1(new_n370_), .C2(new_n377_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n647_), .A2(new_n547_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n649_), .A2(G57gat), .A3(new_n280_), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n647_), .A2(new_n545_), .A3(new_n506_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(new_n279_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n650_), .B1(G57gat), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT105), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(G1332gat));
  OR3_X1    g454(.A1(new_n649_), .A2(G64gat), .A3(new_n375_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n651_), .A2(new_n583_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(G64gat), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n658_), .A2(KEYINPUT48), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(KEYINPUT48), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n656_), .B1(new_n659_), .B2(new_n660_), .ZN(G1333gat));
  OR3_X1    g460(.A1(new_n649_), .A2(G71gat), .A3(new_n243_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n651_), .A2(new_n591_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(G71gat), .ZN(new_n664_));
  AND2_X1   g463(.A1(new_n664_), .A2(KEYINPUT49), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(KEYINPUT49), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n662_), .B1(new_n665_), .B2(new_n666_), .ZN(G1334gat));
  OR3_X1    g466(.A1(new_n649_), .A2(G78gat), .A3(new_n353_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n651_), .A2(new_n354_), .ZN(new_n669_));
  XOR2_X1   g468(.A(KEYINPUT106), .B(KEYINPUT50), .Z(new_n670_));
  AND3_X1   g469(.A1(new_n669_), .A2(G78gat), .A3(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n670_), .B1(new_n669_), .B2(G78gat), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n668_), .B1(new_n671_), .B2(new_n672_), .ZN(G1335gat));
  AND2_X1   g472(.A1(new_n647_), .A2(new_n607_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n674_), .A2(new_n402_), .A3(new_n279_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n613_), .A2(new_n614_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n476_), .A2(new_n545_), .A3(new_n570_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n678_), .A2(new_n279_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n675_), .B1(new_n679_), .B2(new_n402_), .ZN(G1336gat));
  NAND3_X1  g479(.A1(new_n674_), .A2(new_n403_), .A3(new_n583_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n678_), .A2(new_n583_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n682_), .B2(new_n403_), .ZN(G1337gat));
  AND3_X1   g482(.A1(new_n591_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n674_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT107), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n685_), .B(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n676_), .A2(new_n591_), .A3(new_n677_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(G99gat), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(KEYINPUT51), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT51), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n687_), .A2(new_n692_), .A3(new_n689_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1338gat));
  NAND3_X1  g493(.A1(new_n674_), .A2(new_n391_), .A3(new_n354_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n613_), .A2(new_n354_), .A3(new_n614_), .A4(new_n677_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT52), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n696_), .A2(new_n697_), .A3(G106gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n696_), .B2(G106gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n695_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n700_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g500(.A(KEYINPUT117), .ZN(new_n702_));
  NOR3_X1   g501(.A1(new_n570_), .A2(new_n544_), .A3(new_n543_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n466_), .A2(new_n472_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n466_), .A2(new_n703_), .A3(new_n472_), .A4(KEYINPUT108), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n706_), .A2(new_n612_), .A3(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT109), .B(KEYINPUT54), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT110), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n708_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT111), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n709_), .A2(new_n710_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n708_), .A2(KEYINPUT111), .A3(new_n711_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n714_), .A2(new_n715_), .A3(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n715_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n711_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n511_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n720_));
  AOI211_X1 g519(.A(new_n713_), .B(new_n719_), .C1(new_n720_), .C2(new_n707_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT111), .B1(new_n708_), .B2(new_n711_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n718_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n717_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT112), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT55), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n725_), .B1(new_n459_), .B2(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n451_), .A2(KEYINPUT112), .A3(KEYINPUT55), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n459_), .A2(new_n726_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n432_), .B1(new_n457_), .B2(new_n458_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(new_n455_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n727_), .A2(new_n728_), .A3(new_n729_), .A4(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n732_), .A2(KEYINPUT56), .A3(new_n384_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT115), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT56), .B1(new_n732_), .B2(new_n384_), .ZN(new_n736_));
  INV_X1    g535(.A(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n732_), .A2(KEYINPUT115), .A3(KEYINPUT56), .A4(new_n384_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n735_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n556_), .A2(new_n557_), .A3(new_n559_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n558_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n741_));
  OR3_X1    g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n553_), .ZN(new_n742_));
  AND2_X1   g541(.A1(new_n567_), .A2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(new_n463_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(KEYINPUT58), .B1(new_n739_), .B2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT116), .B1(new_n746_), .B2(new_n612_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT116), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n736_), .B1(new_n734_), .B2(new_n733_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n744_), .B1(new_n749_), .B2(new_n738_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n748_), .B(new_n511_), .C1(new_n750_), .C2(KEYINPUT58), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(KEYINPUT58), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n747_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT114), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT57), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n754_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n757_));
  AND2_X1   g556(.A1(new_n570_), .A2(new_n463_), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n732_), .A2(KEYINPUT56), .A3(new_n384_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n759_), .B2(new_n736_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n743_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n757_), .B1(new_n762_), .B2(new_n507_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n507_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n755_), .B1(new_n764_), .B2(new_n754_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n763_), .B1(new_n765_), .B2(KEYINPUT57), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n545_), .B1(new_n753_), .B2(new_n766_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n702_), .B1(new_n724_), .B2(new_n767_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n753_), .A2(new_n766_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n546_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n770_), .A2(KEYINPUT117), .A3(new_n717_), .A4(new_n723_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n768_), .A2(new_n771_), .ZN(new_n772_));
  NOR4_X1   g571(.A1(new_n583_), .A2(new_n280_), .A3(new_n354_), .A4(new_n243_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(G113gat), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n774_), .A2(new_n775_), .A3(new_n570_), .ZN(new_n776_));
  AND2_X1   g575(.A1(new_n717_), .A2(new_n723_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(new_n770_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n773_), .B1(KEYINPUT118), .B2(KEYINPUT59), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n778_), .B(new_n779_), .C1(KEYINPUT118), .C2(new_n773_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT59), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n570_), .B(new_n780_), .C1(new_n774_), .C2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n776_), .B1(new_n783_), .B2(new_n775_), .ZN(G1340gat));
  INV_X1    g583(.A(KEYINPUT60), .ZN(new_n785_));
  AOI21_X1  g584(.A(G120gat), .B1(new_n475_), .B2(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n785_), .B2(G120gat), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n774_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n780_), .B1(new_n774_), .B2(new_n781_), .ZN(new_n791_));
  OAI21_X1  g590(.A(G120gat), .B1(new_n791_), .B2(new_n476_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n790_), .A2(new_n792_), .ZN(G1341gat));
  INV_X1    g592(.A(G127gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n774_), .A2(new_n794_), .A3(new_n545_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n545_), .B(new_n780_), .C1(new_n774_), .C2(new_n781_), .ZN(new_n796_));
  INV_X1    g595(.A(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n797_), .B2(new_n794_), .ZN(G1342gat));
  INV_X1    g597(.A(G134gat), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n774_), .A2(new_n799_), .A3(new_n507_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n511_), .B(new_n780_), .C1(new_n774_), .C2(new_n781_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n802_), .B2(new_n799_), .ZN(G1343gat));
  NOR4_X1   g602(.A1(new_n583_), .A2(new_n280_), .A3(new_n353_), .A4(new_n591_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n805_), .B1(new_n768_), .B2(new_n771_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n570_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n475_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g609(.A1(new_n806_), .A2(new_n545_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(KEYINPUT61), .B(G155gat), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n811_), .B(new_n812_), .ZN(G1346gat));
  NAND3_X1  g612(.A1(new_n806_), .A2(G162gat), .A3(new_n511_), .ZN(new_n814_));
  AOI211_X1 g613(.A(KEYINPUT120), .B(G162gat), .C1(new_n806_), .C2(new_n507_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n816_));
  AOI21_X1  g615(.A(KEYINPUT117), .B1(new_n777_), .B2(new_n770_), .ZN(new_n817_));
  NOR3_X1   g616(.A1(new_n724_), .A2(new_n767_), .A3(new_n702_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n507_), .B(new_n804_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(G162gat), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n816_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n814_), .B1(new_n815_), .B2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT121), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n822_), .A2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(KEYINPUT121), .B(new_n814_), .C1(new_n815_), .C2(new_n821_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(G1347gat));
  NOR3_X1   g625(.A1(new_n375_), .A2(new_n279_), .A3(new_n243_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n827_), .A2(new_n353_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n570_), .A2(new_n217_), .ZN(new_n829_));
  XOR2_X1   g628(.A(new_n829_), .B(KEYINPUT122), .Z(new_n830_));
  NAND3_X1  g629(.A1(new_n778_), .A2(new_n828_), .A3(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n778_), .A2(new_n570_), .A3(new_n828_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT62), .ZN(new_n833_));
  AND3_X1   g632(.A1(new_n832_), .A2(new_n833_), .A3(G169gat), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n833_), .B1(new_n832_), .B2(G169gat), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(G1348gat));
  NAND2_X1  g635(.A1(new_n772_), .A2(new_n353_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT123), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n772_), .A2(KEYINPUT123), .A3(new_n353_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n839_), .A2(new_n827_), .A3(new_n840_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n475_), .A2(G176gat), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n778_), .A2(new_n475_), .A3(new_n828_), .ZN(new_n843_));
  AOI22_X1  g642(.A1(new_n841_), .A2(new_n842_), .B1(new_n216_), .B2(new_n843_), .ZN(G1349gat));
  NOR2_X1   g643(.A1(new_n546_), .A2(new_n302_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n778_), .A2(new_n828_), .A3(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n841_), .A2(new_n545_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n202_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n847_), .B1(new_n848_), .B2(new_n849_), .ZN(G1350gat));
  NAND4_X1  g649(.A1(new_n778_), .A2(new_n507_), .A3(new_n205_), .A4(new_n828_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n778_), .A2(new_n511_), .A3(new_n828_), .ZN(new_n852_));
  AND3_X1   g651(.A1(new_n852_), .A2(KEYINPUT124), .A3(G190gat), .ZN(new_n853_));
  AOI21_X1  g652(.A(KEYINPUT124), .B1(new_n852_), .B2(G190gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n851_), .B1(new_n853_), .B2(new_n854_), .ZN(G1351gat));
  NAND4_X1  g654(.A1(new_n583_), .A2(new_n280_), .A3(new_n354_), .A4(new_n243_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n856_), .B1(new_n768_), .B2(new_n771_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n570_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g658(.A1(new_n857_), .A2(new_n475_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n281_), .A2(KEYINPUT125), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n281_), .A2(KEYINPUT125), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n860_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n863_), .B1(new_n860_), .B2(new_n862_), .ZN(G1353gat));
  AND2_X1   g663(.A1(new_n857_), .A2(new_n545_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n865_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT63), .B(G211gat), .Z(new_n867_));
  AOI21_X1  g666(.A(new_n866_), .B1(new_n865_), .B2(new_n867_), .ZN(G1354gat));
  NAND2_X1  g667(.A1(new_n857_), .A2(new_n507_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT126), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT127), .B(G218gat), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n612_), .A2(new_n871_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n870_), .A2(new_n871_), .B1(new_n857_), .B2(new_n872_), .ZN(G1355gat));
endmodule


