//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 1 0 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n769_, new_n770_,
    new_n771_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n953_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_;
  NOR2_X1   g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n203_));
  XOR2_X1   g002(.A(new_n202_), .B(new_n203_), .Z(new_n204_));
  NAND2_X1  g003(.A1(G99gat), .A2(G106gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n205_), .B(KEYINPUT6), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G85gat), .B(G92gat), .Z(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT8), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n207_), .A2(KEYINPUT8), .A3(new_n208_), .ZN(new_n212_));
  XOR2_X1   g011(.A(KEYINPUT10), .B(G99gat), .Z(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n208_), .A2(KEYINPUT9), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT9), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(G85gat), .A3(G92gat), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n215_), .A2(new_n216_), .A3(new_n206_), .A4(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n211_), .A2(new_n212_), .A3(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(G29gat), .B(G36gat), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n221_), .A2(KEYINPUT67), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(KEYINPUT67), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G43gat), .B(G50gat), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n224_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n222_), .A2(new_n223_), .A3(new_n225_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT15), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(KEYINPUT15), .B1(new_n227_), .B2(new_n228_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n220_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(KEYINPUT8), .B1(new_n207_), .B2(new_n208_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n219_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n236_), .A2(new_n228_), .A3(new_n227_), .A4(new_n212_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n233_), .A2(KEYINPUT71), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT35), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n233_), .A2(new_n241_), .A3(KEYINPUT71), .A4(new_n237_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G232gat), .A2(G233gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n243_), .B(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n240_), .A2(new_n242_), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT71), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n229_), .B(new_n230_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n248_), .B2(new_n220_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n245_), .ZN(new_n250_));
  NAND4_X1  g049(.A1(new_n249_), .A2(new_n241_), .A3(new_n237_), .A4(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G190gat), .B(G218gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G134gat), .B(G162gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n252_), .B(new_n253_), .ZN(new_n254_));
  XOR2_X1   g053(.A(KEYINPUT69), .B(KEYINPUT36), .Z(new_n255_));
  NOR2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(new_n256_), .B(KEYINPUT70), .Z(new_n257_));
  NAND3_X1  g056(.A1(new_n246_), .A2(new_n251_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT73), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT35), .B1(new_n249_), .B2(new_n237_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n242_), .A2(new_n245_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n251_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT72), .B(KEYINPUT36), .ZN(new_n263_));
  XOR2_X1   g062(.A(new_n254_), .B(new_n263_), .Z(new_n264_));
  AOI22_X1  g063(.A1(new_n258_), .A2(new_n259_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n262_), .A2(new_n259_), .A3(new_n264_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT37), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT37), .ZN(new_n268_));
  AND3_X1   g067(.A1(new_n262_), .A2(KEYINPUT74), .A3(new_n264_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT74), .B1(new_n262_), .B2(new_n264_), .ZN(new_n270_));
  OAI211_X1 g069(.A(new_n268_), .B(new_n258_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G57gat), .B(G64gat), .ZN(new_n274_));
  OR2_X1    g073(.A1(new_n274_), .A2(KEYINPUT11), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(KEYINPUT11), .ZN(new_n276_));
  XOR2_X1   g075(.A(G71gat), .B(G78gat), .Z(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(new_n276_), .A3(new_n277_), .ZN(new_n278_));
  OR2_X1    g077(.A1(new_n276_), .A2(new_n277_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G231gat), .A2(G233gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G1gat), .B(G8gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT75), .ZN(new_n284_));
  INV_X1    g083(.A(G15gat), .ZN(new_n285_));
  INV_X1    g084(.A(G22gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G15gat), .A2(G22gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(G1gat), .A2(G8gat), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n287_), .A2(new_n288_), .B1(KEYINPUT14), .B2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n284_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n282_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n294_), .A2(KEYINPUT77), .ZN(new_n295_));
  XOR2_X1   g094(.A(G127gat), .B(G155gat), .Z(new_n296_));
  XNOR2_X1  g095(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n296_), .B(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G183gat), .B(G211gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT17), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT78), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n294_), .A2(KEYINPUT77), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n295_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n300_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n294_), .A2(KEYINPUT17), .A3(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n273_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n280_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n220_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n220_), .A2(new_n309_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(KEYINPUT65), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n310_), .B1(new_n312_), .B2(KEYINPUT12), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G230gat), .A2(G233gat), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT12), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n311_), .A2(KEYINPUT65), .A3(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n313_), .A2(KEYINPUT66), .A3(new_n314_), .A4(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n280_), .B1(new_n236_), .B2(new_n212_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT65), .ZN(new_n319_));
  OAI21_X1  g118(.A(KEYINPUT12), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n310_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n320_), .A2(new_n316_), .A3(new_n314_), .A4(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT66), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n314_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n325_), .B1(new_n310_), .B2(new_n318_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n317_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G120gat), .B(G148gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT5), .ZN(new_n329_));
  XNOR2_X1  g128(.A(G176gat), .B(G204gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  XNOR2_X1  g130(.A(new_n327_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(KEYINPUT13), .ZN(new_n333_));
  AND2_X1   g132(.A1(new_n308_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G197gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(G204gat), .ZN(new_n336_));
  INV_X1    g135(.A(G204gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(G197gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT21), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n336_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n340_), .A2(KEYINPUT95), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT95), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n336_), .A2(new_n338_), .A3(new_n342_), .A4(new_n339_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G211gat), .B(G218gat), .Z(new_n345_));
  INV_X1    g144(.A(KEYINPUT94), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n346_), .B1(new_n337_), .B2(G197gat), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n335_), .A2(KEYINPUT94), .A3(G204gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n347_), .A2(new_n338_), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n345_), .B1(new_n349_), .B2(KEYINPUT21), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n339_), .B1(new_n336_), .B2(new_n338_), .ZN(new_n351_));
  AOI22_X1  g150(.A1(new_n344_), .A2(new_n350_), .B1(new_n345_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(G155gat), .ZN(new_n354_));
  INV_X1    g153(.A(G162gat), .ZN(new_n355_));
  OAI21_X1  g154(.A(KEYINPUT1), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT88), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n357_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT88), .B1(G155gat), .B2(G162gat), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT1), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n360_), .A2(G155gat), .A3(G162gat), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n356_), .A2(new_n358_), .A3(new_n359_), .A4(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n363_), .A2(KEYINPUT87), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT87), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(G141gat), .A3(G148gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n364_), .A2(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(G141gat), .A2(G148gat), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n362_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n372_), .B1(new_n367_), .B2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT90), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT3), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(new_n368_), .B2(KEYINPUT89), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT89), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n378_), .A2(G141gat), .A3(G148gat), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n375_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT91), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n368_), .A2(KEYINPUT89), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n378_), .B1(G141gat), .B2(G148gat), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n383_), .A2(KEYINPUT90), .A3(new_n384_), .A4(new_n376_), .ZN(new_n385_));
  NAND4_X1  g184(.A1(new_n374_), .A2(new_n380_), .A3(new_n382_), .A4(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n358_), .B(new_n359_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n370_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT29), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n353_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT93), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n344_), .A2(new_n350_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n351_), .A2(new_n345_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n392_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(G228gat), .ZN(new_n396_));
  INV_X1    g195(.A(G233gat), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(G78gat), .B1(new_n395_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(G78gat), .ZN(new_n400_));
  OAI221_X1 g199(.A(new_n400_), .B1(new_n396_), .B2(new_n397_), .C1(new_n352_), .C2(new_n392_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n399_), .A2(new_n401_), .A3(G106gat), .ZN(new_n402_));
  AOI21_X1  g201(.A(G106gat), .B1(new_n399_), .B2(new_n401_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n391_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n399_), .A2(new_n401_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n405_), .A2(new_n214_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n391_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n399_), .A2(new_n401_), .A3(G106gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT92), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n404_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n389_), .A2(new_n390_), .ZN(new_n412_));
  XOR2_X1   g211(.A(new_n412_), .B(KEYINPUT28), .Z(new_n413_));
  NAND2_X1  g212(.A1(new_n411_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(new_n413_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n404_), .A2(new_n409_), .A3(new_n415_), .A4(new_n410_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G22gat), .B(G50gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n414_), .A2(new_n418_), .A3(new_n416_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G57gat), .B(G85gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT102), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(G1gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT101), .B(KEYINPUT0), .Z(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(G29gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n425_), .B(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n386_), .A2(new_n388_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT98), .ZN(new_n430_));
  INV_X1    g229(.A(new_n370_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(G134gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(G127gat), .ZN(new_n434_));
  INV_X1    g233(.A(G127gat), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(G134gat), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n434_), .A2(new_n436_), .A3(KEYINPUT86), .ZN(new_n437_));
  INV_X1    g236(.A(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G113gat), .B(G120gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT86), .B1(new_n434_), .B2(new_n436_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n438_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n434_), .A2(new_n436_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT86), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n439_), .B1(new_n445_), .B2(new_n437_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n442_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n432_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n389_), .A2(new_n430_), .A3(new_n447_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G225gat), .A2(G233gat), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n428_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT99), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n440_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n445_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n456_));
  AOI21_X1  g255(.A(KEYINPUT4), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n380_), .A2(new_n385_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT91), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n381_), .B(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(KEYINPUT2), .B1(new_n364_), .B2(new_n366_), .ZN(new_n461_));
  NOR3_X1   g260(.A1(new_n460_), .A2(new_n461_), .A3(new_n372_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n387_), .B1(new_n458_), .B2(new_n462_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n454_), .B(new_n457_), .C1(new_n463_), .C2(new_n370_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT4), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n465_), .B1(new_n442_), .B2(new_n446_), .ZN(new_n466_));
  OAI21_X1  g265(.A(KEYINPUT99), .B1(new_n389_), .B2(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n452_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n449_), .A2(KEYINPUT4), .A3(new_n450_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n468_), .A2(new_n469_), .A3(KEYINPUT100), .ZN(new_n470_));
  AOI21_X1  g269(.A(KEYINPUT100), .B1(new_n468_), .B2(new_n469_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n453_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT103), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  OAI211_X1 g273(.A(KEYINPUT103), .B(new_n453_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n451_), .A2(new_n452_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n476_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n477_));
  AOI22_X1  g276(.A1(new_n474_), .A2(new_n475_), .B1(new_n477_), .B2(new_n428_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G227gat), .A2(G233gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(new_n285_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT30), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(KEYINPUT31), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(G169gat), .ZN(new_n485_));
  AND2_X1   g284(.A1(G183gat), .A2(G190gat), .ZN(new_n486_));
  OR2_X1    g285(.A1(new_n486_), .A2(KEYINPUT23), .ZN(new_n487_));
  AND2_X1   g286(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n488_));
  NOR2_X1   g287(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n486_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  NOR2_X1   g290(.A1(G183gat), .A2(G190gat), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n485_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  OR3_X1    g292(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT84), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G183gat), .A2(G190gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n496_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(KEYINPUT23), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n495_), .B1(new_n497_), .B2(new_n499_), .ZN(new_n500_));
  NOR2_X1   g299(.A1(new_n498_), .A2(KEYINPUT84), .ZN(new_n501_));
  OAI211_X1 g300(.A(KEYINPUT85), .B(new_n494_), .C1(new_n500_), .C2(new_n501_), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(G169gat), .ZN(new_n505_));
  INV_X1    g304(.A(G176gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n504_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT26), .B(G190gat), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT25), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT82), .B1(new_n510_), .B2(G183gat), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT25), .B(G183gat), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n513_), .A2(KEYINPUT82), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n508_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n502_), .A2(new_n515_), .ZN(new_n516_));
  OR2_X1    g315(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n517_));
  NAND2_X1  g316(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n486_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT84), .B1(new_n519_), .B2(new_n498_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n501_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(KEYINPUT85), .B1(new_n522_), .B2(new_n494_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n493_), .B1(new_n516_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G71gat), .B(G99gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(G43gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n524_), .B(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(new_n448_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n527_), .A2(new_n448_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n483_), .B1(new_n529_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n530_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(new_n482_), .A3(new_n528_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n478_), .A2(new_n534_), .ZN(new_n535_));
  OAI22_X1  g334(.A1(new_n500_), .A2(new_n501_), .B1(G183gat), .B2(G190gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n509_), .A2(new_n513_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n537_), .A2(new_n507_), .A3(new_n494_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n491_), .ZN(new_n539_));
  AOI22_X1  g338(.A1(new_n536_), .A2(new_n485_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT96), .B1(new_n540_), .B2(new_n352_), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n539_), .A2(new_n537_), .A3(new_n494_), .A4(new_n507_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n492_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n485_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n542_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT96), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(new_n353_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n541_), .A2(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(G226gat), .A2(G233gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n549_), .B(KEYINPUT19), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n352_), .B(new_n493_), .C1(new_n516_), .C2(new_n523_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n548_), .A2(KEYINPUT20), .A3(new_n551_), .A4(new_n552_), .ZN(new_n553_));
  OAI21_X1  g352(.A(new_n494_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT85), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n556_), .A2(new_n502_), .A3(new_n515_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n352_), .B1(new_n557_), .B2(new_n493_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT20), .B1(new_n545_), .B2(new_n353_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n550_), .B1(new_n558_), .B2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n553_), .A2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G8gat), .B(G36gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G64gat), .B(G92gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n561_), .A2(new_n567_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n540_), .A2(KEYINPUT96), .A3(new_n352_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n546_), .B1(new_n545_), .B2(new_n353_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n552_), .A2(KEYINPUT20), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n550_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n558_), .A2(new_n559_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(new_n551_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n575_), .A3(new_n566_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n568_), .A2(new_n576_), .A3(KEYINPUT27), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n552_), .A2(KEYINPUT20), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n551_), .B1(new_n578_), .B2(new_n548_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n558_), .A2(new_n550_), .A3(new_n559_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n579_), .A2(new_n567_), .A3(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n566_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n577_), .B1(new_n583_), .B2(KEYINPUT27), .ZN(new_n584_));
  NOR3_X1   g383(.A1(new_n422_), .A2(new_n535_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT27), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n567_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n588_), .A2(new_n576_), .ZN(new_n589_));
  AOI22_X1  g388(.A1(new_n587_), .A2(new_n568_), .B1(new_n589_), .B2(new_n586_), .ZN(new_n590_));
  AND3_X1   g389(.A1(new_n414_), .A2(new_n418_), .A3(new_n416_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n418_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n590_), .B(new_n478_), .C1(new_n591_), .C2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n477_), .A2(new_n428_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n468_), .A2(new_n469_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT100), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n468_), .A2(new_n469_), .A3(KEYINPUT100), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(KEYINPUT103), .B1(new_n599_), .B2(new_n453_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n475_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n594_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n561_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n566_), .A2(KEYINPUT32), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n579_), .A2(new_n580_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n605_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT33), .B1(new_n599_), .B2(new_n453_), .ZN(new_n608_));
  OAI211_X1 g407(.A(KEYINPUT33), .B(new_n453_), .C1(new_n470_), .C2(new_n471_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n452_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n451_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n612_), .B1(new_n464_), .B2(new_n467_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(new_n469_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n613_), .A2(new_n615_), .A3(new_n428_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n588_), .A2(new_n576_), .A3(new_n616_), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n602_), .A2(new_n607_), .B1(new_n611_), .B2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n593_), .B1(new_n618_), .B2(new_n422_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n534_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n585_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT79), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n229_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n227_), .A2(KEYINPUT79), .A3(new_n228_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n623_), .A2(new_n291_), .A3(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(KEYINPUT80), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT80), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n623_), .A2(new_n627_), .A3(new_n291_), .A4(new_n624_), .ZN(new_n628_));
  AOI22_X1  g427(.A1(new_n626_), .A2(new_n628_), .B1(new_n292_), .B2(new_n248_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(G229gat), .A2(G233gat), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n626_), .A2(new_n628_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n623_), .A2(new_n624_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(new_n292_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n632_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n631_), .B1(new_n636_), .B2(new_n630_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G113gat), .B(G141gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(G169gat), .B(G197gat), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n638_), .B(new_n639_), .Z(new_n640_));
  INV_X1    g439(.A(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n637_), .A2(new_n641_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n631_), .B(new_n640_), .C1(new_n636_), .C2(new_n630_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(KEYINPUT81), .A3(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT81), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n637_), .A2(new_n645_), .A3(new_n641_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n621_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n334_), .A2(new_n648_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n649_), .A2(G1gat), .A3(new_n478_), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT38), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(KEYINPUT38), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n258_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT104), .B(new_n258_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n621_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n647_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n307_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n658_), .A2(new_n659_), .A3(new_n333_), .A4(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G1gat), .B1(new_n661_), .B2(new_n478_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n651_), .A2(new_n652_), .A3(new_n662_), .ZN(G1324gat));
  OAI21_X1  g462(.A(G8gat), .B1(new_n661_), .B2(new_n590_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT39), .ZN(new_n665_));
  OR2_X1    g464(.A1(new_n590_), .A2(G8gat), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n665_), .B1(new_n649_), .B2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT105), .B(KEYINPUT40), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(G1325gat));
  OAI21_X1  g468(.A(G15gat), .B1(new_n661_), .B2(new_n620_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT41), .Z(new_n671_));
  INV_X1    g470(.A(new_n649_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n285_), .A3(new_n534_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n671_), .A2(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT106), .ZN(G1326gat));
  NOR2_X1   g474(.A1(new_n591_), .A2(new_n592_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G22gat), .B1(new_n661_), .B2(new_n676_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT42), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n672_), .A2(new_n286_), .A3(new_n422_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1327gat));
  INV_X1    g479(.A(new_n333_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n657_), .A2(new_n307_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n648_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(G29gat), .B1(new_n685_), .B2(new_n602_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n333_), .A2(new_n659_), .A3(new_n307_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n267_), .A2(new_n271_), .A3(KEYINPUT107), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(KEYINPUT43), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n691_), .B1(new_n621_), .B2(new_n272_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT33), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n472_), .A2(new_n693_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n583_), .A2(new_n694_), .A3(new_n616_), .A4(new_n609_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n606_), .A2(new_n604_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n696_), .B1(new_n604_), .B2(new_n603_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n695_), .B1(new_n478_), .B2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(new_n676_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n534_), .B1(new_n699_), .B2(new_n593_), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n273_), .B(new_n690_), .C1(new_n700_), .C2(new_n585_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n688_), .B1(new_n692_), .B2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n687_), .B1(new_n702_), .B2(KEYINPUT108), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704_));
  AOI211_X1 g503(.A(new_n704_), .B(new_n688_), .C1(new_n692_), .C2(new_n701_), .ZN(new_n705_));
  OAI21_X1  g504(.A(KEYINPUT109), .B1(new_n703_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n688_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n585_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n584_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n709_));
  AOI22_X1  g508(.A1(new_n709_), .A2(new_n478_), .B1(new_n698_), .B2(new_n676_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n708_), .B1(new_n710_), .B2(new_n534_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n690_), .B1(new_n711_), .B2(new_n273_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n701_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n707_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(new_n704_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n702_), .A2(KEYINPUT108), .ZN(new_n717_));
  NAND4_X1  g516(.A1(new_n715_), .A2(new_n716_), .A3(new_n687_), .A4(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n706_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n702_), .A2(KEYINPUT44), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n602_), .A2(G29gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n686_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  INV_X1    g523(.A(KEYINPUT46), .ZN(new_n725_));
  INV_X1    g524(.A(G36gat), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n720_), .A2(new_n584_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n726_), .B1(new_n719_), .B2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n584_), .A2(new_n726_), .ZN(new_n730_));
  OR3_X1    g529(.A1(new_n684_), .A2(KEYINPUT110), .A3(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT110), .B1(new_n684_), .B2(new_n730_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n725_), .B1(new_n729_), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n733_), .B(KEYINPUT45), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n727_), .B1(new_n706_), .B2(new_n718_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n737_), .B(KEYINPUT46), .C1(new_n738_), .C2(new_n726_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n736_), .A2(new_n739_), .ZN(G1329gat));
  INV_X1    g539(.A(new_n720_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n534_), .A2(G43gat), .ZN(new_n742_));
  AOI211_X1 g541(.A(new_n741_), .B(new_n742_), .C1(new_n706_), .C2(new_n718_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(KEYINPUT111), .B(G43gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n744_), .B1(new_n684_), .B2(new_n620_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT47), .B1(new_n743_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT47), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n748_), .B(new_n745_), .C1(new_n721_), .C2(new_n742_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1330gat));
  AOI21_X1  g549(.A(G50gat), .B1(new_n685_), .B2(new_n422_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n422_), .A2(G50gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n722_), .B2(new_n752_), .ZN(G1331gat));
  NAND4_X1  g552(.A1(new_n658_), .A2(new_n647_), .A3(new_n681_), .A4(new_n660_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G57gat), .B1(new_n754_), .B2(new_n478_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n621_), .A2(new_n659_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n681_), .A3(new_n308_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT112), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n478_), .A2(G57gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n755_), .B1(new_n758_), .B2(new_n759_), .ZN(G1332gat));
  OAI21_X1  g559(.A(G64gat), .B1(new_n754_), .B2(new_n590_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT48), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n590_), .A2(G64gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n758_), .B2(new_n763_), .ZN(G1333gat));
  OAI21_X1  g563(.A(G71gat), .B1(new_n754_), .B2(new_n620_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(KEYINPUT49), .ZN(new_n766_));
  OR2_X1    g565(.A1(new_n620_), .A2(G71gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n766_), .B1(new_n758_), .B2(new_n767_), .ZN(G1334gat));
  OAI21_X1  g567(.A(G78gat), .B1(new_n754_), .B2(new_n676_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT50), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n422_), .A2(new_n400_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n770_), .B1(new_n758_), .B2(new_n771_), .ZN(G1335gat));
  NOR2_X1   g571(.A1(new_n682_), .A2(new_n333_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n756_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(G85gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n602_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n681_), .A2(new_n647_), .A3(new_n307_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n692_), .B2(new_n701_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n779_), .A2(new_n602_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n777_), .B1(new_n780_), .B2(new_n776_), .ZN(G1336gat));
  NOR3_X1   g580(.A1(new_n774_), .A2(G92gat), .A3(new_n590_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n779_), .A2(new_n584_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(G92gat), .B2(new_n783_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(new_n784_), .B(KEYINPUT113), .ZN(G1337gat));
  NAND2_X1  g584(.A1(new_n779_), .A2(new_n534_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n534_), .A2(new_n213_), .ZN(new_n787_));
  AOI22_X1  g586(.A1(new_n786_), .A2(G99gat), .B1(new_n775_), .B2(new_n787_), .ZN(new_n788_));
  XOR2_X1   g587(.A(new_n788_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g588(.A1(new_n775_), .A2(new_n214_), .A3(new_n422_), .ZN(new_n790_));
  AOI211_X1 g589(.A(new_n676_), .B(new_n778_), .C1(new_n692_), .C2(new_n701_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT114), .B1(new_n791_), .B2(new_n214_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n779_), .A2(new_n422_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(G106gat), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT52), .ZN(new_n796_));
  AND3_X1   g595(.A1(new_n792_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n792_), .B2(new_n795_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n790_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT53), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n801_), .B(new_n790_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1339gat));
  INV_X1    g602(.A(new_n657_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n331_), .ZN(new_n805_));
  AND4_X1   g604(.A1(new_n326_), .A2(new_n317_), .A3(new_n324_), .A4(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n644_), .A2(new_n646_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n317_), .A2(new_n324_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT116), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n317_), .A2(new_n324_), .A3(KEYINPUT116), .A4(new_n809_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n313_), .A2(KEYINPUT55), .A3(new_n314_), .A4(new_n316_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n320_), .A2(new_n321_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n316_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n325_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n812_), .A2(new_n813_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n820_), .A2(new_n331_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT56), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT117), .ZN(new_n823_));
  INV_X1    g622(.A(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n821_), .A2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n818_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n805_), .B1(new_n826_), .B2(new_n813_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n823_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n808_), .B1(new_n825_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT119), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n248_), .A2(new_n292_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n632_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n630_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n629_), .A2(KEYINPUT118), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n834_), .A2(new_n835_), .A3(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n640_), .B1(new_n635_), .B2(new_n630_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n830_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n836_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n835_), .B1(new_n629_), .B2(KEYINPUT118), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n838_), .B(new_n830_), .C1(new_n841_), .C2(new_n842_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n843_), .A2(new_n643_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n332_), .A2(new_n840_), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n804_), .B1(new_n829_), .B2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  INV_X1    g648(.A(new_n808_), .ZN(new_n850_));
  AOI211_X1 g649(.A(new_n805_), .B(new_n824_), .C1(new_n826_), .C2(new_n813_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n823_), .B1(new_n820_), .B2(new_n331_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n853_), .A2(new_n845_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n854_), .A2(KEYINPUT57), .A3(new_n804_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n821_), .A2(KEYINPUT56), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n827_), .A2(new_n822_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n843_), .A2(new_n643_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n858_), .A2(new_n839_), .A3(new_n806_), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n856_), .A2(new_n857_), .A3(KEYINPUT58), .A4(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(KEYINPUT121), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n844_), .A2(new_n807_), .A3(new_n840_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(KEYINPUT56), .B2(new_n821_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864_));
  NAND4_X1  g663(.A1(new_n863_), .A2(new_n864_), .A3(KEYINPUT58), .A4(new_n857_), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n861_), .A2(new_n865_), .A3(new_n273_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n859_), .B1(new_n827_), .B2(new_n822_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n821_), .A2(KEYINPUT56), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n867_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n856_), .A2(new_n857_), .A3(KEYINPUT120), .A4(new_n859_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n849_), .B(new_n855_), .C1(new_n866_), .C2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n307_), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n308_), .A2(new_n647_), .A3(new_n333_), .ZN(new_n876_));
  XOR2_X1   g675(.A(KEYINPUT115), .B(KEYINPUT54), .Z(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n478_), .B1(new_n875_), .B2(new_n878_), .ZN(new_n879_));
  NOR3_X1   g678(.A1(new_n422_), .A2(new_n584_), .A3(new_n620_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(KEYINPUT59), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n854_), .B2(new_n804_), .ZN(new_n882_));
  AOI211_X1 g681(.A(new_n848_), .B(new_n657_), .C1(new_n853_), .C2(new_n845_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n870_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n885_), .A2(new_n273_), .A3(new_n861_), .A4(new_n865_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n660_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n878_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n602_), .B(new_n880_), .C1(new_n887_), .C2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT59), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n647_), .B1(new_n881_), .B2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(G113gat), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n659_), .A2(new_n893_), .ZN(new_n894_));
  OAI22_X1  g693(.A1(new_n892_), .A2(new_n893_), .B1(new_n889_), .B2(new_n894_), .ZN(G1340gat));
  AOI21_X1  g694(.A(new_n333_), .B1(new_n881_), .B2(new_n891_), .ZN(new_n896_));
  INV_X1    g695(.A(G120gat), .ZN(new_n897_));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n898_));
  AOI21_X1  g697(.A(G120gat), .B1(new_n681_), .B2(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n899_), .B1(new_n898_), .B2(G120gat), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n889_), .A2(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n902_), .A2(KEYINPUT122), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT122), .ZN(new_n904_));
  NOR3_X1   g703(.A1(new_n889_), .A2(new_n904_), .A3(new_n901_), .ZN(new_n905_));
  OAI22_X1  g704(.A1(new_n896_), .A2(new_n897_), .B1(new_n903_), .B2(new_n905_), .ZN(G1341gat));
  NAND2_X1  g705(.A1(new_n881_), .A2(new_n891_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n307_), .A2(new_n435_), .ZN(new_n908_));
  XNOR2_X1  g707(.A(new_n908_), .B(KEYINPUT123), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n879_), .A2(new_n660_), .A3(new_n880_), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n907_), .A2(new_n909_), .B1(new_n435_), .B2(new_n910_), .ZN(G1342gat));
  AOI21_X1  g710(.A(new_n272_), .B1(new_n881_), .B2(new_n891_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n657_), .A2(new_n433_), .ZN(new_n913_));
  OAI22_X1  g712(.A1(new_n912_), .A2(new_n433_), .B1(new_n889_), .B2(new_n913_), .ZN(G1343gat));
  NAND2_X1  g713(.A1(new_n709_), .A2(new_n620_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n915_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n602_), .B(new_n916_), .C1(new_n887_), .C2(new_n888_), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n917_), .A2(new_n647_), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g718(.A1(new_n917_), .A2(new_n333_), .ZN(new_n920_));
  XOR2_X1   g719(.A(new_n920_), .B(G148gat), .Z(G1345gat));
  OAI21_X1  g720(.A(KEYINPUT124), .B1(new_n917_), .B2(new_n307_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT124), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n879_), .A2(new_n923_), .A3(new_n660_), .A4(new_n916_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT61), .B(G155gat), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n922_), .A2(new_n924_), .A3(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n922_), .B2(new_n924_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1346gat));
  NOR3_X1   g727(.A1(new_n917_), .A2(new_n355_), .A3(new_n272_), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n355_), .B1(new_n917_), .B2(new_n804_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n930_), .A2(KEYINPUT125), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932_));
  OAI211_X1 g731(.A(new_n932_), .B(new_n355_), .C1(new_n917_), .C2(new_n804_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n929_), .B1(new_n931_), .B2(new_n933_), .ZN(G1347gat));
  INV_X1    g733(.A(KEYINPUT126), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n887_), .A2(new_n888_), .ZN(new_n936_));
  NOR3_X1   g735(.A1(new_n422_), .A2(new_n535_), .A3(new_n590_), .ZN(new_n937_));
  INV_X1    g736(.A(new_n937_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n935_), .B1(new_n936_), .B2(new_n938_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n875_), .A2(new_n878_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n940_), .A2(KEYINPUT126), .A3(new_n937_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n939_), .A2(new_n941_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(KEYINPUT22), .B(G169gat), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n942_), .A2(new_n659_), .A3(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT62), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n940_), .A2(new_n659_), .A3(new_n937_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n945_), .B1(new_n946_), .B2(G169gat), .ZN(new_n947_));
  AND3_X1   g746(.A1(new_n946_), .A2(new_n945_), .A3(G169gat), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n944_), .B1(new_n947_), .B2(new_n948_), .ZN(G1348gat));
  NAND3_X1  g748(.A1(new_n942_), .A2(new_n506_), .A3(new_n681_), .ZN(new_n950_));
  NOR3_X1   g749(.A1(new_n936_), .A2(new_n333_), .A3(new_n938_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n506_), .B2(new_n951_), .ZN(G1349gat));
  NOR2_X1   g751(.A1(new_n307_), .A2(new_n513_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n940_), .A2(new_n660_), .A3(new_n937_), .ZN(new_n954_));
  INV_X1    g753(.A(G183gat), .ZN(new_n955_));
  AOI22_X1  g754(.A1(new_n942_), .A2(new_n953_), .B1(new_n954_), .B2(new_n955_), .ZN(G1350gat));
  NAND3_X1  g755(.A1(new_n942_), .A2(new_n509_), .A3(new_n657_), .ZN(new_n957_));
  INV_X1    g756(.A(G190gat), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n272_), .B1(new_n939_), .B2(new_n941_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n957_), .B1(new_n958_), .B2(new_n959_), .ZN(G1351gat));
  NOR4_X1   g759(.A1(new_n676_), .A2(new_n602_), .A3(new_n590_), .A4(new_n534_), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n940_), .A2(new_n961_), .ZN(new_n962_));
  NOR2_X1   g761(.A1(new_n962_), .A2(new_n647_), .ZN(new_n963_));
  XNOR2_X1  g762(.A(new_n963_), .B(new_n335_), .ZN(G1352gat));
  NOR2_X1   g763(.A1(new_n962_), .A2(new_n333_), .ZN(new_n965_));
  XNOR2_X1  g764(.A(new_n965_), .B(new_n337_), .ZN(G1353gat));
  AOI21_X1  g765(.A(new_n307_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n940_), .A2(new_n961_), .A3(new_n967_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n969_));
  XNOR2_X1  g768(.A(new_n969_), .B(KEYINPUT127), .ZN(new_n970_));
  XOR2_X1   g769(.A(new_n968_), .B(new_n970_), .Z(G1354gat));
  OAI21_X1  g770(.A(G218gat), .B1(new_n962_), .B2(new_n272_), .ZN(new_n972_));
  OR2_X1    g771(.A1(new_n804_), .A2(G218gat), .ZN(new_n973_));
  OAI21_X1  g772(.A(new_n972_), .B1(new_n962_), .B2(new_n973_), .ZN(G1355gat));
endmodule


