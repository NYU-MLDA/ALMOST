//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:30 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n829_, new_n830_, new_n831_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n943_, new_n944_, new_n945_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n956_, new_n957_, new_n959_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n966_, new_n967_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n977_, new_n978_, new_n979_, new_n980_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT36), .Z(new_n205_));
  OR2_X1    g004(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n206_));
  INV_X1    g005(.A(G106gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT67), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n213_));
  AND2_X1   g012(.A1(G99gat), .A2(G106gat), .ZN(new_n214_));
  AND3_X1   g013(.A1(new_n211_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n214_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n209_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(G85gat), .B2(G92gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n220_));
  AND2_X1   g019(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n221_));
  AND2_X1   g020(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(KEYINPUT66), .A2(G92gat), .ZN(new_n223_));
  OAI22_X1  g022(.A1(new_n220_), .A2(new_n221_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT9), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n219_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n217_), .A2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G43gat), .B(G50gat), .ZN(new_n228_));
  INV_X1    g027(.A(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(G36gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(G29gat), .ZN(new_n231_));
  INV_X1    g030(.A(G29gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G36gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT71), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n231_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n234_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n229_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n231_), .A2(new_n233_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT71), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(new_n235_), .A3(new_n228_), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n238_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT7), .ZN(new_n243_));
  INV_X1    g042(.A(G99gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n244_), .A3(new_n207_), .ZN(new_n245_));
  OAI21_X1  g044(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n214_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n212_), .A2(KEYINPUT6), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n210_), .A2(KEYINPUT67), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n248_), .B1(new_n249_), .B2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n211_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n247_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  XOR2_X1   g052(.A(G85gat), .B(G92gat), .Z(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NOR3_X1   g054(.A1(new_n253_), .A2(KEYINPUT8), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT8), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n245_), .A2(new_n246_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n258_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n257_), .B1(new_n259_), .B2(new_n254_), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n227_), .B(new_n242_), .C1(new_n256_), .C2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT73), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n217_), .A2(new_n226_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT8), .B1(new_n253_), .B2(new_n255_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n259_), .A2(new_n257_), .A3(new_n254_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT73), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n267_), .A3(new_n242_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n262_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G232gat), .A2(G233gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT35), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n227_), .B1(new_n256_), .B2(new_n260_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n238_), .A2(new_n241_), .ZN(new_n277_));
  XOR2_X1   g076(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n238_), .A2(new_n241_), .A3(new_n278_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n276_), .A2(new_n282_), .B1(new_n273_), .B2(new_n272_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n269_), .A2(new_n275_), .A3(new_n283_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n275_), .B1(new_n269_), .B2(new_n283_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n205_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n261_), .A2(KEYINPUT73), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n267_), .B1(new_n266_), .B2(new_n242_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n283_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n274_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n269_), .A2(new_n275_), .A3(new_n283_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n286_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT100), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G225gat), .A2(G233gat), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G127gat), .B(G134gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(G113gat), .B(G120gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n299_), .B(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  OR2_X1    g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G155gat), .A2(G162gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G141gat), .A2(G148gat), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT3), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT86), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n305_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n306_), .B(KEYINPUT85), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT1), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n303_), .A2(new_n317_), .A3(new_n304_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n304_), .ZN(new_n319_));
  AOI22_X1  g118(.A1(new_n319_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n320_));
  AND3_X1   g119(.A1(new_n316_), .A2(new_n318_), .A3(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n302_), .B1(new_n315_), .B2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n305_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n313_), .B(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n323_), .B1(new_n325_), .B2(new_n311_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n316_), .A2(new_n320_), .A3(new_n318_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n326_), .A2(new_n327_), .A3(new_n301_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n298_), .B1(new_n322_), .B2(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n322_), .A2(KEYINPUT4), .A3(new_n328_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n327_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n332_), .A3(new_n302_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n329_), .B1(new_n334_), .B2(new_n298_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G1gat), .B(G29gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(G85gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(KEYINPUT0), .B(G57gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n296_), .B1(new_n335_), .B2(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n297_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n342_));
  NOR4_X1   g141(.A1(new_n342_), .A2(KEYINPUT100), .A3(new_n339_), .A4(new_n329_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n339_), .B1(new_n342_), .B2(new_n329_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT99), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  OAI211_X1 g146(.A(KEYINPUT99), .B(new_n339_), .C1(new_n342_), .C2(new_n329_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT18), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT32), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G226gat), .A2(G233gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(KEYINPUT19), .ZN(new_n356_));
  INV_X1    g155(.A(new_n356_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G197gat), .B(G204gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT90), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT21), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G211gat), .B(G218gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n359_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT90), .ZN(new_n363_));
  OR2_X1    g162(.A1(G197gat), .A2(G204gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G197gat), .A2(G204gat), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n363_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(G211gat), .B(G218gat), .Z(new_n367_));
  OAI21_X1  g166(.A(KEYINPUT21), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n364_), .A2(KEYINPUT91), .A3(new_n365_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT91), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n361_), .B1(new_n370_), .B2(new_n358_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n362_), .A2(new_n368_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  NOR2_X1   g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G183gat), .A2(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT82), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT82), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(G183gat), .A3(G190gat), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT23), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n375_), .A2(KEYINPUT23), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n374_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G169gat), .A2(G176gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT93), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT22), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(G169gat), .ZN(new_n385_));
  INV_X1    g184(.A(G169gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT22), .ZN(new_n387_));
  INV_X1    g186(.A(G176gat), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n385_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n383_), .A2(KEYINPUT94), .A3(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(KEYINPUT94), .B1(new_n383_), .B2(new_n389_), .ZN(new_n392_));
  OAI211_X1 g191(.A(KEYINPUT95), .B(new_n381_), .C1(new_n391_), .C2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n376_), .A2(new_n378_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n394_), .B1(new_n395_), .B2(KEYINPUT23), .ZN(new_n396_));
  NOR2_X1   g195(.A1(G169gat), .A2(G176gat), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(KEYINPUT24), .A3(new_n382_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT24), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n397_), .A2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT25), .B(G183gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT26), .B(G190gat), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n396_), .A2(new_n399_), .A3(new_n401_), .A4(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n393_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n392_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n407_), .A2(new_n390_), .ZN(new_n408_));
  AOI21_X1  g207(.A(KEYINPUT95), .B1(new_n408_), .B2(new_n381_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n372_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n396_), .A2(new_n374_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n384_), .A2(KEYINPUT83), .A3(G169gat), .ZN(new_n412_));
  AND2_X1   g211(.A1(KEYINPUT83), .A2(G169gat), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n388_), .B(new_n412_), .C1(new_n413_), .C2(new_n384_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(new_n382_), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n379_), .A2(new_n380_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n404_), .A2(new_n399_), .A3(new_n401_), .ZN(new_n417_));
  OAI22_X1  g216(.A1(new_n411_), .A2(new_n415_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT20), .B1(new_n418_), .B2(new_n372_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n357_), .B1(new_n410_), .B2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n381_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT95), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n371_), .A2(new_n369_), .ZN(new_n425_));
  NOR3_X1   g224(.A1(new_n366_), .A2(new_n367_), .A3(KEYINPUT21), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n360_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n425_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n424_), .A2(new_n428_), .A3(new_n405_), .A4(new_n393_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT20), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n430_), .B1(new_n418_), .B2(new_n372_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n429_), .A2(new_n357_), .A3(new_n431_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n421_), .A2(new_n432_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n344_), .A2(new_n349_), .B1(new_n354_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT98), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n428_), .A2(KEYINPUT92), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT92), .ZN(new_n437_));
  OAI211_X1 g236(.A(new_n437_), .B(new_n425_), .C1(new_n426_), .C2(new_n427_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n436_), .A2(new_n422_), .A3(new_n405_), .A4(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n431_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n356_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n410_), .A2(new_n420_), .A3(new_n357_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n435_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n424_), .A2(new_n405_), .A3(new_n393_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n419_), .B1(new_n444_), .B2(new_n372_), .ZN(new_n445_));
  AOI21_X1  g244(.A(KEYINPUT98), .B1(new_n445_), .B2(new_n357_), .ZN(new_n446_));
  OAI211_X1 g245(.A(KEYINPUT32), .B(new_n353_), .C1(new_n443_), .C2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n434_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n353_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(new_n421_), .B2(new_n432_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n429_), .A2(new_n431_), .A3(new_n357_), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n353_), .B(new_n451_), .C1(new_n445_), .C2(new_n357_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT96), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT96), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n450_), .A2(new_n455_), .A3(new_n452_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n330_), .A2(new_n297_), .A3(new_n333_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n322_), .A2(new_n298_), .A3(new_n328_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n457_), .A2(new_n340_), .A3(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT97), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n457_), .A2(KEYINPUT97), .A3(new_n340_), .A4(new_n458_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n345_), .A2(KEYINPUT33), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT33), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n465_), .B(new_n339_), .C1(new_n342_), .C2(new_n329_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  NAND4_X1  g266(.A1(new_n454_), .A2(new_n456_), .A3(new_n463_), .A4(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n448_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n331_), .A2(KEYINPUT29), .ZN(new_n470_));
  NAND2_X1  g269(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n473_));
  OAI21_X1  g272(.A(G228gat), .B1(new_n472_), .B2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n470_), .A2(new_n372_), .A3(new_n474_), .ZN(new_n475_));
  AOI22_X1  g274(.A1(new_n436_), .A2(new_n438_), .B1(KEYINPUT29), .B2(new_n331_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n475_), .B1(new_n476_), .B2(new_n474_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT29), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n326_), .A2(new_n327_), .A3(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(KEYINPUT88), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n479_), .B(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n477_), .A2(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G22gat), .B(G50gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G78gat), .B(G106gat), .ZN(new_n486_));
  XOR2_X1   g285(.A(new_n485_), .B(new_n486_), .Z(new_n487_));
  OAI211_X1 g286(.A(new_n482_), .B(new_n475_), .C1(new_n476_), .C2(new_n474_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n484_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n487_), .B1(new_n484_), .B2(new_n488_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  OAI221_X1 g290(.A(KEYINPUT30), .B1(new_n416_), .B2(new_n417_), .C1(new_n411_), .C2(new_n415_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G227gat), .A2(G233gat), .ZN(new_n493_));
  INV_X1    g292(.A(G15gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(G71gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n496_), .A2(G99gat), .ZN(new_n497_));
  INV_X1    g296(.A(G71gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n495_), .B(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n244_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n497_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT30), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n415_), .B1(new_n374_), .B2(new_n396_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n417_), .A2(new_n416_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n502_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n492_), .A2(new_n501_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n501_), .B1(new_n505_), .B2(new_n492_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n302_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n492_), .A2(new_n505_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n501_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n492_), .A2(new_n501_), .A3(new_n505_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n301_), .A3(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(KEYINPUT84), .B(G43gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT31), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n508_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n515_), .B1(new_n508_), .B2(new_n513_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n491_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n469_), .A2(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n508_), .A2(new_n513_), .A3(new_n515_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n508_), .A2(new_n513_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n515_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  OAI211_X1 g324(.A(new_n522_), .B(new_n525_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n487_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n372_), .A2(new_n437_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n438_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n470_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n474_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n482_), .B1(new_n532_), .B2(new_n475_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n488_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n527_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n484_), .A2(new_n487_), .A3(new_n488_), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n535_), .B(new_n536_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n526_), .A2(new_n537_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n344_), .A2(new_n349_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n449_), .B1(new_n443_), .B2(new_n446_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n452_), .A2(KEYINPUT27), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT27), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n540_), .A2(new_n541_), .B1(new_n453_), .B2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n538_), .A2(new_n539_), .A3(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n295_), .B1(new_n521_), .B2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G120gat), .B(G148gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT5), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G176gat), .B(G204gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(new_n548_), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G230gat), .A2(G233gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT64), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(G64gat), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n554_), .A2(G57gat), .ZN(new_n555_));
  INV_X1    g354(.A(G57gat), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(G64gat), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n555_), .A2(new_n557_), .A3(KEYINPUT68), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(KEYINPUT68), .B1(new_n555_), .B2(new_n557_), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT11), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n555_), .A2(new_n557_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT68), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT11), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n565_), .A3(new_n558_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G71gat), .B(G78gat), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n561_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(KEYINPUT11), .B(new_n567_), .C1(new_n559_), .C2(new_n560_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n276_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n264_), .A2(new_n265_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n570_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n574_), .A3(new_n227_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n572_), .A2(KEYINPUT12), .A3(new_n575_), .ZN(new_n576_));
  OR3_X1    g375(.A1(new_n266_), .A2(KEYINPUT12), .A3(new_n574_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n553_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n552_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n550_), .B1(new_n579_), .B2(new_n581_), .ZN(new_n582_));
  NOR3_X1   g381(.A1(new_n578_), .A2(new_n580_), .A3(new_n549_), .ZN(new_n583_));
  XOR2_X1   g382(.A(KEYINPUT69), .B(KEYINPUT13), .Z(new_n584_));
  NOR3_X1   g383(.A1(new_n582_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  OAI22_X1  g385(.A1(new_n582_), .A2(new_n583_), .B1(KEYINPUT69), .B2(KEYINPUT13), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G15gat), .B(G22gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(KEYINPUT76), .B(G1gat), .ZN(new_n590_));
  INV_X1    g389(.A(G8gat), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT14), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n589_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G1gat), .B(G8gat), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n596_), .ZN(new_n597_));
  OAI211_X1 g396(.A(new_n589_), .B(new_n595_), .C1(new_n592_), .C2(new_n593_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n282_), .A2(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n242_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n601_), .A2(new_n602_), .A3(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n597_), .A2(new_n277_), .A3(new_n598_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n602_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n603_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT80), .B1(new_n606_), .B2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT80), .ZN(new_n609_));
  AOI211_X1 g408(.A(new_n609_), .B(new_n603_), .C1(new_n602_), .C2(new_n605_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n604_), .B1(new_n608_), .B2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(G113gat), .B(G141gat), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n612_), .B(KEYINPUT81), .ZN(new_n613_));
  XNOR2_X1  g412(.A(G169gat), .B(G197gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n613_), .B(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n611_), .A2(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n615_), .ZN(new_n617_));
  OAI211_X1 g416(.A(new_n604_), .B(new_n617_), .C1(new_n608_), .C2(new_n610_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n588_), .A2(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT77), .Z(new_n622_));
  XNOR2_X1  g421(.A(G127gat), .B(G155gat), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT16), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G183gat), .B(G211gat), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n624_), .A2(new_n625_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT17), .ZN(new_n629_));
  OAI21_X1  g428(.A(KEYINPUT78), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n630_), .A2(new_n600_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n600_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(new_n571_), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n571_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n622_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n635_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n622_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(new_n633_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n628_), .A2(new_n629_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n636_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n620_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n545_), .A2(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(KEYINPUT102), .ZN(new_n645_));
  INV_X1    g444(.A(new_n539_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT37), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n286_), .A2(new_n293_), .A3(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n649_), .A2(KEYINPUT75), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT74), .ZN(new_n651_));
  OAI211_X1 g450(.A(new_n651_), .B(new_n205_), .C1(new_n284_), .C2(new_n285_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n652_), .A2(new_n293_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n290_), .A2(new_n291_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n651_), .B1(new_n654_), .B2(new_n205_), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT37), .B1(new_n653_), .B2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n650_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT75), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n658_), .B(KEYINPUT37), .C1(new_n653_), .C2(new_n655_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n657_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(new_n642_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT79), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n620_), .B1(new_n521_), .B2(new_n544_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n539_), .B(KEYINPUT101), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AND4_X1   g464(.A1(new_n590_), .A2(new_n662_), .A3(new_n663_), .A4(new_n665_), .ZN(new_n666_));
  AOI22_X1  g465(.A1(G1gat), .A2(new_n647_), .B1(new_n666_), .B2(KEYINPUT38), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(KEYINPUT38), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(KEYINPUT103), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT103), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n666_), .A2(new_n670_), .A3(KEYINPUT38), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n667_), .B1(new_n669_), .B2(new_n671_), .ZN(G1324gat));
  INV_X1    g471(.A(KEYINPUT39), .ZN(new_n673_));
  INV_X1    g472(.A(new_n644_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n543_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n673_), .B1(new_n676_), .B2(G8gat), .ZN(new_n677_));
  AOI211_X1 g476(.A(KEYINPUT39), .B(new_n591_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n662_), .A2(new_n663_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n675_), .A2(new_n591_), .ZN(new_n680_));
  OAI22_X1  g479(.A1(new_n677_), .A2(new_n678_), .B1(new_n679_), .B2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT40), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(G1325gat));
  INV_X1    g482(.A(new_n679_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n518_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n494_), .A3(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n645_), .A2(new_n685_), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n687_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT41), .B1(new_n687_), .B2(G15gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n686_), .B1(new_n688_), .B2(new_n689_), .ZN(G1326gat));
  INV_X1    g489(.A(G22gat), .ZN(new_n691_));
  INV_X1    g490(.A(new_n491_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n684_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n645_), .A2(new_n692_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n694_), .B1(new_n695_), .B2(G22gat), .ZN(new_n696_));
  AOI211_X1 g495(.A(KEYINPUT42), .B(new_n691_), .C1(new_n645_), .C2(new_n692_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n693_), .B1(new_n696_), .B2(new_n697_), .ZN(G1327gat));
  NOR2_X1   g497(.A1(new_n641_), .A2(new_n294_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT106), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n663_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G29gat), .B1(new_n702_), .B2(new_n646_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n467_), .A2(new_n463_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n455_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AOI22_X1  g505(.A1(new_n706_), .A2(new_n456_), .B1(new_n434_), .B2(new_n447_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n544_), .B1(new_n707_), .B2(new_n519_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT43), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(new_n709_), .A3(new_n660_), .ZN(new_n710_));
  AOI22_X1  g509(.A1(new_n521_), .A2(new_n544_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(KEYINPUT104), .B(KEYINPUT43), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n710_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n620_), .A2(new_n641_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT44), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  AND3_X1   g515(.A1(new_n708_), .A2(new_n709_), .A3(new_n660_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n713_), .B1(new_n708_), .B2(new_n660_), .ZN(new_n718_));
  OAI211_X1 g517(.A(KEYINPUT44), .B(new_n715_), .C1(new_n717_), .C2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n714_), .A2(KEYINPUT105), .A3(KEYINPUT44), .A4(new_n715_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n716_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n664_), .A2(new_n232_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n703_), .B1(new_n723_), .B2(new_n724_), .ZN(G1328gat));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n721_), .A2(new_n722_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n716_), .A2(new_n543_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n230_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n543_), .A2(G36gat), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(KEYINPUT107), .B1(new_n701_), .B2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT107), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n663_), .A2(new_n733_), .A3(new_n700_), .A4(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT45), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n732_), .A2(KEYINPUT45), .A3(new_n734_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n726_), .B1(new_n729_), .B2(new_n739_), .ZN(new_n740_));
  AND3_X1   g539(.A1(new_n732_), .A2(KEYINPUT45), .A3(new_n734_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT45), .B1(new_n732_), .B2(new_n734_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n715_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n708_), .A2(new_n660_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n712_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n746_), .B2(new_n710_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n675_), .B1(new_n747_), .B2(KEYINPUT44), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n749_));
  OAI211_X1 g548(.A(new_n743_), .B(KEYINPUT46), .C1(new_n749_), .C2(new_n230_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n740_), .A2(new_n750_), .ZN(G1329gat));
  INV_X1    g550(.A(G43gat), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n518_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n754_), .B(new_n716_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n752_), .B1(new_n701_), .B2(new_n518_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  OAI21_X1  g556(.A(KEYINPUT47), .B1(new_n755_), .B2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n723_), .A2(new_n753_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(new_n756_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n758_), .A2(new_n761_), .ZN(G1330gat));
  AOI21_X1  g561(.A(G50gat), .B1(new_n702_), .B2(new_n692_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n692_), .A2(G50gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n723_), .B2(new_n764_), .ZN(G1331gat));
  NOR2_X1   g564(.A1(new_n588_), .A2(new_n619_), .ZN(new_n766_));
  AND2_X1   g565(.A1(new_n708_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n662_), .A2(new_n767_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n556_), .B1(new_n768_), .B2(new_n664_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n545_), .A2(new_n641_), .A3(new_n766_), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n770_), .A2(KEYINPUT108), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(KEYINPUT108), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(KEYINPUT109), .A2(G57gat), .ZN(new_n774_));
  AND2_X1   g573(.A1(KEYINPUT109), .A2(G57gat), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n646_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n769_), .B1(new_n773_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n769_), .B(KEYINPUT110), .C1(new_n773_), .C2(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1332gat));
  INV_X1    g580(.A(new_n768_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n782_), .A2(new_n554_), .A3(new_n675_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n771_), .A2(new_n675_), .A3(new_n772_), .ZN(new_n784_));
  XNOR2_X1  g583(.A(KEYINPUT111), .B(KEYINPUT48), .ZN(new_n785_));
  AND3_X1   g584(.A1(new_n784_), .A2(G64gat), .A3(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n785_), .B1(new_n784_), .B2(G64gat), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n783_), .B1(new_n786_), .B2(new_n787_), .ZN(G1333gat));
  NAND3_X1  g587(.A1(new_n782_), .A2(new_n498_), .A3(new_n685_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n771_), .A2(new_n685_), .A3(new_n772_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n790_), .A2(new_n791_), .A3(G71gat), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n791_), .B1(new_n790_), .B2(G71gat), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(G1334gat));
  OR3_X1    g593(.A1(new_n768_), .A2(G78gat), .A3(new_n491_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n771_), .A2(new_n692_), .A3(new_n772_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n797_));
  AND3_X1   g596(.A1(new_n796_), .A2(new_n797_), .A3(G78gat), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n796_), .B2(G78gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n795_), .B1(new_n798_), .B2(new_n799_), .ZN(G1335gat));
  AND2_X1   g599(.A1(new_n767_), .A2(new_n700_), .ZN(new_n801_));
  AOI21_X1  g600(.A(G85gat), .B1(new_n801_), .B2(new_n665_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT112), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n714_), .A2(new_n803_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n746_), .A2(KEYINPUT112), .A3(new_n710_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n588_), .A2(new_n619_), .A3(new_n641_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n804_), .A2(new_n805_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  OR2_X1    g607(.A1(new_n221_), .A2(new_n220_), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n646_), .A2(new_n809_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n802_), .B1(new_n808_), .B2(new_n810_), .ZN(G1336gat));
  AOI21_X1  g610(.A(G92gat), .B1(new_n801_), .B2(new_n675_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n222_), .A2(new_n223_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n543_), .A2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n812_), .B1(new_n808_), .B2(new_n814_), .ZN(G1337gat));
  OAI21_X1  g614(.A(G99gat), .B1(new_n807_), .B2(new_n518_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n801_), .A2(new_n206_), .A3(new_n208_), .A4(new_n685_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT51), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n816_), .A2(new_n820_), .A3(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1338gat));
  NAND3_X1  g621(.A1(new_n801_), .A2(new_n207_), .A3(new_n692_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n714_), .A2(new_n692_), .A3(new_n806_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n824_), .A2(new_n825_), .A3(G106gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n824_), .B2(G106gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n823_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT53), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n823_), .B(new_n830_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(G1339gat));
  AOI21_X1  g631(.A(new_n619_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n833_), .A2(new_n657_), .A3(new_n659_), .A4(new_n641_), .ZN(new_n834_));
  XNOR2_X1  g633(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n834_), .B(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n583_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n619_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n576_), .A2(new_n577_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(KEYINPUT55), .A3(new_n552_), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n576_), .A2(new_n577_), .A3(new_n553_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  XOR2_X1   g642(.A(KEYINPUT114), .B(KEYINPUT55), .Z(new_n844_));
  NOR2_X1   g643(.A1(new_n578_), .A2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n549_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT56), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n841_), .B(new_n842_), .C1(new_n578_), .C2(new_n844_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n849_), .A2(KEYINPUT56), .A3(new_n549_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n839_), .B1(new_n848_), .B2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n582_), .A2(new_n583_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n601_), .A2(new_n602_), .A3(new_n607_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n606_), .A2(new_n603_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n854_), .A3(new_n615_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n618_), .A2(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n852_), .A2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n294_), .B1(new_n851_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT115), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861_));
  OAI211_X1 g660(.A(KEYINPUT115), .B(new_n294_), .C1(new_n851_), .C2(new_n857_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n295_), .A2(new_n861_), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n864_), .B1(new_n851_), .B2(new_n857_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT117), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n867_), .B(new_n864_), .C1(new_n851_), .C2(new_n857_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n838_), .A2(KEYINPUT116), .A3(new_n618_), .A4(new_n855_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT116), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n856_), .B2(new_n583_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n850_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT56), .B1(new_n849_), .B2(new_n549_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT58), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n876_), .A2(new_n877_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n873_), .B(KEYINPUT58), .C1(new_n875_), .C2(new_n874_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n863_), .A2(new_n869_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n837_), .B1(new_n881_), .B2(new_n642_), .ZN(new_n882_));
  OR3_X1    g681(.A1(new_n664_), .A2(new_n675_), .A3(new_n537_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(KEYINPUT118), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n882_), .A2(new_n885_), .ZN(new_n886_));
  AOI21_X1  g685(.A(G113gat), .B1(new_n886_), .B2(new_n619_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT59), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n888_), .B1(new_n882_), .B2(new_n885_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n866_), .A2(new_n868_), .B1(new_n878_), .B2(new_n879_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n641_), .B1(new_n890_), .B2(new_n863_), .ZN(new_n891_));
  OAI211_X1 g690(.A(KEYINPUT59), .B(new_n884_), .C1(new_n891_), .C2(new_n837_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n889_), .A2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n619_), .A2(G113gat), .ZN(new_n894_));
  XOR2_X1   g693(.A(new_n894_), .B(KEYINPUT119), .Z(new_n895_));
  AOI21_X1  g694(.A(new_n887_), .B1(new_n893_), .B2(new_n895_), .ZN(G1340gat));
  XNOR2_X1  g695(.A(KEYINPUT120), .B(G120gat), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n588_), .B2(KEYINPUT60), .ZN(new_n898_));
  OAI211_X1 g697(.A(new_n886_), .B(new_n898_), .C1(KEYINPUT60), .C2(new_n897_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n588_), .B1(new_n889_), .B2(new_n892_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n900_), .B2(new_n897_), .ZN(G1341gat));
  INV_X1    g700(.A(G127gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n886_), .A2(new_n902_), .A3(new_n641_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n642_), .B1(new_n889_), .B2(new_n892_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n902_), .ZN(G1342gat));
  OAI211_X1 g704(.A(new_n295_), .B(new_n884_), .C1(new_n891_), .C2(new_n837_), .ZN(new_n906_));
  INV_X1    g705(.A(G134gat), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT121), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n906_), .A2(KEYINPUT121), .A3(new_n907_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n660_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n907_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n910_), .A2(new_n911_), .B1(new_n893_), .B2(new_n913_), .ZN(G1343gat));
  NAND2_X1  g713(.A1(new_n881_), .A2(new_n642_), .ZN(new_n915_));
  INV_X1    g714(.A(new_n837_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n664_), .A2(new_n675_), .A3(new_n526_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n917_), .A2(new_n619_), .A3(new_n918_), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n919_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g719(.A(new_n588_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n917_), .A2(new_n921_), .A3(new_n918_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g722(.A1(new_n917_), .A2(new_n641_), .A3(new_n918_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT61), .B(G155gat), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n924_), .B(new_n925_), .ZN(G1346gat));
  NAND2_X1  g725(.A1(new_n917_), .A2(new_n918_), .ZN(new_n927_));
  OAI21_X1  g726(.A(G162gat), .B1(new_n927_), .B2(new_n912_), .ZN(new_n928_));
  INV_X1    g727(.A(G162gat), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n295_), .A2(new_n929_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n928_), .B1(new_n927_), .B2(new_n930_), .ZN(G1347gat));
  AND3_X1   g730(.A1(new_n664_), .A2(new_n685_), .A3(new_n675_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n619_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n933_), .B(new_n934_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n935_), .B(new_n491_), .C1(new_n891_), .C2(new_n837_), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT62), .ZN(new_n937_));
  AND3_X1   g736(.A1(new_n936_), .A2(new_n937_), .A3(G169gat), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n937_), .B1(new_n936_), .B2(G169gat), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n491_), .B(new_n932_), .C1(new_n891_), .C2(new_n837_), .ZN(new_n940_));
  NAND3_X1  g739(.A1(new_n619_), .A2(new_n385_), .A3(new_n387_), .ZN(new_n941_));
  OAI22_X1  g740(.A1(new_n938_), .A2(new_n939_), .B1(new_n940_), .B2(new_n941_), .ZN(G1348gat));
  NOR2_X1   g741(.A1(new_n882_), .A2(new_n692_), .ZN(new_n943_));
  NAND4_X1  g742(.A1(new_n943_), .A2(G176gat), .A3(new_n921_), .A4(new_n932_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n388_), .B1(new_n940_), .B2(new_n588_), .ZN(new_n945_));
  AND2_X1   g744(.A1(new_n944_), .A2(new_n945_), .ZN(G1349gat));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n947_));
  INV_X1    g746(.A(new_n402_), .ZN(new_n948_));
  AND2_X1   g747(.A1(new_n932_), .A2(new_n641_), .ZN(new_n949_));
  NAND4_X1  g748(.A1(new_n943_), .A2(new_n947_), .A3(new_n948_), .A4(new_n949_), .ZN(new_n950_));
  OAI211_X1 g749(.A(new_n491_), .B(new_n949_), .C1(new_n891_), .C2(new_n837_), .ZN(new_n951_));
  OAI21_X1  g750(.A(KEYINPUT123), .B1(new_n951_), .B2(new_n402_), .ZN(new_n952_));
  INV_X1    g751(.A(G183gat), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n951_), .A2(new_n953_), .ZN(new_n954_));
  AND3_X1   g753(.A1(new_n950_), .A2(new_n952_), .A3(new_n954_), .ZN(G1350gat));
  OAI21_X1  g754(.A(G190gat), .B1(new_n940_), .B2(new_n912_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n295_), .A2(new_n403_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n940_), .B2(new_n957_), .ZN(G1351gat));
  OR3_X1    g757(.A1(new_n646_), .A2(KEYINPUT124), .A3(new_n526_), .ZN(new_n959_));
  OAI21_X1  g758(.A(KEYINPUT124), .B1(new_n646_), .B2(new_n526_), .ZN(new_n960_));
  AND3_X1   g759(.A1(new_n959_), .A2(new_n675_), .A3(new_n960_), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n917_), .A2(new_n619_), .A3(new_n961_), .ZN(new_n962_));
  XNOR2_X1  g761(.A(KEYINPUT125), .B(G197gat), .ZN(new_n963_));
  INV_X1    g762(.A(new_n963_), .ZN(new_n964_));
  XNOR2_X1  g763(.A(new_n962_), .B(new_n964_), .ZN(G1352gat));
  NAND3_X1  g764(.A1(new_n917_), .A2(new_n921_), .A3(new_n961_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(KEYINPUT126), .B(G204gat), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n966_), .B(new_n967_), .ZN(G1353gat));
  AOI21_X1  g767(.A(new_n642_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n969_));
  OAI211_X1 g768(.A(new_n961_), .B(new_n969_), .C1(new_n891_), .C2(new_n837_), .ZN(new_n970_));
  NOR3_X1   g769(.A1(KEYINPUT127), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n971_));
  NOR2_X1   g770(.A1(new_n970_), .A2(new_n971_), .ZN(new_n972_));
  INV_X1    g771(.A(new_n971_), .ZN(new_n973_));
  OAI21_X1  g772(.A(KEYINPUT127), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n973_), .A2(new_n974_), .ZN(new_n975_));
  AOI21_X1  g774(.A(new_n972_), .B1(new_n970_), .B2(new_n975_), .ZN(G1354gat));
  NAND2_X1  g775(.A1(new_n917_), .A2(new_n961_), .ZN(new_n977_));
  OAI21_X1  g776(.A(G218gat), .B1(new_n977_), .B2(new_n912_), .ZN(new_n978_));
  INV_X1    g777(.A(G218gat), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n295_), .A2(new_n979_), .ZN(new_n980_));
  OAI21_X1  g779(.A(new_n978_), .B1(new_n977_), .B2(new_n980_), .ZN(G1355gat));
endmodule


