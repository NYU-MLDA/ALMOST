//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n899_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n921_, new_n922_,
    new_n923_, new_n924_;
  XNOR2_X1  g000(.A(G190gat), .B(G218gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n204_), .B(KEYINPUT36), .Z(new_n205_));
  INV_X1    g004(.A(KEYINPUT66), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NOR3_X1   g007(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(new_n206_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G99gat), .ZN(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT6), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n213_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT7), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(KEYINPUT66), .A3(new_n207_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n210_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G85gat), .ZN(new_n221_));
  INV_X1    g020(.A(G92gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G85gat), .A2(G92gat), .ZN(new_n224_));
  AND2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n220_), .A2(KEYINPUT67), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT8), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT67), .B1(new_n220_), .B2(new_n225_), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT68), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n220_), .A2(new_n225_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n232_), .A2(new_n233_), .A3(KEYINPUT8), .A4(new_n226_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n216_), .A2(new_n218_), .A3(new_n207_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT8), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n225_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT65), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n229_), .A2(new_n234_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT9), .ZN(new_n241_));
  AND3_X1   g040(.A1(new_n224_), .A2(KEYINPUT64), .A3(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(KEYINPUT64), .B1(new_n224_), .B2(new_n241_), .ZN(new_n243_));
  OAI221_X1 g042(.A(new_n223_), .B1(new_n241_), .B2(new_n224_), .C1(new_n242_), .C2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT10), .B(G99gat), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n244_), .B(new_n216_), .C1(G106gat), .C2(new_n245_), .ZN(new_n246_));
  AND3_X1   g045(.A1(new_n240_), .A2(KEYINPUT71), .A3(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT71), .B1(new_n240_), .B2(new_n246_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G43gat), .B(G50gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G29gat), .B(G36gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT73), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  NOR2_X1   g054(.A1(new_n252_), .A2(new_n253_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n251_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G29gat), .B(G36gat), .Z(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT73), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n259_), .A2(new_n254_), .A3(new_n250_), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n257_), .A2(KEYINPUT15), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT15), .B1(new_n257_), .B2(new_n260_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n249_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G232gat), .A2(G233gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT35), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n240_), .A2(new_n246_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NOR3_X1   g070(.A1(new_n255_), .A2(new_n256_), .A3(new_n251_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n250_), .B1(new_n259_), .B2(new_n254_), .ZN(new_n273_));
  NOR2_X1   g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  AOI22_X1  g073(.A1(new_n271_), .A2(new_n274_), .B1(new_n267_), .B2(new_n266_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n263_), .A2(new_n269_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n269_), .B1(new_n263_), .B2(new_n275_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n205_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n278_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n204_), .A2(KEYINPUT36), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n280_), .A2(new_n281_), .A3(new_n276_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n279_), .A2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n283_), .A2(KEYINPUT37), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT37), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n285_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n284_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G15gat), .B(G22gat), .ZN(new_n288_));
  INV_X1    g087(.A(G1gat), .ZN(new_n289_));
  INV_X1    g088(.A(G8gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT14), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G1gat), .B(G8gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G231gat), .A2(G233gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n295_), .B(KEYINPUT74), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n294_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G57gat), .B(G64gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(KEYINPUT11), .ZN(new_n300_));
  XOR2_X1   g099(.A(G71gat), .B(G78gat), .Z(new_n301_));
  OR2_X1    g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n300_), .A2(new_n301_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n299_), .A2(KEYINPUT11), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT75), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n298_), .A2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G127gat), .B(G155gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G183gat), .B(G211gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n312_), .A2(KEYINPUT17), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n298_), .A2(new_n306_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n307_), .A2(new_n313_), .A3(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT77), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n312_), .A2(KEYINPUT17), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n305_), .B(KEYINPUT69), .Z(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI211_X1 g118(.A(new_n317_), .B(new_n313_), .C1(new_n319_), .C2(new_n298_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n320_), .B1(new_n319_), .B2(new_n298_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n316_), .A2(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n287_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT78), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT71), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n270_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n240_), .A2(KEYINPUT71), .A3(new_n246_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n305_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT12), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n326_), .A2(new_n327_), .A3(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n240_), .A2(new_n246_), .A3(new_n318_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(KEYINPUT12), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n270_), .A2(new_n319_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G230gat), .A2(G233gat), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n331_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n336_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n332_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n318_), .B1(new_n240_), .B2(new_n246_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT70), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OAI211_X1 g142(.A(KEYINPUT70), .B(new_n338_), .C1(new_n339_), .C2(new_n340_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n337_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G120gat), .B(G148gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT5), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G176gat), .B(G204gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  AND2_X1   g148(.A1(new_n345_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n349_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n337_), .A2(new_n343_), .A3(new_n344_), .A4(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n350_), .A2(new_n353_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n354_), .A2(KEYINPUT13), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(KEYINPUT13), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n324_), .A2(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT87), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT1), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n364_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(G141gat), .ZN(new_n369_));
  INV_X1    g168(.A(G148gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(G141gat), .A2(G148gat), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n368_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT88), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT3), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT2), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n378_), .B(new_n379_), .C1(new_n380_), .C2(new_n372_), .ZN(new_n381_));
  OAI211_X1 g180(.A(new_n364_), .B(new_n365_), .C1(new_n376_), .C2(new_n381_), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n373_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT29), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT89), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n385_), .B(KEYINPUT89), .ZN(new_n390_));
  INV_X1    g189(.A(new_n388_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  XOR2_X1   g191(.A(G22gat), .B(G50gat), .Z(new_n393_));
  AND3_X1   g192(.A1(new_n389_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n393_), .B1(new_n389_), .B2(new_n392_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(G78gat), .B(G106gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT21), .ZN(new_n398_));
  XNOR2_X1  g197(.A(G211gat), .B(G218gat), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n399_), .A2(KEYINPUT92), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(KEYINPUT92), .ZN(new_n401_));
  XOR2_X1   g200(.A(G197gat), .B(G204gat), .Z(new_n402_));
  OR3_X1    g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT91), .ZN(new_n404_));
  OAI22_X1  g203(.A1(new_n400_), .A2(new_n401_), .B1(new_n404_), .B2(new_n402_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n398_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n405_), .A2(new_n398_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n384_), .B2(new_n383_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n409_), .A2(new_n411_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n397_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  OAI22_X1  g213(.A1(new_n394_), .A2(new_n395_), .B1(new_n414_), .B2(KEYINPUT93), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(KEYINPUT94), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT94), .ZN(new_n417_));
  INV_X1    g216(.A(new_n393_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n390_), .A2(new_n391_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n387_), .A2(new_n388_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n418_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n389_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n409_), .B(new_n411_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n396_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT93), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n417_), .B1(new_n423_), .B2(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n424_), .A2(new_n396_), .ZN(new_n429_));
  OAI22_X1  g228(.A1(new_n416_), .A2(new_n428_), .B1(new_n414_), .B2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n415_), .A2(KEYINPUT94), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n429_), .A2(new_n414_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n423_), .A2(new_n427_), .A3(new_n417_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n431_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n373_), .A2(new_n382_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G127gat), .B(G134gat), .Z(new_n437_));
  XOR2_X1   g236(.A(G113gat), .B(G120gat), .Z(new_n438_));
  XOR2_X1   g237(.A(new_n437_), .B(new_n438_), .Z(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(KEYINPUT4), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(KEYINPUT98), .B1(new_n436_), .B2(new_n439_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(new_n440_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT4), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n442_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G225gat), .A2(G233gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n446_), .A2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n447_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  XOR2_X1   g250(.A(G1gat), .B(G29gat), .Z(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT99), .B(KEYINPUT0), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G57gat), .B(G85gat), .ZN(new_n455_));
  XOR2_X1   g254(.A(new_n454_), .B(new_n455_), .Z(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n451_), .A2(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n449_), .A2(new_n456_), .A3(new_n450_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G183gat), .A2(G190gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT23), .ZN(new_n463_));
  OR2_X1    g262(.A1(G183gat), .A2(G190gat), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G169gat), .A2(G176gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT22), .B(G169gat), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n466_), .B1(new_n468_), .B2(G176gat), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n465_), .B1(KEYINPUT84), .B2(new_n469_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(KEYINPUT84), .B2(new_n469_), .ZN(new_n471_));
  OR2_X1    g270(.A1(G169gat), .A2(G176gat), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n472_), .A2(KEYINPUT24), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(KEYINPUT24), .A3(new_n466_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n463_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(KEYINPUT26), .B(G190gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT25), .B(G183gat), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n475_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n471_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G71gat), .B(G99gat), .ZN(new_n481_));
  INV_X1    g280(.A(G43gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n481_), .B(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n480_), .B(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(G227gat), .A2(G233gat), .ZN(new_n486_));
  INV_X1    g285(.A(G15gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT30), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT31), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NOR2_X1   g291(.A1(new_n485_), .A2(new_n490_), .ZN(new_n493_));
  OAI21_X1  g292(.A(KEYINPUT85), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  OR2_X1    g293(.A1(new_n485_), .A2(new_n490_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT85), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(new_n496_), .A3(new_n491_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n494_), .A2(new_n439_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n439_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n461_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n465_), .A2(new_n469_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n477_), .B(KEYINPUT96), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n476_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n503_), .B1(new_n475_), .B2(new_n505_), .ZN(new_n506_));
  OR3_X1    g305(.A1(new_n506_), .A2(new_n406_), .A3(new_n407_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n507_), .B(KEYINPUT20), .C1(new_n408_), .C2(new_n480_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G226gat), .A2(G233gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n506_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT97), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n514_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n480_), .A2(new_n408_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n511_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n518_), .A2(KEYINPUT20), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .A4(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G8gat), .B(G36gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT18), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G64gat), .B(G92gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n522_), .B(new_n523_), .Z(new_n524_));
  NAND3_X1  g323(.A1(new_n512_), .A2(new_n520_), .A3(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n525_), .A2(KEYINPUT102), .ZN(new_n526_));
  INV_X1    g325(.A(new_n524_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n508_), .A2(new_n511_), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n513_), .A2(KEYINPUT20), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n518_), .B1(new_n529_), .B2(new_n517_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n527_), .B1(new_n528_), .B2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n526_), .A2(new_n531_), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n525_), .A2(KEYINPUT102), .ZN(new_n533_));
  OAI21_X1  g332(.A(KEYINPUT27), .B1(new_n532_), .B2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n512_), .A2(new_n520_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(new_n527_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT27), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n525_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n534_), .A2(new_n538_), .ZN(new_n539_));
  AND3_X1   g338(.A1(new_n435_), .A2(new_n502_), .A3(new_n539_), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n539_), .A2(new_n430_), .A3(new_n461_), .A4(new_n434_), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n444_), .A2(new_n447_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n542_), .B(new_n456_), .C1(new_n446_), .C2(new_n448_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n536_), .A2(new_n543_), .A3(new_n525_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT101), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT33), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n458_), .A2(new_n545_), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n456_), .B1(new_n449_), .B2(new_n450_), .ZN(new_n548_));
  OAI21_X1  g347(.A(KEYINPUT101), .B1(new_n548_), .B2(KEYINPUT33), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n544_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT100), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n551_), .B1(new_n458_), .B2(new_n546_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(KEYINPUT100), .A3(KEYINPUT33), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n528_), .A2(new_n530_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n524_), .A2(KEYINPUT32), .ZN(new_n556_));
  MUX2_X1   g355(.A(new_n555_), .B(new_n535_), .S(new_n556_), .Z(new_n557_));
  AOI22_X1  g356(.A1(new_n550_), .A2(new_n554_), .B1(new_n460_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n434_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n432_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  OAI21_X1  g360(.A(new_n541_), .B1(new_n558_), .B2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n500_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n563_), .A2(new_n498_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT86), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(KEYINPUT86), .B1(new_n563_), .B2(new_n498_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n540_), .B1(new_n562_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n294_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT80), .ZN(new_n572_));
  NOR3_X1   g371(.A1(new_n272_), .A2(new_n273_), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT80), .B1(new_n257_), .B2(new_n260_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n571_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n294_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G229gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT81), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n575_), .A2(new_n576_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n579_), .A2(KEYINPUT82), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n573_), .A2(new_n574_), .A3(new_n571_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n572_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n257_), .A2(KEYINPUT80), .A3(new_n260_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n294_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(G229gat), .B(G233gat), .C1(new_n581_), .C2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT82), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n575_), .A2(new_n576_), .A3(new_n586_), .A4(new_n578_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n580_), .A2(new_n585_), .A3(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G169gat), .B(G197gat), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n589_), .B(new_n590_), .Z(new_n591_));
  NOR2_X1   g390(.A1(new_n591_), .A2(KEYINPUT83), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n588_), .B(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OR3_X1    g393(.A1(new_n570_), .A2(KEYINPUT103), .A3(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(KEYINPUT103), .B1(new_n570_), .B2(new_n594_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n324_), .A2(KEYINPUT79), .A3(new_n358_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n461_), .A2(G1gat), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n361_), .A2(new_n597_), .A3(new_n598_), .A4(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT38), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n600_), .A2(new_n601_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n283_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(new_n570_), .A2(new_n604_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n357_), .A2(new_n322_), .A3(new_n594_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(G1gat), .B1(new_n607_), .B2(new_n461_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n602_), .A2(new_n603_), .A3(new_n608_), .ZN(G1324gat));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n610_));
  INV_X1    g409(.A(new_n607_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n539_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n610_), .B1(new_n613_), .B2(G8gat), .ZN(new_n614_));
  AOI211_X1 g413(.A(KEYINPUT39), .B(new_n290_), .C1(new_n611_), .C2(new_n612_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n361_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n612_), .A2(new_n290_), .ZN(new_n617_));
  OAI22_X1  g416(.A1(new_n614_), .A2(new_n615_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT40), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(G1325gat));
  OAI21_X1  g419(.A(G15gat), .B1(new_n607_), .B2(new_n569_), .ZN(new_n621_));
  XOR2_X1   g420(.A(new_n621_), .B(KEYINPUT41), .Z(new_n622_));
  NAND2_X1  g421(.A1(new_n568_), .A2(new_n487_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n622_), .B1(new_n616_), .B2(new_n623_), .ZN(G1326gat));
  OR2_X1    g423(.A1(new_n435_), .A2(G22gat), .ZN(new_n625_));
  OAI21_X1  g424(.A(G22gat), .B1(new_n607_), .B2(new_n435_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(KEYINPUT42), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n626_), .A2(KEYINPUT42), .ZN(new_n628_));
  OAI22_X1  g427(.A1(new_n616_), .A2(new_n625_), .B1(new_n627_), .B2(new_n628_), .ZN(G1327gat));
  INV_X1    g428(.A(new_n322_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n283_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n358_), .A2(new_n631_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n633_));
  AOI21_X1  g432(.A(G29gat), .B1(new_n633_), .B2(new_n460_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n287_), .ZN(new_n635_));
  OAI21_X1  g434(.A(KEYINPUT43), .B1(new_n570_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT43), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n550_), .A2(new_n554_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n557_), .A2(new_n460_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n435_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n568_), .B1(new_n641_), .B2(new_n541_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n637_), .B(new_n287_), .C1(new_n642_), .C2(new_n540_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n636_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n358_), .A2(new_n322_), .A3(new_n593_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n644_), .A2(KEYINPUT44), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(KEYINPUT44), .B1(new_n644_), .B2(new_n646_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n460_), .A2(G29gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n634_), .B1(new_n649_), .B2(new_n650_), .ZN(G1328gat));
  INV_X1    g450(.A(G36gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n633_), .A2(new_n652_), .A3(new_n612_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT45), .ZN(new_n654_));
  XNOR2_X1  g453(.A(KEYINPUT104), .B(KEYINPUT46), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n647_), .A2(new_n648_), .A3(new_n539_), .ZN(new_n656_));
  OAI211_X1 g455(.A(new_n654_), .B(new_n655_), .C1(new_n656_), .C2(new_n652_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n655_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT45), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n653_), .B(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n656_), .A2(new_n652_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n657_), .A2(new_n662_), .ZN(G1329gat));
  AOI21_X1  g462(.A(G43gat), .B1(new_n633_), .B2(new_n568_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n564_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(new_n482_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n664_), .B1(new_n649_), .B2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(G1330gat));
  NOR3_X1   g468(.A1(new_n647_), .A2(new_n648_), .A3(new_n435_), .ZN(new_n670_));
  INV_X1    g469(.A(G50gat), .ZN(new_n671_));
  INV_X1    g470(.A(new_n633_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n561_), .A2(new_n671_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT106), .ZN(new_n674_));
  OAI22_X1  g473(.A1(new_n670_), .A2(new_n671_), .B1(new_n672_), .B2(new_n674_), .ZN(G1331gat));
  OR3_X1    g474(.A1(new_n570_), .A2(KEYINPUT107), .A3(new_n593_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(new_n357_), .ZN(new_n677_));
  OAI21_X1  g476(.A(KEYINPUT107), .B1(new_n570_), .B2(new_n593_), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n324_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT108), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n679_), .A2(KEYINPUT108), .A3(new_n324_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n461_), .A2(G57gat), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n682_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n322_), .A2(new_n593_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n605_), .A2(new_n357_), .A3(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G57gat), .B1(new_n687_), .B2(new_n461_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n685_), .A2(new_n688_), .ZN(G1332gat));
  NOR2_X1   g488(.A1(new_n539_), .A2(G64gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n682_), .A2(new_n683_), .A3(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(G64gat), .B1(new_n687_), .B2(new_n539_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT48), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1333gat));
  NOR2_X1   g493(.A1(new_n569_), .A2(G71gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n682_), .A2(new_n683_), .A3(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G71gat), .B1(new_n687_), .B2(new_n569_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT49), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n696_), .A2(new_n698_), .ZN(G1334gat));
  NOR2_X1   g498(.A1(new_n435_), .A2(G78gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n682_), .A2(new_n683_), .A3(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(G78gat), .B1(new_n687_), .B2(new_n435_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT50), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(G1335gat));
  NAND3_X1  g503(.A1(new_n357_), .A2(new_n322_), .A3(new_n594_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n705_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n636_), .A2(new_n643_), .A3(KEYINPUT109), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT109), .B1(new_n636_), .B2(new_n643_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n706_), .B1(new_n707_), .B2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(G85gat), .B1(new_n709_), .B2(new_n461_), .ZN(new_n710_));
  AND4_X1   g509(.A1(new_n357_), .A2(new_n676_), .A3(new_n631_), .A4(new_n678_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n711_), .A2(new_n221_), .A3(new_n460_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1336gat));
  OAI21_X1  g512(.A(G92gat), .B1(new_n709_), .B2(new_n539_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(new_n222_), .A3(new_n612_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(G1337gat));
  OAI211_X1 g515(.A(new_n568_), .B(new_n706_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(G99gat), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(KEYINPUT110), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT110), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n717_), .A2(new_n720_), .A3(G99gat), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n665_), .A2(new_n245_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n711_), .B2(new_n723_), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n719_), .A2(new_n721_), .A3(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT51), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n719_), .A2(new_n727_), .A3(new_n721_), .A4(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n726_), .A2(new_n728_), .ZN(G1338gat));
  NAND3_X1  g528(.A1(new_n711_), .A2(new_n212_), .A3(new_n561_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT52), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n705_), .A2(new_n435_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n644_), .A2(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n733_), .B2(G106gat), .ZN(new_n734_));
  AOI211_X1 g533(.A(KEYINPUT52), .B(new_n212_), .C1(new_n644_), .C2(new_n732_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n730_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g536(.A1(new_n635_), .A2(new_n358_), .A3(new_n686_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT113), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n738_), .A2(new_n740_), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n739_), .A2(KEYINPUT113), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n635_), .A2(new_n358_), .A3(new_n686_), .A4(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n353_), .A2(new_n594_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT114), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n247_), .A2(new_n248_), .A3(new_n329_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n340_), .B1(KEYINPUT12), .B2(new_n332_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n748_), .B2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n331_), .A2(new_n335_), .A3(KEYINPUT114), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n750_), .A2(new_n338_), .A3(new_n751_), .ZN(new_n752_));
  AOI22_X1  g551(.A1(new_n249_), .A2(new_n330_), .B1(new_n334_), .B2(new_n333_), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n753_), .A2(KEYINPUT115), .A3(KEYINPUT55), .A4(new_n336_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT55), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n337_), .A2(new_n755_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n331_), .A2(new_n335_), .A3(KEYINPUT55), .A4(new_n336_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT115), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n752_), .A2(new_n754_), .A3(new_n756_), .A4(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n349_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT56), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n760_), .A2(KEYINPUT56), .A3(new_n349_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n746_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n766_));
  INV_X1    g565(.A(new_n578_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n582_), .A2(new_n294_), .A3(new_n583_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n575_), .B2(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n766_), .B1(new_n769_), .B2(new_n591_), .ZN(new_n770_));
  OAI21_X1  g569(.A(new_n578_), .B1(new_n581_), .B2(new_n584_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n591_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(KEYINPUT116), .A3(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n575_), .A2(new_n576_), .A3(new_n767_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n770_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n580_), .A2(new_n591_), .A3(new_n585_), .A4(new_n587_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT117), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(KEYINPUT117), .A3(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n350_), .B2(new_n353_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n283_), .B1(new_n765_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT58), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n760_), .A2(KEYINPUT56), .A3(new_n349_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT56), .B1(new_n760_), .B2(new_n349_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n781_), .A2(new_n352_), .A3(KEYINPUT118), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT118), .B1(new_n781_), .B2(new_n352_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n787_), .B1(new_n790_), .B2(new_n793_), .ZN(new_n794_));
  OR2_X1    g593(.A1(new_n791_), .A2(new_n792_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n795_), .B(KEYINPUT58), .C1(new_n789_), .C2(new_n788_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n794_), .A2(new_n287_), .A3(new_n796_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n745_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n604_), .B1(new_n798_), .B2(new_n782_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT57), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n786_), .A2(new_n797_), .A3(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT120), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n322_), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n802_), .B1(new_n801_), .B2(new_n322_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n744_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n561_), .A2(new_n612_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n665_), .A2(new_n461_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  XOR2_X1   g609(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n812_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n801_), .A2(new_n322_), .ZN(new_n814_));
  INV_X1    g613(.A(new_n744_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n810_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  AOI22_X1  g615(.A1(new_n806_), .A2(new_n813_), .B1(new_n816_), .B2(KEYINPUT59), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n593_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(G113gat), .ZN(new_n819_));
  OR3_X1    g618(.A1(new_n816_), .A2(G113gat), .A3(new_n594_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(G1340gat));
  NAND2_X1  g620(.A1(new_n817_), .A2(new_n357_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(G120gat), .ZN(new_n823_));
  INV_X1    g622(.A(new_n816_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT60), .ZN(new_n825_));
  AOI21_X1  g624(.A(G120gat), .B1(new_n357_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n825_), .B2(G120gat), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n824_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT121), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT121), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n824_), .A2(new_n830_), .A3(new_n827_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n823_), .A2(new_n832_), .ZN(G1341gat));
  AOI21_X1  g632(.A(G127gat), .B1(new_n824_), .B2(new_n630_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n322_), .A2(KEYINPUT122), .ZN(new_n835_));
  MUX2_X1   g634(.A(KEYINPUT122), .B(new_n835_), .S(G127gat), .Z(new_n836_));
  AOI21_X1  g635(.A(new_n834_), .B1(new_n817_), .B2(new_n836_), .ZN(G1342gat));
  NAND2_X1  g636(.A1(new_n817_), .A2(new_n287_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G134gat), .ZN(new_n839_));
  OR3_X1    g638(.A1(new_n816_), .A2(G134gat), .A3(new_n283_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(G1343gat));
  NOR2_X1   g640(.A1(new_n814_), .A2(new_n815_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n568_), .ZN(new_n843_));
  NOR3_X1   g642(.A1(new_n435_), .A2(new_n612_), .A3(new_n461_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT123), .B(G141gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n593_), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n847_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n849_), .B1(new_n845_), .B2(new_n594_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(G1344gat));
  NAND3_X1  g650(.A1(new_n846_), .A2(new_n370_), .A3(new_n357_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G148gat), .B1(new_n845_), .B2(new_n358_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1345gat));
  XNOR2_X1  g653(.A(KEYINPUT61), .B(G155gat), .ZN(new_n855_));
  OR3_X1    g654(.A1(new_n845_), .A2(new_n322_), .A3(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n845_), .B2(new_n322_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1346gat));
  OR3_X1    g657(.A1(new_n845_), .A2(G162gat), .A3(new_n283_), .ZN(new_n859_));
  OAI21_X1  g658(.A(G162gat), .B1(new_n845_), .B2(new_n635_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1347gat));
  NOR2_X1   g660(.A1(new_n539_), .A2(new_n460_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  NOR3_X1   g662(.A1(new_n569_), .A2(new_n561_), .A3(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n806_), .A2(new_n593_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(G169gat), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n864_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n793_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n287_), .B1(new_n870_), .B2(KEYINPUT58), .ZN(new_n871_));
  INV_X1    g670(.A(new_n796_), .ZN(new_n872_));
  OAI22_X1  g671(.A1(new_n871_), .A2(new_n872_), .B1(new_n799_), .B2(KEYINPUT57), .ZN(new_n873_));
  NOR2_X1   g672(.A1(new_n784_), .A2(new_n785_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n322_), .B1(new_n873_), .B2(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT120), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(new_n803_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n869_), .B1(new_n877_), .B2(new_n744_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n467_), .A3(new_n593_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n865_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n868_), .A2(new_n879_), .A3(new_n880_), .ZN(G1348gat));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882_));
  AOI21_X1  g681(.A(G176gat), .B1(new_n878_), .B2(new_n357_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n842_), .A2(new_n869_), .ZN(new_n884_));
  INV_X1    g683(.A(G176gat), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n358_), .A2(new_n885_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n884_), .A2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n882_), .B1(new_n883_), .B2(new_n887_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n806_), .A2(new_n357_), .A3(new_n864_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n885_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n884_), .A2(new_n886_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n890_), .A2(KEYINPUT124), .A3(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n888_), .A2(new_n892_), .ZN(G1349gat));
  AOI21_X1  g692(.A(G183gat), .B1(new_n884_), .B2(new_n630_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n322_), .A2(new_n504_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n894_), .B1(new_n878_), .B2(new_n895_), .ZN(G1350gat));
  NAND2_X1  g695(.A1(new_n878_), .A2(new_n287_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(G190gat), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n878_), .A2(new_n604_), .A3(new_n476_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1351gat));
  XOR2_X1   g699(.A(KEYINPUT125), .B(G197gat), .Z(new_n901_));
  NOR2_X1   g700(.A1(new_n863_), .A2(new_n435_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n843_), .A2(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n901_), .B1(new_n903_), .B2(new_n594_), .ZN(new_n904_));
  INV_X1    g703(.A(G197gat), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT125), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n843_), .A2(new_n593_), .A3(new_n902_), .A4(new_n906_), .ZN(new_n907_));
  AND2_X1   g706(.A1(new_n904_), .A2(new_n907_), .ZN(G1352gat));
  OR3_X1    g707(.A1(new_n903_), .A2(G204gat), .A3(new_n358_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G204gat), .B1(new_n903_), .B2(new_n358_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1353gat));
  INV_X1    g710(.A(new_n903_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(KEYINPUT126), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n322_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n912_), .A2(new_n914_), .A3(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n914_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n915_), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n903_), .B2(new_n918_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n916_), .A2(new_n919_), .ZN(G1354gat));
  NAND2_X1  g719(.A1(new_n912_), .A2(new_n604_), .ZN(new_n921_));
  INV_X1    g720(.A(G218gat), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n287_), .A2(G218gat), .ZN(new_n923_));
  XOR2_X1   g722(.A(new_n923_), .B(KEYINPUT127), .Z(new_n924_));
  AOI22_X1  g723(.A1(new_n921_), .A2(new_n922_), .B1(new_n912_), .B2(new_n924_), .ZN(G1355gat));
endmodule


