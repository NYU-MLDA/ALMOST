//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n865_, new_n867_, new_n868_, new_n870_, new_n871_, new_n872_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n901_, new_n902_, new_n904_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  INV_X1    g001(.A(G113gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G120gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(G141gat), .ZN(new_n208_));
  INV_X1    g007(.A(G148gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G155gat), .A2(G162gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT1), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT82), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(KEYINPUT1), .B2(new_n211_), .ZN(new_n216_));
  OAI211_X1 g015(.A(new_n207_), .B(new_n210_), .C1(new_n213_), .C2(new_n216_), .ZN(new_n217_));
  AND2_X1   g016(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n218_));
  NOR2_X1   g017(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n210_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  OAI21_X1  g019(.A(new_n220_), .B1(new_n210_), .B2(new_n218_), .ZN(new_n221_));
  XOR2_X1   g020(.A(new_n207_), .B(KEYINPUT2), .Z(new_n222_));
  OAI211_X1 g021(.A(new_n211_), .B(new_n215_), .C1(new_n221_), .C2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n206_), .A2(new_n217_), .A3(new_n223_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n204_), .B(G120gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n217_), .A2(new_n223_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(KEYINPUT4), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT90), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n229_), .B1(new_n227_), .B2(KEYINPUT4), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G225gat), .A2(G233gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT4), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n225_), .A2(new_n226_), .A3(KEYINPUT90), .A4(new_n233_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n228_), .A2(new_n230_), .A3(new_n232_), .A4(new_n234_), .ZN(new_n235_));
  AND2_X1   g034(.A1(new_n224_), .A2(new_n227_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT91), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n231_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n224_), .A2(new_n227_), .ZN(new_n239_));
  OAI21_X1  g038(.A(KEYINPUT91), .B1(new_n239_), .B2(new_n232_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n235_), .A2(new_n238_), .A3(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G57gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(G85gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(G1gat), .B(G29gat), .Z(new_n244_));
  XOR2_X1   g043(.A(new_n243_), .B(new_n244_), .Z(new_n245_));
  NAND2_X1  g044(.A1(new_n241_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT93), .ZN(new_n247_));
  INV_X1    g046(.A(new_n245_), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n235_), .A2(new_n238_), .A3(new_n240_), .A4(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n246_), .A2(new_n247_), .A3(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n241_), .A2(KEYINPUT93), .A3(new_n245_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT84), .B(G197gat), .ZN(new_n252_));
  INV_X1    g051(.A(G204gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G197gat), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n254_), .B(KEYINPUT21), .C1(new_n255_), .C2(new_n253_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G211gat), .B(G218gat), .Z(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(G204gat), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n259_), .B1(new_n255_), .B2(G204gat), .ZN(new_n260_));
  OAI211_X1 g059(.A(new_n256_), .B(new_n258_), .C1(new_n260_), .C2(KEYINPUT21), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(KEYINPUT21), .A3(new_n257_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT85), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT22), .B(G169gat), .ZN(new_n266_));
  INV_X1    g065(.A(G176gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT79), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n269_), .B(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT23), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n273_), .B1(G183gat), .B2(G190gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n273_), .A2(G183gat), .A3(G190gat), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n275_), .A2(KEYINPUT81), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(KEYINPUT81), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n274_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NOR2_X1   g077(.A1(G183gat), .A2(G190gat), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n272_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(new_n275_), .A2(KEYINPUT80), .ZN(new_n281_));
  INV_X1    g080(.A(new_n274_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n275_), .A2(KEYINPUT80), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n281_), .A2(new_n282_), .A3(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(G169gat), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(new_n267_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n271_), .A2(KEYINPUT24), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(G183gat), .ZN(new_n288_));
  OR3_X1    g087(.A1(new_n288_), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G190gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT25), .B1(new_n288_), .B2(KEYINPUT78), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n289_), .A2(new_n290_), .A3(new_n291_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n286_), .A2(KEYINPUT24), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n284_), .A2(new_n287_), .A3(new_n292_), .A4(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n280_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n261_), .A2(KEYINPUT85), .A3(new_n262_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n265_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(KEYINPUT25), .B(G183gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT88), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n290_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n278_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n286_), .A2(KEYINPUT24), .A3(new_n269_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n301_), .A2(new_n302_), .A3(new_n293_), .A4(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n284_), .B1(G183gat), .B2(G190gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(new_n272_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n304_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n263_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n298_), .A2(KEYINPUT20), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G226gat), .A2(G233gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT19), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT18), .B(G64gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(G92gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G8gat), .B(G36gat), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n315_), .B(new_n316_), .Z(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT32), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT20), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n265_), .A2(new_n297_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n320_), .B1(new_n321_), .B2(new_n295_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n307_), .A2(new_n263_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n313_), .B(new_n319_), .C1(new_n324_), .C2(new_n312_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n309_), .A2(new_n311_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT89), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n322_), .A2(new_n312_), .A3(new_n323_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT89), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n309_), .A2(new_n329_), .A3(new_n311_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n327_), .A2(new_n328_), .A3(new_n318_), .A4(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n250_), .A2(new_n251_), .A3(new_n325_), .A4(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n327_), .A2(new_n328_), .A3(new_n330_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n317_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND4_X1  g134(.A1(new_n327_), .A2(new_n328_), .A3(new_n317_), .A4(new_n330_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n236_), .A2(new_n232_), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n228_), .A2(new_n230_), .A3(new_n234_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n245_), .B(new_n337_), .C1(new_n338_), .C2(new_n232_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n335_), .A2(new_n336_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT92), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n249_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT33), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT33), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n249_), .A2(new_n341_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  OAI21_X1  g145(.A(new_n332_), .B1(new_n340_), .B2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G15gat), .B(G43gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n348_), .B(KEYINPUT31), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n295_), .A2(KEYINPUT30), .ZN(new_n350_));
  INV_X1    g149(.A(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n295_), .A2(KEYINPUT30), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n351_), .A2(new_n225_), .A3(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n295_), .A2(KEYINPUT30), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n206_), .B1(new_n354_), .B2(new_n350_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n349_), .B1(new_n353_), .B2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n225_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n354_), .A2(new_n206_), .A3(new_n350_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n349_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n356_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G71gat), .B(G99gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G227gat), .A2(G233gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n361_), .A2(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n356_), .A2(new_n364_), .A3(new_n360_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NOR2_X1   g168(.A1(new_n226_), .A2(KEYINPUT29), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G22gat), .B(G50gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT28), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n370_), .B(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n226_), .A2(KEYINPUT29), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(new_n263_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n375_), .A2(G228gat), .A3(G233gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G228gat), .A2(G233gat), .ZN(new_n377_));
  AND3_X1   g176(.A1(new_n261_), .A2(KEYINPUT85), .A3(new_n262_), .ZN(new_n378_));
  AOI21_X1  g177(.A(KEYINPUT85), .B1(new_n261_), .B2(new_n262_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n377_), .B(new_n374_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(G78gat), .B(G106gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n381_), .B(KEYINPUT86), .ZN(new_n382_));
  AND3_X1   g181(.A1(new_n376_), .A2(new_n380_), .A3(new_n382_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n382_), .B1(new_n376_), .B2(new_n380_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n373_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT87), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT87), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n387_), .B(new_n373_), .C1(new_n383_), .C2(new_n384_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n376_), .A2(new_n380_), .ZN(new_n390_));
  AND2_X1   g189(.A1(new_n390_), .A2(new_n381_), .ZN(new_n391_));
  OR3_X1    g190(.A1(new_n391_), .A2(new_n383_), .A3(new_n373_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n369_), .A2(new_n389_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n347_), .A2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n250_), .A2(new_n251_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n389_), .A2(new_n368_), .A3(new_n392_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n368_), .B1(new_n389_), .B2(new_n392_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n396_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n335_), .A2(new_n336_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT27), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OAI211_X1 g201(.A(new_n334_), .B(new_n313_), .C1(new_n324_), .C2(new_n312_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n336_), .A2(KEYINPUT27), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n395_), .B1(new_n399_), .B2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT16), .B(G183gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(G211gat), .ZN(new_n408_));
  XOR2_X1   g207(.A(G127gat), .B(G155gat), .Z(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G57gat), .B(G64gat), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n411_), .A2(KEYINPUT11), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(KEYINPUT11), .ZN(new_n413_));
  XOR2_X1   g212(.A(G71gat), .B(G78gat), .Z(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  OR2_X1    g214(.A1(new_n413_), .A2(new_n414_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G231gat), .A2(G233gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(G1gat), .B(G8gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G1gat), .A2(G8gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(KEYINPUT14), .ZN(new_n422_));
  INV_X1    g221(.A(G15gat), .ZN(new_n423_));
  INV_X1    g222(.A(G22gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NOR2_X1   g224(.A1(G15gat), .A2(G22gat), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n422_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(KEYINPUT74), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n427_), .A2(KEYINPUT74), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n420_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n430_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n420_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(new_n433_), .A3(new_n428_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n431_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n419_), .B(new_n436_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n410_), .B1(new_n437_), .B2(KEYINPUT17), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(KEYINPUT17), .B2(new_n410_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n437_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(KEYINPUT75), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n439_), .B(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT9), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT65), .B(G85gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT66), .B(G92gat), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n443_), .B1(new_n444_), .B2(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(G85gat), .A2(G92gat), .ZN(new_n447_));
  NAND3_X1  g246(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT67), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n446_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G99gat), .A2(G106gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT6), .ZN(new_n452_));
  INV_X1    g251(.A(G106gat), .ZN(new_n453_));
  INV_X1    g252(.A(G99gat), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT10), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT10), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(G99gat), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT64), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n455_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n453_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n450_), .A2(new_n452_), .A3(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(G29gat), .ZN(new_n463_));
  INV_X1    g262(.A(G36gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G43gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G29gat), .A2(G36gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G50gat), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n466_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n469_), .A2(new_n470_), .A3(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G29gat), .B(G36gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(G43gat), .ZN(new_n474_));
  AOI21_X1  g273(.A(G50gat), .B1(new_n474_), .B2(new_n468_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n472_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NOR3_X1   g278(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n482_));
  NOR2_X1   g281(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n451_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT69), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AND2_X1   g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(KEYINPUT69), .A2(KEYINPUT6), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n481_), .A2(new_n484_), .A3(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G85gat), .B(G92gat), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n477_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n481_), .A2(new_n452_), .ZN(new_n495_));
  XNOR2_X1  g294(.A(KEYINPUT68), .B(KEYINPUT8), .ZN(new_n496_));
  AND3_X1   g295(.A1(new_n495_), .A2(new_n493_), .A3(new_n496_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n462_), .B(new_n476_), .C1(new_n494_), .C2(new_n497_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n450_), .A2(new_n452_), .A3(new_n461_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n484_), .A2(new_n490_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n480_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n478_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n493_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n492_), .B1(new_n481_), .B2(new_n452_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n503_), .A2(KEYINPUT8), .B1(new_n504_), .B2(new_n496_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n499_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT15), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n472_), .A2(new_n475_), .A3(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n470_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n474_), .A2(G50gat), .A3(new_n468_), .ZN(new_n510_));
  AOI21_X1  g309(.A(KEYINPUT15), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n498_), .B1(new_n506_), .B2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(G232gat), .A2(G233gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT34), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n513_), .A2(KEYINPUT35), .A3(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(KEYINPUT71), .B(G134gat), .ZN(new_n517_));
  INV_X1    g316(.A(G162gat), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n517_), .B(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G190gat), .B(G218gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n519_), .B(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT36), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n507_), .B1(new_n472_), .B2(new_n475_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n509_), .A2(KEYINPUT15), .A3(new_n510_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n526_), .B1(new_n505_), .B2(new_n499_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n515_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT35), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n515_), .A2(KEYINPUT35), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND4_X1  g332(.A1(new_n527_), .A2(new_n531_), .A3(new_n533_), .A4(new_n498_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n516_), .A2(new_n523_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT72), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n516_), .A2(KEYINPUT72), .A3(new_n523_), .A4(new_n534_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n521_), .B(KEYINPUT36), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n516_), .B2(new_n534_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT37), .ZN(new_n544_));
  OR2_X1    g343(.A1(new_n544_), .A2(KEYINPUT73), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(KEYINPUT73), .ZN(new_n546_));
  AND4_X1   g345(.A1(new_n539_), .A2(new_n543_), .A3(new_n545_), .A4(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n542_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n546_), .B1(new_n548_), .B2(new_n545_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n547_), .A2(new_n549_), .ZN(new_n550_));
  AND3_X1   g349(.A1(new_n406_), .A2(new_n442_), .A3(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT13), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G120gat), .B(G148gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(new_n253_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT5), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(new_n267_), .ZN(new_n556_));
  INV_X1    g355(.A(new_n417_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n557_), .B1(new_n499_), .B2(new_n505_), .ZN(new_n558_));
  OAI211_X1 g357(.A(new_n462_), .B(new_n417_), .C1(new_n494_), .C2(new_n497_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n558_), .A2(KEYINPUT12), .A3(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT12), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n561_), .B(new_n557_), .C1(new_n499_), .C2(new_n505_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(G230gat), .A2(G233gat), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT70), .ZN(new_n566_));
  INV_X1    g365(.A(new_n564_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n567_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT70), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n566_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n558_), .A2(new_n559_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n567_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n556_), .B1(new_n571_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n569_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n576_));
  AOI211_X1 g375(.A(KEYINPUT70), .B(new_n567_), .C1(new_n560_), .C2(new_n562_), .ZN(new_n577_));
  OAI211_X1 g376(.A(new_n573_), .B(new_n556_), .C1(new_n576_), .C2(new_n577_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n552_), .B1(new_n575_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n578_), .ZN(new_n580_));
  NOR3_X1   g379(.A1(new_n574_), .A2(new_n580_), .A3(KEYINPUT13), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G229gat), .A2(G233gat), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n431_), .A2(new_n434_), .A3(new_n476_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n476_), .B1(new_n431_), .B2(new_n434_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n585_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n526_), .A2(new_n435_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n590_), .A2(new_n584_), .A3(new_n586_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G113gat), .B(G141gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(new_n285_), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(new_n255_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n589_), .A2(new_n591_), .A3(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT77), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n589_), .A2(new_n591_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT76), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT76), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n589_), .A2(new_n591_), .A3(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n599_), .A2(new_n594_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n597_), .A2(new_n602_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n551_), .A2(new_n583_), .A3(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(G1gat), .ZN(new_n605_));
  INV_X1    g404(.A(new_n396_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT38), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n548_), .B(KEYINPUT95), .Z(new_n609_));
  NAND2_X1  g408(.A1(new_n406_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT96), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n603_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n442_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n582_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n615_), .B(KEYINPUT94), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n612_), .A2(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n617_), .B2(new_n396_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n608_), .A2(new_n618_), .ZN(G1324gat));
  XOR2_X1   g418(.A(KEYINPUT98), .B(KEYINPUT40), .Z(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n612_), .A2(new_n405_), .A3(new_n616_), .ZN(new_n623_));
  XOR2_X1   g422(.A(KEYINPUT97), .B(KEYINPUT39), .Z(new_n624_));
  AND3_X1   g423(.A1(new_n623_), .A2(G8gat), .A3(new_n624_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n624_), .B1(new_n623_), .B2(G8gat), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(G8gat), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n604_), .A2(new_n628_), .A3(new_n405_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n622_), .B1(new_n627_), .B2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n623_), .A2(G8gat), .ZN(new_n631_));
  INV_X1    g430(.A(new_n624_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n623_), .A2(G8gat), .A3(new_n624_), .ZN(new_n634_));
  AND4_X1   g433(.A1(new_n622_), .A2(new_n633_), .A3(new_n629_), .A4(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n621_), .B1(new_n630_), .B2(new_n635_), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n627_), .A2(new_n622_), .A3(new_n629_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n633_), .A2(new_n629_), .A3(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT99), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n637_), .A2(new_n639_), .A3(new_n620_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(G1325gat));
  OAI21_X1  g440(.A(G15gat), .B1(new_n617_), .B2(new_n369_), .ZN(new_n642_));
  XOR2_X1   g441(.A(new_n642_), .B(KEYINPUT41), .Z(new_n643_));
  NAND3_X1  g442(.A1(new_n604_), .A2(new_n423_), .A3(new_n368_), .ZN(new_n644_));
  XOR2_X1   g443(.A(new_n644_), .B(KEYINPUT100), .Z(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(G1326gat));
  NAND2_X1  g445(.A1(new_n389_), .A2(new_n392_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n604_), .A2(new_n424_), .A3(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n612_), .A2(new_n647_), .A3(new_n616_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n649_), .A2(G22gat), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT101), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(KEYINPUT101), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n651_), .A2(KEYINPUT42), .A3(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(KEYINPUT42), .B1(new_n651_), .B2(new_n652_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n648_), .B1(new_n653_), .B2(new_n654_), .ZN(G1327gat));
  AND2_X1   g454(.A1(new_n406_), .A2(new_n548_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n582_), .A2(new_n613_), .A3(new_n442_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(new_n463_), .A3(new_n606_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  INV_X1    g460(.A(new_n550_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n406_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT103), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n406_), .A2(new_n665_), .A3(new_n661_), .A4(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n550_), .B1(new_n406_), .B2(KEYINPUT102), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT102), .ZN(new_n669_));
  OAI211_X1 g468(.A(new_n395_), .B(new_n669_), .C1(new_n399_), .C2(new_n405_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n661_), .B1(new_n668_), .B2(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n657_), .B1(new_n667_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT104), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n672_), .A2(new_n673_), .A3(KEYINPUT44), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT44), .B1(new_n672_), .B2(new_n673_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n396_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n660_), .B1(new_n678_), .B2(new_n463_), .ZN(G1328gat));
  INV_X1    g478(.A(KEYINPUT46), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(KEYINPUT106), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT107), .Z(new_n682_));
  OAI21_X1  g481(.A(new_n405_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G36gat), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n405_), .A2(KEYINPUT105), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n405_), .A2(KEYINPUT105), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n659_), .A2(new_n464_), .A3(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT45), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n688_), .B(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n682_), .B1(new_n684_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n682_), .ZN(new_n693_));
  AOI211_X1 g492(.A(new_n693_), .B(new_n690_), .C1(new_n683_), .C2(G36gat), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1329gat));
  INV_X1    g494(.A(KEYINPUT47), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n368_), .B1(new_n674_), .B2(new_n676_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G43gat), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n658_), .A2(G43gat), .A3(new_n369_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n696_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n701_));
  AOI211_X1 g500(.A(KEYINPUT47), .B(new_n699_), .C1(new_n697_), .C2(G43gat), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1330gat));
  NAND3_X1  g502(.A1(new_n659_), .A2(new_n470_), .A3(new_n647_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n647_), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n705_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n704_), .B1(new_n706_), .B2(new_n470_), .ZN(G1331gat));
  NOR2_X1   g506(.A1(new_n583_), .A2(new_n603_), .ZN(new_n708_));
  AND2_X1   g507(.A1(new_n551_), .A2(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(G57gat), .B1(new_n709_), .B2(new_n606_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n612_), .A2(new_n442_), .A3(new_n708_), .ZN(new_n711_));
  INV_X1    g510(.A(G57gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n606_), .B2(KEYINPUT108), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(KEYINPUT108), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n710_), .B1(new_n714_), .B2(new_n715_), .ZN(G1332gat));
  INV_X1    g515(.A(new_n711_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n687_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n718_), .A2(G64gat), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT109), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n718_), .A2(new_n721_), .A3(G64gat), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n720_), .A2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT48), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(G64gat), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n709_), .A2(new_n726_), .A3(new_n687_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n720_), .A2(KEYINPUT48), .A3(new_n722_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n725_), .A2(new_n727_), .A3(new_n728_), .ZN(G1333gat));
  OAI21_X1  g528(.A(G71gat), .B1(new_n711_), .B2(new_n369_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT49), .ZN(new_n731_));
  INV_X1    g530(.A(G71gat), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n709_), .A2(new_n732_), .A3(new_n368_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n731_), .A2(new_n733_), .ZN(G1334gat));
  INV_X1    g533(.A(G78gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n709_), .A2(new_n735_), .A3(new_n647_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT50), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n717_), .A2(new_n647_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n738_), .B2(G78gat), .ZN(new_n739_));
  AOI211_X1 g538(.A(KEYINPUT50), .B(new_n735_), .C1(new_n717_), .C2(new_n647_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT110), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(new_n743_));
  OAI211_X1 g542(.A(KEYINPUT110), .B(new_n736_), .C1(new_n739_), .C2(new_n740_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1335gat));
  NOR3_X1   g544(.A1(new_n583_), .A2(new_n603_), .A3(new_n442_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n656_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  AOI21_X1  g547(.A(G85gat), .B1(new_n748_), .B2(new_n606_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n746_), .B1(new_n667_), .B2(new_n671_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT111), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  OAI211_X1 g551(.A(KEYINPUT111), .B(new_n746_), .C1(new_n667_), .C2(new_n671_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n396_), .A2(new_n444_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n749_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n756_), .B(new_n757_), .ZN(G1336gat));
  AOI21_X1  g557(.A(G92gat), .B1(new_n748_), .B2(new_n405_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n687_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n760_), .A2(new_n445_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT113), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n759_), .B1(new_n754_), .B2(new_n762_), .ZN(G1337gat));
  NAND3_X1  g562(.A1(new_n752_), .A2(new_n368_), .A3(new_n753_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(G99gat), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n748_), .B(new_n368_), .C1(new_n460_), .C2(new_n459_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  XOR2_X1   g566(.A(KEYINPUT114), .B(KEYINPUT51), .Z(new_n768_));
  XNOR2_X1  g567(.A(new_n767_), .B(new_n768_), .ZN(G1338gat));
  XNOR2_X1  g568(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n748_), .A2(new_n453_), .A3(new_n647_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n647_), .B(new_n746_), .C1(new_n667_), .C2(new_n671_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(G106gat), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n773_), .A2(KEYINPUT52), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(KEYINPUT52), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n770_), .B(new_n771_), .C1(new_n774_), .C2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n773_), .B(KEYINPUT52), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n770_), .B1(new_n778_), .B2(new_n771_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n777_), .A2(new_n779_), .ZN(G1339gat));
  OAI21_X1  g579(.A(new_n584_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n590_), .A2(new_n585_), .A3(new_n586_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n781_), .A2(new_n782_), .A3(new_n594_), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n578_), .A2(new_n597_), .A3(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n785_), .B1(new_n576_), .B2(new_n577_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n560_), .A2(new_n567_), .A3(new_n562_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(KEYINPUT55), .B2(new_n568_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n556_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT56), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT56), .ZN(new_n792_));
  AOI211_X1 g591(.A(new_n792_), .B(new_n556_), .C1(new_n786_), .C2(new_n788_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n784_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n550_), .B1(new_n794_), .B2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT55), .B1(new_n566_), .B2(new_n570_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n568_), .A2(KEYINPUT55), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n798_), .B1(new_n564_), .B2(new_n563_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n790_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n792_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n789_), .A2(KEYINPUT56), .A3(new_n790_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n803_), .A2(KEYINPUT116), .A3(KEYINPUT58), .A4(new_n784_), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT58), .B(new_n784_), .C1(new_n791_), .C2(new_n793_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n796_), .A2(new_n804_), .A3(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT57), .ZN(new_n809_));
  AND2_X1   g608(.A1(new_n603_), .A2(new_n578_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n810_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n811_));
  OAI211_X1 g610(.A(new_n597_), .B(new_n783_), .C1(new_n574_), .C2(new_n580_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n548_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n809_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  AOI211_X1 g614(.A(KEYINPUT57), .B(new_n548_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n808_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(new_n808_), .B(KEYINPUT117), .C1(new_n815_), .C2(new_n816_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n614_), .A3(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n550_), .A2(new_n613_), .A3(new_n442_), .ZN(new_n822_));
  OR3_X1    g621(.A1(new_n822_), .A2(new_n582_), .A3(KEYINPUT54), .ZN(new_n823_));
  OAI21_X1  g622(.A(KEYINPUT54), .B1(new_n822_), .B2(new_n582_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n821_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n821_), .A2(KEYINPUT118), .A3(new_n825_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n397_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n405_), .A2(new_n830_), .A3(new_n396_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n828_), .A2(new_n829_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT119), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n828_), .A2(new_n834_), .A3(new_n829_), .A4(new_n831_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(G113gat), .B1(new_n836_), .B2(new_n603_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n832_), .A2(KEYINPUT59), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n817_), .A2(new_n614_), .B1(new_n824_), .B2(new_n823_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n831_), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n841_));
  NOR3_X1   g640(.A1(new_n839_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  AND4_X1   g642(.A1(G113gat), .A2(new_n838_), .A3(new_n603_), .A4(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n837_), .A2(new_n844_), .ZN(G1340gat));
  OAI21_X1  g644(.A(new_n205_), .B1(new_n583_), .B2(KEYINPUT60), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n836_), .B(new_n846_), .C1(KEYINPUT60), .C2(new_n205_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n842_), .B1(new_n832_), .B2(KEYINPUT59), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n582_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n849_), .A2(G120gat), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n847_), .A2(new_n850_), .ZN(G1341gat));
  NAND2_X1  g650(.A1(new_n836_), .A2(new_n442_), .ZN(new_n852_));
  INV_X1    g651(.A(G127gat), .ZN(new_n853_));
  AOI211_X1 g652(.A(new_n853_), .B(new_n842_), .C1(new_n832_), .C2(KEYINPUT59), .ZN(new_n854_));
  AOI22_X1  g653(.A1(new_n852_), .A2(new_n853_), .B1(new_n442_), .B2(new_n854_), .ZN(G1342gat));
  INV_X1    g654(.A(new_n609_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n836_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(G134gat), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n550_), .A2(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT121), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n857_), .A2(new_n858_), .B1(new_n848_), .B2(new_n860_), .ZN(G1343gat));
  NAND4_X1  g660(.A1(new_n828_), .A2(new_n606_), .A3(new_n398_), .A4(new_n829_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n862_), .A2(new_n613_), .A3(new_n687_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(new_n208_), .ZN(G1344gat));
  NOR3_X1   g663(.A1(new_n862_), .A2(new_n583_), .A3(new_n687_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(new_n209_), .ZN(G1345gat));
  NOR3_X1   g665(.A1(new_n862_), .A2(new_n614_), .A3(new_n687_), .ZN(new_n867_));
  XOR2_X1   g666(.A(KEYINPUT61), .B(G155gat), .Z(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(G1346gat));
  NOR4_X1   g668(.A1(new_n862_), .A2(new_n518_), .A3(new_n550_), .A4(new_n687_), .ZN(new_n870_));
  AND3_X1   g669(.A1(new_n828_), .A2(new_n398_), .A3(new_n829_), .ZN(new_n871_));
  NAND4_X1  g670(.A1(new_n871_), .A2(new_n606_), .A3(new_n856_), .A4(new_n760_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n518_), .B2(new_n872_), .ZN(G1347gat));
  NAND2_X1  g672(.A1(new_n687_), .A2(new_n396_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(new_n397_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n839_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n877_), .A2(new_n603_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(G169gat), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT122), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n881_), .A3(G169gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n880_), .A2(KEYINPUT62), .A3(new_n882_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n266_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n885_), .B(new_n886_), .C1(new_n887_), .C2(new_n878_), .ZN(G1348gat));
  AND3_X1   g687(.A1(new_n821_), .A2(KEYINPUT118), .A3(new_n825_), .ZN(new_n889_));
  AOI21_X1  g688(.A(KEYINPUT118), .B1(new_n821_), .B2(new_n825_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n889_), .A2(new_n890_), .A3(new_n876_), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n891_), .A2(G176gat), .A3(new_n582_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT123), .ZN(new_n893_));
  INV_X1    g692(.A(new_n877_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n267_), .B1(new_n894_), .B2(new_n583_), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT123), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n891_), .A2(new_n896_), .A3(G176gat), .A4(new_n582_), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n893_), .A2(new_n895_), .A3(new_n897_), .ZN(G1349gat));
  NOR3_X1   g697(.A1(new_n894_), .A2(new_n300_), .A3(new_n614_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n876_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n828_), .A2(new_n442_), .A3(new_n829_), .A4(new_n900_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT124), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n899_), .B1(new_n902_), .B2(new_n288_), .ZN(G1350gat));
  OAI21_X1  g702(.A(G190gat), .B1(new_n894_), .B2(new_n550_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n856_), .A2(new_n290_), .ZN(new_n905_));
  XOR2_X1   g704(.A(new_n905_), .B(KEYINPUT125), .Z(new_n906_));
  OAI21_X1  g705(.A(new_n904_), .B1(new_n894_), .B2(new_n906_), .ZN(G1351gat));
  NAND2_X1  g706(.A1(new_n871_), .A2(new_n875_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(new_n255_), .A3(new_n603_), .ZN(new_n910_));
  OAI21_X1  g709(.A(G197gat), .B1(new_n908_), .B2(new_n613_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1352gat));
  NOR2_X1   g711(.A1(new_n253_), .A2(KEYINPUT126), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n909_), .A2(new_n582_), .A3(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n913_), .B1(new_n908_), .B2(new_n583_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1353gat));
  XNOR2_X1  g716(.A(KEYINPUT63), .B(G211gat), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n871_), .A2(new_n442_), .A3(new_n875_), .A4(new_n918_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n908_), .A2(new_n614_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n919_), .B1(new_n920_), .B2(new_n921_), .ZN(G1354gat));
  INV_X1    g721(.A(G218gat), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n550_), .A2(new_n923_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(KEYINPUT127), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n871_), .A2(new_n856_), .A3(new_n875_), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n909_), .A2(new_n925_), .B1(new_n926_), .B2(new_n923_), .ZN(G1355gat));
endmodule


