//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n867_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n887_, new_n888_, new_n890_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_;
  XNOR2_X1  g000(.A(G29gat), .B(G36gat), .ZN(new_n202_));
  INV_X1    g001(.A(G43gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G50gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT71), .B(KEYINPUT72), .Z(new_n208_));
  XNOR2_X1  g007(.A(G1gat), .B(G8gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G15gat), .ZN(new_n211_));
  INV_X1    g010(.A(G22gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G15gat), .A2(G22gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G1gat), .A2(G8gat), .ZN(new_n215_));
  AOI22_X1  g014(.A1(new_n213_), .A2(new_n214_), .B1(KEYINPUT14), .B2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n210_), .B(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n207_), .A2(new_n217_), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n206_), .B(KEYINPUT15), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n218_), .B1(new_n219_), .B2(new_n217_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G229gat), .A2(G233gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n207_), .B(new_n217_), .ZN(new_n223_));
  INV_X1    g022(.A(new_n221_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G113gat), .B(G141gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT76), .ZN(new_n227_));
  INV_X1    g026(.A(G169gat), .ZN(new_n228_));
  XNOR2_X1  g027(.A(new_n227_), .B(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G197gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n222_), .A2(new_n225_), .A3(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT77), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n222_), .A2(new_n225_), .ZN(new_n233_));
  INV_X1    g032(.A(new_n230_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT100), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT99), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G8gat), .B(G36gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT18), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(G64gat), .ZN(new_n242_));
  AND2_X1   g041(.A1(new_n242_), .A2(G92gat), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n242_), .A2(G92gat), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(G197gat), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n246_), .A2(G204gat), .ZN(new_n247_));
  INV_X1    g046(.A(G204gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n248_), .A2(G197gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT21), .B1(new_n247_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(G197gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n246_), .A2(G204gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT21), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G211gat), .B(G218gat), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n250_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G211gat), .B(G218gat), .Z(new_n257_));
  OAI211_X1 g056(.A(new_n257_), .B(KEYINPUT21), .C1(new_n247_), .C2(new_n249_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT78), .ZN(new_n260_));
  INV_X1    g059(.A(G176gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n228_), .A3(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT78), .B1(G169gat), .B2(G176gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT24), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT25), .B(G183gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(G190gat), .ZN(new_n267_));
  AOI22_X1  g066(.A1(new_n264_), .A2(new_n265_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n265_), .B1(G169gat), .B2(G176gat), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n269_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT79), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G183gat), .A2(G190gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT23), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(KEYINPUT80), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT80), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(G183gat), .A3(G190gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n274_), .B1(new_n278_), .B2(KEYINPUT23), .ZN(new_n279_));
  NAND4_X1  g078(.A1(new_n269_), .A2(new_n262_), .A3(KEYINPUT79), .A4(new_n263_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n268_), .A2(new_n272_), .A3(new_n279_), .A4(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n273_), .ZN(new_n282_));
  OR2_X1    g081(.A1(new_n282_), .A2(KEYINPUT23), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n275_), .A2(new_n277_), .A3(KEYINPUT23), .ZN(new_n284_));
  OR2_X1    g083(.A1(G183gat), .A2(G190gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n283_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(G169gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n259_), .A2(new_n281_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT20), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n279_), .A2(new_n285_), .ZN(new_n292_));
  OR2_X1    g091(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n294_));
  AND3_X1   g093(.A1(new_n293_), .A2(KEYINPUT93), .A3(new_n294_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT93), .B1(new_n293_), .B2(new_n294_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n261_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  OR3_X1    g096(.A1(new_n228_), .A2(new_n261_), .A3(KEYINPUT92), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT92), .B1(new_n228_), .B2(new_n261_), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n292_), .A2(new_n297_), .A3(new_n298_), .A4(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n267_), .A2(KEYINPUT91), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT91), .ZN(new_n302_));
  OR2_X1    g101(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n302_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n266_), .B1(new_n301_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n264_), .A2(new_n265_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n283_), .A2(new_n284_), .ZN(new_n308_));
  NAND4_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .A4(new_n270_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n259_), .B1(new_n300_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G226gat), .A2(G233gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n311_), .B(KEYINPUT90), .Z(new_n312_));
  XOR2_X1   g111(.A(new_n312_), .B(KEYINPUT19), .Z(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NOR3_X1   g113(.A1(new_n291_), .A2(new_n310_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT20), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n281_), .A2(new_n289_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n259_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n316_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n300_), .A2(new_n309_), .A3(new_n259_), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n313_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  OAI211_X1 g120(.A(KEYINPUT32), .B(new_n245_), .C1(new_n315_), .C2(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT98), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n314_), .B1(new_n291_), .B2(new_n310_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(KEYINPUT94), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n319_), .A2(new_n313_), .A3(new_n320_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT94), .ZN(new_n328_));
  OAI211_X1 g127(.A(new_n328_), .B(new_n314_), .C1(new_n291_), .C2(new_n310_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n326_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n245_), .A2(KEYINPUT32), .ZN(new_n332_));
  AOI22_X1  g131(.A1(new_n331_), .A2(new_n332_), .B1(new_n323_), .B2(new_n322_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G1gat), .B(G29gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(G85gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT0), .ZN(new_n336_));
  INV_X1    g135(.A(G57gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(G141gat), .A2(G148gat), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(G155gat), .A2(G162gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT83), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT1), .ZN(new_n345_));
  NOR2_X1   g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n341_), .B(new_n342_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n342_), .A2(KEYINPUT2), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT2), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(G141gat), .A3(G148gat), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(KEYINPUT84), .B(KEYINPUT3), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT85), .B1(new_n354_), .B2(new_n341_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT85), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT84), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(KEYINPUT3), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT3), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n359_), .A2(KEYINPUT84), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n356_), .B(new_n340_), .C1(new_n358_), .C2(new_n360_), .ZN(new_n361_));
  AOI211_X1 g160(.A(new_n349_), .B(new_n353_), .C1(new_n355_), .C2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n344_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n346_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n353_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n354_), .A2(KEYINPUT85), .A3(new_n341_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n359_), .A2(KEYINPUT84), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n357_), .A2(KEYINPUT3), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n356_), .B1(new_n370_), .B2(new_n340_), .ZN(new_n371_));
  OAI211_X1 g170(.A(new_n348_), .B(new_n366_), .C1(new_n367_), .C2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n365_), .B1(new_n372_), .B2(KEYINPUT86), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n347_), .B1(new_n364_), .B2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G127gat), .B(G134gat), .ZN(new_n375_));
  INV_X1    g174(.A(G113gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(new_n377_), .B(G120gat), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n374_), .A2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n372_), .A2(KEYINPUT86), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n349_), .B1(new_n355_), .B2(new_n361_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(new_n363_), .A3(new_n366_), .ZN(new_n383_));
  NAND4_X1  g182(.A1(new_n381_), .A2(new_n383_), .A3(new_n365_), .A4(new_n344_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(new_n378_), .A3(new_n347_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n380_), .A2(KEYINPUT4), .A3(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n374_), .A2(new_n387_), .A3(new_n379_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n386_), .A2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(G225gat), .A2(G233gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n389_), .A2(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(new_n380_), .B2(new_n385_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n339_), .B1(new_n392_), .B2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n390_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n396_), .A2(new_n338_), .A3(new_n393_), .ZN(new_n397_));
  OAI211_X1 g196(.A(new_n324_), .B(new_n333_), .C1(new_n395_), .C2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n386_), .A2(new_n390_), .A3(new_n388_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT97), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n380_), .A2(new_n391_), .A3(new_n385_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n402_), .A2(new_n339_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n386_), .A2(KEYINPUT97), .A3(new_n390_), .A4(new_n388_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n401_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n245_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n330_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT95), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n409_), .B1(new_n330_), .B2(new_n406_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n330_), .A2(new_n409_), .A3(new_n406_), .ZN(new_n412_));
  NAND4_X1  g211(.A1(new_n405_), .A2(new_n408_), .A3(new_n411_), .A4(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n338_), .B1(new_n396_), .B2(new_n393_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT96), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(KEYINPUT33), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  OAI221_X1 g216(.A(new_n338_), .B1(new_n415_), .B2(KEYINPUT33), .C1(new_n396_), .C2(new_n393_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  OAI21_X1  g218(.A(new_n398_), .B1(new_n413_), .B2(new_n419_), .ZN(new_n420_));
  OAI21_X1  g219(.A(G50gat), .B1(new_n374_), .B2(KEYINPUT29), .ZN(new_n421_));
  XOR2_X1   g220(.A(KEYINPUT28), .B(G22gat), .Z(new_n422_));
  INV_X1    g221(.A(KEYINPUT29), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n384_), .A2(new_n423_), .A3(new_n205_), .A4(new_n347_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n421_), .A2(new_n422_), .A3(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n422_), .B1(new_n421_), .B2(new_n424_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n259_), .B1(new_n374_), .B2(KEYINPUT29), .ZN(new_n428_));
  INV_X1    g227(.A(G228gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT87), .ZN(new_n430_));
  OR2_X1    g229(.A1(new_n430_), .A2(G233gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(G233gat), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n429_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT88), .ZN(new_n434_));
  XOR2_X1   g233(.A(G78gat), .B(G106gat), .Z(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n428_), .A2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n423_), .B1(new_n384_), .B2(new_n347_), .ZN(new_n439_));
  NOR3_X1   g238(.A1(new_n439_), .A2(new_n259_), .A3(new_n436_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT89), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n428_), .A2(new_n437_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT89), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n436_), .B1(new_n439_), .B2(new_n259_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n427_), .A2(new_n441_), .A3(new_n445_), .ZN(new_n446_));
  OAI221_X1 g245(.A(KEYINPUT89), .B1(new_n438_), .B2(new_n440_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n239_), .B1(new_n420_), .B2(new_n448_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n446_), .A2(new_n447_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n330_), .A2(new_n409_), .A3(new_n406_), .ZN(new_n451_));
  NOR3_X1   g250(.A1(new_n451_), .A2(new_n410_), .A3(new_n407_), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n452_), .A2(new_n417_), .A3(new_n405_), .A4(new_n418_), .ZN(new_n453_));
  AOI211_X1 g252(.A(KEYINPUT99), .B(new_n450_), .C1(new_n453_), .C2(new_n398_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n411_), .A2(new_n408_), .A3(new_n412_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT27), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n406_), .B1(new_n321_), .B2(new_n315_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n408_), .A2(KEYINPUT27), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n395_), .A2(new_n397_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NOR3_X1   g261(.A1(new_n460_), .A2(new_n462_), .A3(new_n448_), .ZN(new_n463_));
  NOR3_X1   g262(.A1(new_n449_), .A2(new_n454_), .A3(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n317_), .B(G43gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G71gat), .B(G99gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT30), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G227gat), .A2(G233gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(G15gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n467_), .B(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n465_), .B(new_n470_), .ZN(new_n471_));
  AND2_X1   g270(.A1(new_n471_), .A2(KEYINPUT81), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(KEYINPUT81), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n378_), .B(KEYINPUT31), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR3_X1   g274(.A1(new_n472_), .A2(new_n473_), .A3(new_n475_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n476_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT82), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n238_), .B1(new_n464_), .B2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n420_), .A2(new_n448_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(KEYINPUT99), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n460_), .A2(new_n448_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n461_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n420_), .A2(new_n239_), .A3(new_n448_), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n482_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n486_), .A2(KEYINPUT100), .A3(new_n478_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n480_), .A2(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n460_), .A2(new_n450_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT101), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(new_n461_), .A3(new_n477_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n237_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G99gat), .A2(G106gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT6), .ZN(new_n494_));
  OAI22_X1  g293(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(KEYINPUT65), .A2(KEYINPUT7), .ZN(new_n496_));
  INV_X1    g295(.A(G99gat), .ZN(new_n497_));
  INV_X1    g296(.A(G106gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n496_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n494_), .A2(new_n495_), .A3(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G85gat), .A2(G92gat), .ZN(new_n501_));
  INV_X1    g300(.A(G85gat), .ZN(new_n502_));
  INV_X1    g301(.A(G92gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n500_), .A2(new_n501_), .A3(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT66), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT66), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n500_), .A2(new_n507_), .A3(new_n501_), .A4(new_n504_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n506_), .A2(KEYINPUT8), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT8), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n505_), .A2(KEYINPUT66), .A3(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n504_), .A2(KEYINPUT9), .A3(new_n501_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n512_), .B1(KEYINPUT9), .B2(new_n501_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT64), .ZN(new_n514_));
  OR2_X1    g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT10), .B(G99gat), .Z(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n498_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n513_), .A2(new_n514_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n515_), .A2(new_n494_), .A3(new_n517_), .A4(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n509_), .A2(new_n511_), .A3(new_n519_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n520_), .A2(new_n207_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(KEYINPUT68), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT68), .ZN(new_n523_));
  NAND4_X1  g322(.A1(new_n509_), .A2(new_n523_), .A3(new_n511_), .A4(new_n519_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n522_), .A2(new_n524_), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n521_), .B1(new_n525_), .B2(new_n219_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G232gat), .A2(G233gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT34), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT35), .ZN(new_n530_));
  NOR2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  OR3_X1    g331(.A1(new_n526_), .A2(KEYINPUT70), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n529_), .A2(new_n530_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n526_), .A2(new_n534_), .A3(new_n532_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT70), .B1(new_n526_), .B2(new_n532_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n533_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G190gat), .B(G218gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(G134gat), .ZN(new_n539_));
  INV_X1    g338(.A(G162gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n539_), .B(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(KEYINPUT36), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n537_), .A2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n542_), .A2(KEYINPUT36), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NOR3_X1   g345(.A1(new_n537_), .A2(KEYINPUT36), .A3(new_n542_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n548_), .B(KEYINPUT103), .Z(new_n549_));
  NAND2_X1  g348(.A1(G231gat), .A2(G233gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n217_), .B(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G57gat), .B(G64gat), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(KEYINPUT11), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G71gat), .B(G78gat), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n554_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n555_), .B(new_n556_), .C1(KEYINPUT11), .C2(new_n552_), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n557_), .B(KEYINPUT67), .Z(new_n558_));
  XOR2_X1   g357(.A(new_n551_), .B(new_n558_), .Z(new_n559_));
  XNOR2_X1  g358(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G127gat), .B(G155gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XOR2_X1   g361(.A(G183gat), .B(G211gat), .Z(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n564_), .A2(KEYINPUT17), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(KEYINPUT17), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n559_), .A2(new_n565_), .A3(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(KEYINPUT74), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n551_), .B(new_n557_), .Z(new_n569_));
  NOR2_X1   g368(.A1(new_n569_), .A2(new_n566_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n549_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(G230gat), .A2(G233gat), .ZN(new_n574_));
  OAI21_X1  g373(.A(KEYINPUT12), .B1(new_n558_), .B2(new_n520_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n558_), .A2(new_n520_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT12), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n578_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n579_), .A2(KEYINPUT69), .A3(new_n557_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(KEYINPUT69), .B1(new_n579_), .B2(new_n557_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n574_), .B(new_n577_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n558_), .B(new_n520_), .Z(new_n584_));
  OAI21_X1  g383(.A(new_n583_), .B1(new_n574_), .B2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G120gat), .B(G148gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT5), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(G176gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(new_n248_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n585_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT13), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n492_), .A2(new_n573_), .A3(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(G1gat), .B1(new_n592_), .B2(new_n461_), .ZN(new_n593_));
  AND2_X1   g392(.A1(new_n548_), .A2(KEYINPUT37), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n548_), .A2(KEYINPUT37), .ZN(new_n595_));
  OR2_X1    g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n596_), .A2(new_n572_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n591_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT75), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n599_), .A2(new_n492_), .ZN(new_n600_));
  INV_X1    g399(.A(G1gat), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n462_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT102), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT38), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT102), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n600_), .A2(new_n605_), .A3(new_n601_), .A4(new_n462_), .ZN(new_n606_));
  AND3_X1   g405(.A1(new_n603_), .A2(new_n604_), .A3(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n604_), .B1(new_n603_), .B2(new_n606_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n593_), .B1(new_n607_), .B2(new_n608_), .ZN(G1324gat));
  INV_X1    g408(.A(G8gat), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n600_), .A2(new_n610_), .A3(new_n460_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n460_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G8gat), .B1(new_n592_), .B2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(KEYINPUT104), .B(KEYINPUT39), .Z(new_n614_));
  OR2_X1    g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n613_), .A2(new_n614_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n611_), .B1(new_n616_), .B2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(new_n618_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g418(.A1(new_n600_), .A2(new_n211_), .A3(new_n479_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT105), .Z(new_n621_));
  OAI21_X1  g420(.A(G15gat), .B1(new_n592_), .B2(new_n478_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT41), .Z(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(G1326gat));
  NAND3_X1  g423(.A1(new_n600_), .A2(new_n212_), .A3(new_n450_), .ZN(new_n625_));
  OAI21_X1  g424(.A(G22gat), .B1(new_n592_), .B2(new_n448_), .ZN(new_n626_));
  OR2_X1    g425(.A1(new_n626_), .A2(KEYINPUT106), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(KEYINPUT106), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n627_), .A2(KEYINPUT42), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(KEYINPUT42), .B1(new_n627_), .B2(new_n628_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n625_), .B1(new_n629_), .B2(new_n630_), .ZN(G1327gat));
  INV_X1    g430(.A(new_n549_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n632_), .A2(new_n571_), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n492_), .A2(new_n591_), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(G29gat), .B1(new_n634_), .B2(new_n462_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n486_), .A2(KEYINPUT100), .A3(new_n478_), .ZN(new_n636_));
  AOI21_X1  g435(.A(KEYINPUT100), .B1(new_n486_), .B2(new_n478_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n491_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n596_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT43), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n638_), .A2(KEYINPUT43), .A3(new_n596_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n641_), .A2(new_n572_), .A3(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n643_), .A2(KEYINPUT44), .A3(new_n591_), .A4(new_n236_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n644_), .A2(G29gat), .A3(new_n462_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n643_), .A2(new_n591_), .A3(new_n236_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT44), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n635_), .B1(new_n645_), .B2(new_n648_), .ZN(G1328gat));
  AOI21_X1  g448(.A(new_n612_), .B1(new_n646_), .B2(new_n647_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n644_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G36gat), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT45), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n492_), .A2(new_n591_), .A3(new_n633_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n654_), .A2(G36gat), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT107), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n655_), .A2(new_n656_), .A3(new_n460_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n656_), .B1(new_n655_), .B2(new_n460_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n653_), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n659_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(KEYINPUT45), .A3(new_n657_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n652_), .A2(new_n663_), .A3(KEYINPUT46), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  INV_X1    g464(.A(G36gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(new_n650_), .B2(new_n644_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n660_), .A2(new_n662_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n665_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n664_), .A2(new_n669_), .ZN(G1329gat));
  NAND4_X1  g469(.A1(new_n648_), .A2(G43gat), .A3(new_n477_), .A4(new_n644_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n203_), .B1(new_n654_), .B2(new_n478_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(KEYINPUT47), .ZN(new_n674_));
  INV_X1    g473(.A(KEYINPUT47), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n671_), .A2(new_n675_), .A3(new_n672_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n674_), .A2(new_n676_), .ZN(G1330gat));
  NAND4_X1  g476(.A1(new_n648_), .A2(G50gat), .A3(new_n450_), .A4(new_n644_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n205_), .B1(new_n654_), .B2(new_n448_), .ZN(new_n679_));
  AND2_X1   g478(.A1(new_n678_), .A2(new_n679_), .ZN(G1331gat));
  INV_X1    g479(.A(new_n591_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n597_), .A2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT108), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n236_), .B1(new_n488_), .B2(new_n491_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  AOI21_X1  g485(.A(G57gat), .B1(new_n686_), .B2(new_n462_), .ZN(new_n687_));
  NAND4_X1  g486(.A1(new_n638_), .A2(new_n573_), .A3(new_n681_), .A4(new_n237_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n688_), .A2(KEYINPUT109), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT109), .ZN(new_n690_));
  NAND4_X1  g489(.A1(new_n684_), .A2(new_n690_), .A3(new_n573_), .A4(new_n681_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n461_), .A2(new_n337_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n687_), .B1(new_n692_), .B2(new_n693_), .ZN(G1332gat));
  INV_X1    g493(.A(G64gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n686_), .A2(new_n695_), .A3(new_n460_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT48), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n692_), .A2(new_n460_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n697_), .B1(new_n698_), .B2(G64gat), .ZN(new_n699_));
  AOI211_X1 g498(.A(KEYINPUT48), .B(new_n695_), .C1(new_n692_), .C2(new_n460_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n696_), .B1(new_n699_), .B2(new_n700_), .ZN(G1333gat));
  INV_X1    g500(.A(new_n686_), .ZN(new_n702_));
  OR3_X1    g501(.A1(new_n702_), .A2(G71gat), .A3(new_n478_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n689_), .A2(new_n691_), .A3(new_n479_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT110), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(G71gat), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n705_), .B1(new_n704_), .B2(G71gat), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT49), .ZN(new_n709_));
  NOR3_X1   g508(.A1(new_n707_), .A2(new_n708_), .A3(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n704_), .A2(G71gat), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT110), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT49), .B1(new_n712_), .B2(new_n706_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n703_), .B1(new_n710_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT111), .B(new_n703_), .C1(new_n710_), .C2(new_n713_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(G1334gat));
  OR3_X1    g517(.A1(new_n702_), .A2(G78gat), .A3(new_n448_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n692_), .A2(new_n450_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n720_), .A2(new_n721_), .A3(G78gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n720_), .B2(G78gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1335gat));
  NAND3_X1  g523(.A1(new_n684_), .A2(new_n681_), .A3(new_n633_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n502_), .B1(new_n725_), .B2(new_n461_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n591_), .A2(new_n236_), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n641_), .A2(new_n572_), .A3(new_n642_), .A4(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n462_), .A2(G85gat), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n726_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(G1336gat));
  OAI21_X1  g530(.A(new_n503_), .B1(new_n725_), .B2(new_n612_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n460_), .A2(G92gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n728_), .B2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(G1337gat));
  OAI21_X1  g534(.A(G99gat), .B1(new_n728_), .B2(new_n478_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n477_), .A2(new_n516_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n736_), .B1(new_n725_), .B2(new_n737_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT113), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n738_), .B(new_n740_), .ZN(G1338gat));
  NAND4_X1  g540(.A1(new_n643_), .A2(KEYINPUT115), .A3(new_n450_), .A4(new_n727_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT115), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n743_), .B1(new_n728_), .B2(new_n448_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n742_), .A2(G106gat), .A3(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n725_), .A2(G106gat), .A3(new_n448_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT114), .Z(new_n749_));
  NAND4_X1  g548(.A1(new_n742_), .A2(KEYINPUT52), .A3(new_n744_), .A4(G106gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n747_), .A2(new_n749_), .A3(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(KEYINPUT53), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753_));
  NAND4_X1  g552(.A1(new_n747_), .A2(new_n749_), .A3(new_n753_), .A4(new_n750_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(G1339gat));
  NOR2_X1   g554(.A1(new_n585_), .A2(new_n589_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n525_), .A2(KEYINPUT12), .A3(new_n557_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT69), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(new_n759_));
  AOI22_X1  g558(.A1(new_n759_), .A2(new_n580_), .B1(new_n576_), .B2(new_n575_), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT116), .B1(new_n760_), .B2(new_n574_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n577_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT116), .ZN(new_n763_));
  INV_X1    g562(.A(new_n574_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n762_), .A2(new_n763_), .A3(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n583_), .A2(new_n766_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n760_), .A2(KEYINPUT55), .A3(new_n574_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n761_), .A2(new_n765_), .A3(new_n767_), .A4(new_n768_), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n589_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT56), .B1(new_n769_), .B2(new_n589_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n756_), .B1(new_n772_), .B2(KEYINPUT119), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT119), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n769_), .A2(new_n774_), .A3(KEYINPUT56), .A4(new_n589_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n220_), .A2(new_n224_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n223_), .A2(new_n221_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n234_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n232_), .A2(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT118), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n232_), .A2(KEYINPUT118), .A3(new_n778_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  AND2_X1   g582(.A1(new_n775_), .A2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n773_), .A2(KEYINPUT120), .A3(KEYINPUT58), .A4(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n594_), .A2(new_n595_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n761_), .A2(new_n765_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n767_), .A2(new_n768_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n589_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT56), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n769_), .A2(KEYINPUT56), .A3(new_n589_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(KEYINPUT119), .A3(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n756_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n784_), .A3(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT58), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n786_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n793_), .A2(new_n784_), .A3(KEYINPUT58), .A4(new_n794_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n785_), .A2(new_n797_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n794_), .A2(new_n236_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n791_), .A2(KEYINPUT117), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT117), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n771_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n802_), .B1(new_n806_), .B2(new_n792_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n590_), .A2(new_n783_), .ZN(new_n808_));
  OAI211_X1 g607(.A(KEYINPUT57), .B(new_n632_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n804_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n811_));
  AOI211_X1 g610(.A(KEYINPUT117), .B(KEYINPUT56), .C1(new_n769_), .C2(new_n589_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n792_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n802_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n808_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n810_), .B1(new_n815_), .B2(new_n549_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n801_), .A2(new_n809_), .A3(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(new_n572_), .ZN(new_n818_));
  OAI21_X1  g617(.A(KEYINPUT54), .B1(new_n598_), .B2(new_n236_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n597_), .A2(new_n820_), .A3(new_n591_), .A4(new_n237_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n818_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n490_), .A2(new_n477_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n823_), .A2(new_n462_), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT121), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n461_), .B1(new_n818_), .B2(new_n822_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(KEYINPUT121), .A3(new_n825_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(G113gat), .B1(new_n831_), .B2(new_n236_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT59), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n829_), .A2(new_n833_), .A3(new_n825_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n833_), .B1(new_n829_), .B2(new_n825_), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n237_), .A2(new_n376_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n832_), .B1(new_n837_), .B2(new_n838_), .ZN(G1340gat));
  NOR2_X1   g638(.A1(new_n591_), .A2(G120gat), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(KEYINPUT60), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n826_), .A2(KEYINPUT59), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(new_n681_), .A3(new_n834_), .ZN(new_n844_));
  OAI21_X1  g643(.A(G120gat), .B1(new_n842_), .B2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n842_), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n845_), .B1(new_n846_), .B2(KEYINPUT60), .ZN(G1341gat));
  AOI21_X1  g646(.A(G127gat), .B1(new_n831_), .B2(new_n571_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n571_), .A2(G127gat), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n848_), .B1(new_n837_), .B2(new_n849_), .ZN(G1342gat));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n786_), .A2(new_n851_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT123), .ZN(new_n853_));
  NOR3_X1   g652(.A1(new_n835_), .A2(new_n836_), .A3(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n632_), .B1(new_n828_), .B2(new_n830_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(G134gat), .ZN(new_n857_));
  AOI21_X1  g656(.A(KEYINPUT121), .B1(new_n829_), .B2(new_n825_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n572_), .A2(new_n817_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n859_));
  NOR4_X1   g658(.A1(new_n859_), .A2(new_n827_), .A3(new_n461_), .A4(new_n824_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n549_), .B1(new_n858_), .B2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(KEYINPUT122), .A3(new_n851_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n854_), .B1(new_n857_), .B2(new_n862_), .ZN(G1343gat));
  AND4_X1   g662(.A1(new_n462_), .A2(new_n823_), .A3(new_n478_), .A4(new_n483_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n236_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n681_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g667(.A1(new_n864_), .A2(new_n571_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(KEYINPUT61), .B(G155gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1346gat));
  AOI21_X1  g670(.A(G162gat), .B1(new_n864_), .B2(new_n549_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n786_), .A2(new_n540_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n872_), .B1(new_n864_), .B2(new_n873_), .ZN(G1347gat));
  NOR3_X1   g673(.A1(new_n859_), .A2(new_n462_), .A3(new_n612_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n295_), .A2(new_n296_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n478_), .A2(new_n450_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n875_), .A2(new_n236_), .A3(new_n876_), .A4(new_n877_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n612_), .A2(new_n462_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n823_), .A2(new_n879_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n877_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n880_), .A2(new_n237_), .A3(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n878_), .B1(new_n882_), .B2(new_n228_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT62), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n882_), .A2(new_n228_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n884_), .B1(KEYINPUT62), .B2(new_n885_), .ZN(G1348gat));
  NOR2_X1   g685(.A1(new_n880_), .A2(new_n881_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n681_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g688(.A1(new_n887_), .A2(new_n571_), .ZN(new_n890_));
  MUX2_X1   g689(.A(new_n266_), .B(G183gat), .S(new_n890_), .Z(G1350gat));
  OAI211_X1 g690(.A(new_n887_), .B(new_n549_), .C1(new_n305_), .C2(new_n301_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n880_), .A2(new_n786_), .A3(new_n881_), .ZN(new_n893_));
  INV_X1    g692(.A(G190gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1351gat));
  NOR2_X1   g694(.A1(new_n479_), .A2(new_n448_), .ZN(new_n896_));
  AND3_X1   g695(.A1(new_n823_), .A2(new_n879_), .A3(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n236_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G197gat), .ZN(G1352gat));
  AND2_X1   g698(.A1(new_n897_), .A2(new_n681_), .ZN(new_n900_));
  AND2_X1   g699(.A1(new_n248_), .A2(KEYINPUT124), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n248_), .A2(KEYINPUT124), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n900_), .B2(new_n901_), .ZN(G1353gat));
  XOR2_X1   g703(.A(KEYINPUT63), .B(G211gat), .Z(new_n905_));
  NAND4_X1  g704(.A1(new_n897_), .A2(KEYINPUT125), .A3(new_n571_), .A4(new_n905_), .ZN(new_n906_));
  NAND4_X1  g705(.A1(new_n823_), .A2(new_n571_), .A3(new_n879_), .A4(new_n896_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(new_n909_));
  INV_X1    g708(.A(KEYINPUT125), .ZN(new_n910_));
  INV_X1    g709(.A(new_n905_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n907_), .B2(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n906_), .A2(new_n909_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(KEYINPUT126), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n915_));
  NAND4_X1  g714(.A1(new_n906_), .A2(new_n915_), .A3(new_n912_), .A4(new_n909_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1354gat));
  XOR2_X1   g716(.A(KEYINPUT127), .B(G218gat), .Z(new_n918_));
  AOI21_X1  g717(.A(new_n918_), .B1(new_n897_), .B2(new_n549_), .ZN(new_n919_));
  AND2_X1   g718(.A1(new_n596_), .A2(new_n918_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n897_), .B2(new_n920_), .ZN(G1355gat));
endmodule


