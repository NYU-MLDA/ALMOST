//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 1 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:41 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n929_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n940_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_;
  INV_X1    g000(.A(KEYINPUT3), .ZN(new_n202_));
  INV_X1    g001(.A(G141gat), .ZN(new_n203_));
  INV_X1    g002(.A(G148gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT2), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G155gat), .B(G162gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  AND2_X1   g013(.A1(G141gat), .A2(G148gat), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n217_), .B(new_n218_), .C1(new_n212_), .C2(KEYINPUT1), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n214_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT89), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT95), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n214_), .A2(KEYINPUT89), .A3(new_n219_), .ZN(new_n224_));
  XNOR2_X1  g023(.A(G127gat), .B(G134gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(G113gat), .B(G120gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .A4(new_n228_), .ZN(new_n229_));
  AND3_X1   g028(.A1(new_n214_), .A2(KEYINPUT89), .A3(new_n219_), .ZN(new_n230_));
  AOI21_X1  g029(.A(KEYINPUT89), .B1(new_n214_), .B2(new_n219_), .ZN(new_n231_));
  NOR3_X1   g030(.A1(new_n230_), .A2(new_n231_), .A3(new_n227_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT95), .B1(new_n228_), .B2(new_n220_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n229_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT4), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G225gat), .A2(G233gat), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n230_), .A2(new_n231_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT4), .ZN(new_n239_));
  NAND4_X1  g038(.A1(new_n238_), .A2(KEYINPUT96), .A3(new_n239_), .A4(new_n228_), .ZN(new_n240_));
  NAND4_X1  g039(.A1(new_n222_), .A2(new_n239_), .A3(new_n224_), .A4(new_n228_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT96), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n240_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n235_), .A2(new_n237_), .A3(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n234_), .A2(new_n236_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G1gat), .B(G29gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(G85gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT0), .B(G57gat), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n248_), .B(new_n249_), .Z(new_n250_));
  NAND3_X1  g049(.A1(new_n245_), .A2(new_n246_), .A3(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT101), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n245_), .A2(new_n246_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n250_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT101), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n245_), .A2(new_n256_), .A3(new_n246_), .A4(new_n250_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n252_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n258_));
  XNOR2_X1  g057(.A(G8gat), .B(G36gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT18), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G64gat), .B(G92gat), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n260_), .B(new_n261_), .Z(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT19), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT84), .ZN(new_n266_));
  INV_X1    g065(.A(G169gat), .ZN(new_n267_));
  INV_X1    g066(.A(G176gat), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(KEYINPUT83), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT83), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n270_), .B1(G169gat), .B2(G176gat), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G169gat), .A2(G176gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT24), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n266_), .B1(new_n272_), .B2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n274_), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n276_), .A2(KEYINPUT84), .A3(new_n269_), .A4(new_n271_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT81), .ZN(new_n279_));
  INV_X1    g078(.A(G183gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n279_), .B1(new_n280_), .B2(KEYINPUT25), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT25), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(KEYINPUT81), .A3(G183gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n281_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n280_), .A2(KEYINPUT80), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT80), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n286_), .A2(G183gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n285_), .A2(new_n287_), .A3(KEYINPUT25), .ZN(new_n288_));
  XNOR2_X1  g087(.A(KEYINPUT26), .B(G190gat), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n284_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT82), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT24), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n294_), .B1(new_n295_), .B2(new_n272_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT82), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n284_), .A2(new_n288_), .A3(new_n297_), .A4(new_n289_), .ZN(new_n298_));
  NAND4_X1  g097(.A1(new_n278_), .A2(new_n291_), .A3(new_n296_), .A4(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(KEYINPUT85), .B(G176gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT22), .B(G169gat), .ZN(new_n301_));
  AOI22_X1  g100(.A1(new_n300_), .A2(new_n301_), .B1(G169gat), .B2(G176gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n285_), .A2(new_n287_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n303_), .A2(G190gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n302_), .B1(new_n294_), .B2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G211gat), .B(G218gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(G204gat), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(KEYINPUT90), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT90), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(G204gat), .ZN(new_n311_));
  INV_X1    g110(.A(G197gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n309_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT21), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n314_), .B1(G197gat), .B2(G204gat), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n307_), .B1(new_n313_), .B2(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n312_), .B1(new_n309_), .B2(new_n311_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(G197gat), .A2(G204gat), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n314_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n317_), .A2(new_n318_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n306_), .A2(new_n314_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n316_), .A2(new_n319_), .B1(new_n320_), .B2(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n299_), .A2(new_n305_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT20), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n273_), .A2(KEYINPUT91), .A3(KEYINPUT24), .ZN(new_n325_));
  AOI21_X1  g124(.A(KEYINPUT91), .B1(new_n273_), .B2(KEYINPUT24), .ZN(new_n326_));
  NOR3_X1   g125(.A1(new_n272_), .A2(new_n325_), .A3(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n282_), .A2(G183gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n280_), .A2(KEYINPUT25), .ZN(new_n329_));
  AND3_X1   g128(.A1(new_n289_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT92), .B1(new_n327_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n326_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n273_), .A2(KEYINPUT91), .A3(KEYINPUT24), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n332_), .A2(new_n271_), .A3(new_n269_), .A4(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT92), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n289_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n334_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  NOR3_X1   g136(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n294_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n331_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G183gat), .A2(G190gat), .ZN(new_n341_));
  OAI21_X1  g140(.A(new_n302_), .B1(new_n294_), .B2(new_n341_), .ZN(new_n342_));
  AOI21_X1  g141(.A(new_n322_), .B1(new_n340_), .B2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n265_), .B1(new_n324_), .B2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n299_), .A2(new_n305_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n322_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n340_), .A2(new_n322_), .A3(new_n342_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT93), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT20), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n265_), .A2(new_n350_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n347_), .A2(new_n348_), .A3(new_n349_), .A4(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n344_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n351_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n349_), .B1(new_n355_), .B2(new_n348_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n263_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n347_), .A2(new_n348_), .A3(new_n351_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT93), .ZN(new_n359_));
  NAND4_X1  g158(.A1(new_n359_), .A2(new_n262_), .A3(new_n344_), .A4(new_n352_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT27), .B1(new_n357_), .B2(new_n360_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n324_), .A2(new_n343_), .A3(new_n265_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n265_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n350_), .B1(new_n345_), .B2(new_n346_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(new_n348_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n263_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n360_), .A2(new_n366_), .A3(KEYINPUT27), .ZN(new_n367_));
  XOR2_X1   g166(.A(G78gat), .B(G106gat), .Z(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  AND2_X1   g168(.A1(new_n214_), .A2(new_n219_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT29), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  OAI211_X1 g171(.A(G228gat), .B(G233gat), .C1(new_n372_), .C2(new_n322_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n222_), .A2(KEYINPUT29), .A3(new_n224_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G228gat), .A2(G233gat), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n375_), .A3(new_n346_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n369_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  OAI21_X1  g177(.A(KEYINPUT28), .B1(new_n238_), .B2(KEYINPUT29), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n222_), .A2(new_n224_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT28), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n380_), .A2(new_n381_), .A3(new_n371_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G22gat), .B(G50gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n384_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n379_), .A2(new_n382_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n373_), .A2(new_n376_), .A3(new_n369_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n378_), .A2(new_n385_), .A3(new_n387_), .A4(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n387_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n386_), .B1(new_n379_), .B2(new_n382_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n373_), .A2(new_n376_), .A3(new_n369_), .ZN(new_n392_));
  OAI22_X1  g191(.A1(new_n390_), .A2(new_n391_), .B1(new_n392_), .B2(new_n377_), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n389_), .A2(new_n393_), .ZN(new_n394_));
  NOR4_X1   g193(.A1(new_n258_), .A2(new_n361_), .A3(new_n367_), .A4(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n262_), .A2(KEYINPUT32), .ZN(new_n396_));
  NOR3_X1   g195(.A1(new_n362_), .A2(new_n365_), .A3(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT100), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n359_), .A2(new_n344_), .A3(new_n352_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n397_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n396_), .B1(new_n399_), .B2(KEYINPUT100), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n258_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n357_), .A2(new_n360_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT94), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n357_), .A2(KEYINPUT94), .A3(new_n360_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT99), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n234_), .A2(KEYINPUT4), .B1(new_n240_), .B2(new_n243_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n409_), .B2(new_n236_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n408_), .A3(new_n236_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n222_), .A2(new_n224_), .A3(new_n228_), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n223_), .B1(new_n370_), .B2(new_n227_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  AOI21_X1  g214(.A(new_n236_), .B1(new_n415_), .B2(new_n229_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT98), .B1(new_n416_), .B2(new_n250_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n234_), .A2(new_n237_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT98), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n418_), .A2(new_n419_), .A3(new_n254_), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n411_), .A2(new_n412_), .A3(new_n417_), .A4(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n406_), .A2(new_n407_), .A3(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n251_), .A2(KEYINPUT97), .A3(KEYINPUT33), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT33), .B1(new_n251_), .B2(KEYINPUT97), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n403_), .B1(new_n422_), .B2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n395_), .B1(new_n426_), .B2(new_n394_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G71gat), .B(G99gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n428_), .B(G43gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n345_), .B(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(G227gat), .A2(G233gat), .ZN(new_n431_));
  INV_X1    g230(.A(G15gat), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT30), .ZN(new_n434_));
  OR2_X1    g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  XOR2_X1   g234(.A(new_n227_), .B(KEYINPUT31), .Z(new_n436_));
  NAND2_X1  g235(.A1(new_n430_), .A2(new_n434_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n435_), .A2(new_n436_), .A3(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(KEYINPUT88), .ZN(new_n439_));
  XOR2_X1   g238(.A(new_n436_), .B(KEYINPUT87), .Z(new_n440_));
  NAND2_X1  g239(.A1(new_n435_), .A2(new_n437_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT86), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n443_), .B1(new_n442_), .B2(new_n441_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(KEYINPUT102), .B1(new_n427_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n445_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n394_), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n258_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n361_), .A2(new_n367_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n449_), .A2(new_n450_), .A3(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT102), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n420_), .A2(new_n417_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n454_), .A2(new_n410_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n405_), .A2(new_n404_), .B1(new_n455_), .B2(new_n412_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n251_), .A2(KEYINPUT97), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT33), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n251_), .A2(KEYINPUT97), .A3(KEYINPUT33), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n456_), .A2(new_n461_), .A3(new_n407_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n448_), .B1(new_n462_), .B2(new_n403_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n453_), .B(new_n447_), .C1(new_n463_), .C2(new_n395_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n446_), .A2(new_n452_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT105), .ZN(new_n466_));
  XOR2_X1   g265(.A(G85gat), .B(G92gat), .Z(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT9), .ZN(new_n468_));
  NAND2_X1  g267(.A1(G99gat), .A2(G106gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT6), .ZN(new_n470_));
  INV_X1    g269(.A(G85gat), .ZN(new_n471_));
  INV_X1    g270(.A(G92gat), .ZN(new_n472_));
  OR3_X1    g271(.A1(new_n471_), .A2(new_n472_), .A3(KEYINPUT9), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n468_), .A2(new_n470_), .A3(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(KEYINPUT10), .B(G99gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT64), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n474_), .B1(G106gat), .B2(new_n476_), .ZN(new_n477_));
  OR3_X1    g276(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(KEYINPUT65), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT65), .ZN(new_n481_));
  OAI211_X1 g280(.A(new_n481_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n470_), .A2(new_n478_), .A3(new_n480_), .A4(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT66), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n483_), .B(new_n467_), .C1(new_n484_), .C2(KEYINPUT8), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n467_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT8), .B1(new_n467_), .B2(new_n484_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n477_), .A2(new_n485_), .A3(new_n488_), .ZN(new_n489_));
  XOR2_X1   g288(.A(G29gat), .B(G36gat), .Z(new_n490_));
  XOR2_X1   g289(.A(G43gat), .B(G50gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT15), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n489_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT70), .ZN(new_n495_));
  XOR2_X1   g294(.A(KEYINPUT69), .B(KEYINPUT34), .Z(new_n496_));
  NAND2_X1  g295(.A1(G232gat), .A2(G233gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT35), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n495_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n492_), .ZN(new_n501_));
  OAI211_X1 g300(.A(new_n494_), .B(new_n500_), .C1(new_n489_), .C2(new_n501_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n498_), .A2(new_n499_), .ZN(new_n503_));
  OR2_X1    g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(G190gat), .B(G218gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G134gat), .B(G162gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n507_), .A2(KEYINPUT36), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n502_), .A2(new_n503_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n504_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT71), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n504_), .A2(new_n509_), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n507_), .B(KEYINPUT36), .Z(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n515_), .A2(KEYINPUT72), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(KEYINPUT72), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n512_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  AND3_X1   g317(.A1(new_n465_), .A2(new_n466_), .A3(new_n518_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n466_), .B1(new_n465_), .B2(new_n518_), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT73), .B(G1gat), .ZN(new_n522_));
  INV_X1    g321(.A(G8gat), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT14), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G1gat), .B(G8gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n524_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n493_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n529_), .A2(new_n530_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(new_n492_), .ZN(new_n535_));
  AND3_X1   g334(.A1(new_n532_), .A2(new_n533_), .A3(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n531_), .A2(new_n501_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n537_), .A2(KEYINPUT76), .A3(new_n535_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n533_), .ZN(new_n539_));
  OR3_X1    g338(.A1(new_n534_), .A2(KEYINPUT76), .A3(new_n492_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT77), .ZN(new_n542_));
  OR2_X1    g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n541_), .A2(new_n542_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n536_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT79), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G113gat), .B(G141gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT78), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G169gat), .B(G197gat), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n548_), .B(new_n549_), .Z(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  OR3_X1    g350(.A1(new_n545_), .A2(new_n546_), .A3(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n545_), .B2(new_n546_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT104), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT11), .ZN(new_n558_));
  XOR2_X1   g357(.A(G71gat), .B(G78gat), .Z(new_n559_));
  OR2_X1    g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n557_), .A2(KEYINPUT11), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n559_), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n560_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n489_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT12), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(G230gat), .A2(G233gat), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n477_), .A2(new_n488_), .A3(new_n485_), .A4(new_n563_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n563_), .A2(KEYINPUT67), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT67), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n560_), .B(new_n571_), .C1(new_n561_), .C2(new_n562_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(new_n489_), .A3(KEYINPUT12), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n567_), .A2(new_n568_), .A3(new_n569_), .A4(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n565_), .A2(new_n569_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n568_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(G120gat), .B(G148gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(G176gat), .B(G204gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n579_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n575_), .A2(new_n578_), .A3(new_n584_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT13), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n586_), .A2(KEYINPUT13), .A3(new_n587_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n555_), .A2(new_n556_), .A3(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(G127gat), .B(G155gat), .Z(new_n595_));
  XNOR2_X1  g394(.A(G183gat), .B(G211gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n595_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT17), .ZN(new_n600_));
  AND2_X1   g399(.A1(G231gat), .A2(G233gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n534_), .B(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n600_), .B1(new_n603_), .B2(new_n563_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n604_), .B1(new_n603_), .B2(new_n563_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n599_), .A2(KEYINPUT17), .ZN(new_n606_));
  INV_X1    g405(.A(new_n573_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n606_), .B1(new_n602_), .B2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n608_), .B1(new_n602_), .B2(new_n607_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n605_), .A2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(KEYINPUT104), .B1(new_n554_), .B2(new_n592_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n594_), .A2(new_n610_), .A3(new_n611_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n521_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(new_n258_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(G1gat), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT37), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n616_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n518_), .A2(new_n616_), .B1(new_n512_), .B2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n610_), .B(KEYINPUT75), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NOR3_X1   g420(.A1(new_n619_), .A2(new_n592_), .A3(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n465_), .A2(new_n555_), .A3(new_n622_), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n258_), .A2(KEYINPUT103), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n258_), .A2(KEYINPUT103), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n623_), .A2(new_n522_), .A3(new_n627_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT38), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n615_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT106), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n615_), .A2(KEYINPUT106), .A3(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(G1324gat));
  INV_X1    g433(.A(new_n451_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n623_), .A2(new_n523_), .A3(new_n635_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n635_), .B(new_n612_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT107), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n637_), .A2(new_n638_), .A3(G8gat), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n638_), .B1(new_n637_), .B2(G8gat), .ZN(new_n641_));
  NOR3_X1   g440(.A1(new_n640_), .A2(new_n641_), .A3(KEYINPUT39), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n637_), .A2(G8gat), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(KEYINPUT107), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n643_), .B1(new_n645_), .B2(new_n639_), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n636_), .B1(new_n642_), .B2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  OAI211_X1 g448(.A(KEYINPUT40), .B(new_n636_), .C1(new_n642_), .C2(new_n646_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1325gat));
  NAND3_X1  g450(.A1(new_n623_), .A2(new_n432_), .A3(new_n445_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n613_), .A2(new_n445_), .ZN(new_n653_));
  AND3_X1   g452(.A1(new_n653_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n654_));
  AOI21_X1  g453(.A(KEYINPUT41), .B1(new_n653_), .B2(G15gat), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n652_), .B1(new_n654_), .B2(new_n655_), .ZN(G1326gat));
  INV_X1    g455(.A(G22gat), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n448_), .A2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT108), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n623_), .A2(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n613_), .A2(new_n448_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n662_), .B2(G22gat), .ZN(new_n663_));
  AOI211_X1 g462(.A(KEYINPUT42), .B(new_n657_), .C1(new_n613_), .C2(new_n448_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n660_), .B1(new_n663_), .B2(new_n664_), .ZN(G1327gat));
  NOR3_X1   g464(.A1(new_n518_), .A2(new_n620_), .A3(new_n592_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n465_), .A2(new_n555_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT112), .ZN(new_n668_));
  OR2_X1    g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n667_), .A2(new_n668_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(G29gat), .B1(new_n671_), .B2(new_n258_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n465_), .A2(new_n619_), .ZN(new_n673_));
  XOR2_X1   g472(.A(KEYINPUT109), .B(KEYINPUT43), .Z(new_n674_));
  NAND2_X1  g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n465_), .B(new_n619_), .C1(KEYINPUT109), .C2(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n594_), .A2(new_n611_), .A3(new_n621_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT44), .ZN(new_n682_));
  OAI21_X1  g481(.A(KEYINPUT111), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n679_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT111), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n684_), .A2(new_n685_), .A3(KEYINPUT44), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n683_), .A2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(KEYINPUT110), .B(KEYINPUT44), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n681_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n687_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n627_), .A2(G29gat), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n672_), .B1(new_n692_), .B2(new_n693_), .ZN(G1328gat));
  INV_X1    g493(.A(G36gat), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n669_), .A2(new_n695_), .A3(new_n635_), .A4(new_n670_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT45), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n684_), .A2(new_n688_), .ZN(new_n698_));
  AOI211_X1 g497(.A(new_n451_), .B(new_n698_), .C1(new_n683_), .C2(new_n686_), .ZN(new_n699_));
  OAI211_X1 g498(.A(new_n697_), .B(KEYINPUT46), .C1(new_n699_), .C2(new_n695_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT46), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n698_), .A2(new_n451_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n695_), .B1(new_n687_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n697_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n701_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n700_), .A2(new_n705_), .ZN(G1329gat));
  NAND2_X1  g505(.A1(new_n445_), .A2(G43gat), .ZN(new_n707_));
  AOI211_X1 g506(.A(new_n698_), .B(new_n707_), .C1(new_n683_), .C2(new_n686_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n671_), .A2(new_n445_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(KEYINPUT113), .B(G43gat), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n711_), .ZN(new_n712_));
  OAI21_X1  g511(.A(KEYINPUT47), .B1(new_n708_), .B2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n714_), .B(new_n711_), .C1(new_n691_), .C2(new_n707_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1330gat));
  INV_X1    g515(.A(G50gat), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n671_), .A2(new_n717_), .A3(new_n448_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n698_), .A2(new_n394_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n687_), .A2(new_n719_), .ZN(new_n720_));
  AOI21_X1  g519(.A(KEYINPUT114), .B1(new_n720_), .B2(G50gat), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT114), .ZN(new_n722_));
  AOI211_X1 g521(.A(new_n722_), .B(new_n717_), .C1(new_n687_), .C2(new_n719_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n718_), .B1(new_n721_), .B2(new_n723_), .ZN(G1331gat));
  NAND2_X1  g523(.A1(new_n465_), .A2(new_n554_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n620_), .A2(new_n592_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n725_), .A2(new_n619_), .A3(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(G57gat), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n727_), .A2(new_n728_), .A3(new_n627_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n726_), .A2(new_n555_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n521_), .A2(new_n258_), .A3(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n729_), .B1(new_n731_), .B2(new_n728_), .ZN(G1332gat));
  INV_X1    g531(.A(G64gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n727_), .A2(new_n733_), .A3(new_n635_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n521_), .A2(new_n635_), .A3(new_n730_), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT48), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(new_n736_), .A3(G64gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n735_), .B2(G64gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n734_), .B1(new_n737_), .B2(new_n738_), .ZN(G1333gat));
  NOR2_X1   g538(.A1(new_n447_), .A2(G71gat), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT115), .Z(new_n741_));
  NAND2_X1  g540(.A1(new_n727_), .A2(new_n741_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n521_), .A2(new_n445_), .A3(new_n730_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT49), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n743_), .A2(new_n744_), .A3(G71gat), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n744_), .B1(new_n743_), .B2(G71gat), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n742_), .B1(new_n745_), .B2(new_n746_), .ZN(G1334gat));
  INV_X1    g546(.A(G78gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n727_), .A2(new_n748_), .A3(new_n448_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n521_), .A2(new_n448_), .A3(new_n730_), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT50), .ZN(new_n751_));
  AND3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(G78gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n751_), .B1(new_n750_), .B2(G78gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n749_), .B1(new_n752_), .B2(new_n753_), .ZN(G1335gat));
  NAND2_X1  g553(.A1(new_n621_), .A2(new_n592_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n755_), .A2(new_n555_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759_), .B2(new_n450_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n725_), .A2(new_n518_), .A3(new_n755_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n471_), .A3(new_n627_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1336gat));
  OAI21_X1  g562(.A(G92gat), .B1(new_n759_), .B2(new_n451_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n761_), .A2(new_n472_), .A3(new_n635_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1337gat));
  INV_X1    g565(.A(G99gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n767_), .B1(new_n758_), .B2(new_n445_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n755_), .A2(new_n518_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n447_), .A2(new_n476_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n465_), .A2(new_n554_), .A3(new_n769_), .A4(new_n770_), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n771_), .A2(KEYINPUT116), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n771_), .A2(KEYINPUT116), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  NOR3_X1   g573(.A1(new_n768_), .A2(new_n774_), .A3(KEYINPUT117), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT117), .B1(new_n768_), .B2(new_n774_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT118), .ZN(new_n778_));
  NAND4_X1  g577(.A1(new_n776_), .A2(new_n777_), .A3(new_n778_), .A4(KEYINPUT51), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n758_), .A2(new_n445_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n780_), .A2(G99gat), .B1(new_n772_), .B2(new_n773_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n778_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n777_), .A2(KEYINPUT51), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n775_), .ZN(new_n785_));
  AND2_X1   g584(.A1(new_n779_), .A2(new_n785_), .ZN(G1338gat));
  INV_X1    g585(.A(G106gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n761_), .A2(new_n787_), .A3(new_n448_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n758_), .A2(new_n448_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(G106gat), .ZN(new_n791_));
  AOI211_X1 g590(.A(KEYINPUT52), .B(new_n787_), .C1(new_n758_), .C2(new_n448_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n788_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g593(.A1(new_n622_), .A2(new_n554_), .ZN(new_n795_));
  XNOR2_X1  g594(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n795_), .B(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n518_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n538_), .A2(new_n540_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(new_n533_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n532_), .A2(new_n535_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n539_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n551_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n545_), .B2(new_n551_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n588_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT121), .ZN(new_n806_));
  XNOR2_X1  g605(.A(new_n805_), .B(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n587_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n808_), .B1(new_n552_), .B2(new_n553_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n574_), .A2(new_n569_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT12), .B1(new_n489_), .B2(new_n564_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n577_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n812_), .A2(KEYINPUT55), .A3(new_n575_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n810_), .A2(new_n811_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n814_), .A2(new_n815_), .A3(new_n568_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT120), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT120), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n813_), .A2(new_n819_), .A3(new_n816_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n818_), .A2(KEYINPUT56), .A3(new_n585_), .A4(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n584_), .B1(new_n817_), .B2(KEYINPUT120), .ZN(new_n823_));
  AOI21_X1  g622(.A(KEYINPUT56), .B1(new_n823_), .B2(new_n820_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n809_), .B1(new_n822_), .B2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n798_), .B1(new_n807_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT57), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n827_), .A2(KEYINPUT124), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT124), .B(KEYINPUT57), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n798_), .B(new_n830_), .C1(new_n807_), .C2(new_n825_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n829_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT122), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n821_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n818_), .A2(new_n585_), .A3(new_n820_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n823_), .A2(KEYINPUT122), .A3(KEYINPUT56), .A4(new_n820_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n834_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n804_), .A2(new_n587_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n618_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n839_), .A2(KEYINPUT58), .A3(new_n840_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n832_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n621_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n797_), .A2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n449_), .A2(new_n627_), .A3(new_n451_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n849_), .A2(KEYINPUT59), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n843_), .A2(KEYINPUT123), .A3(new_n844_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT123), .B1(new_n843_), .B2(new_n844_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n832_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT125), .ZN(new_n855_));
  INV_X1    g654(.A(new_n610_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT125), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n832_), .B(new_n857_), .C1(new_n852_), .C2(new_n853_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n855_), .A2(new_n856_), .A3(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n849_), .B1(new_n859_), .B2(new_n797_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT59), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n851_), .B1(new_n860_), .B2(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(G113gat), .B1(new_n862_), .B2(new_n554_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n830_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n826_), .A2(new_n864_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n845_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n843_), .A2(KEYINPUT123), .A3(new_n844_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n866_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n856_), .B1(new_n870_), .B2(new_n857_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n858_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n797_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n849_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  OR3_X1    g674(.A1(new_n875_), .A2(G113gat), .A3(new_n554_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n863_), .A2(new_n876_), .ZN(G1340gat));
  OAI21_X1  g676(.A(G120gat), .B1(new_n862_), .B2(new_n593_), .ZN(new_n878_));
  INV_X1    g677(.A(G120gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n593_), .B2(KEYINPUT60), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n860_), .B(new_n880_), .C1(KEYINPUT60), .C2(new_n879_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n878_), .A2(new_n881_), .ZN(G1341gat));
  OAI21_X1  g681(.A(G127gat), .B1(new_n862_), .B2(new_n856_), .ZN(new_n883_));
  OR3_X1    g682(.A1(new_n875_), .A2(G127gat), .A3(new_n621_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(G1342gat));
  AOI211_X1 g684(.A(new_n518_), .B(new_n849_), .C1(new_n859_), .C2(new_n797_), .ZN(new_n886_));
  OAI21_X1  g685(.A(KEYINPUT126), .B1(new_n886_), .B2(G134gat), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT126), .ZN(new_n888_));
  INV_X1    g687(.A(G134gat), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n888_), .B(new_n889_), .C1(new_n875_), .C2(new_n518_), .ZN(new_n890_));
  AOI22_X1  g689(.A1(new_n875_), .A2(KEYINPUT59), .B1(new_n848_), .B2(new_n850_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n618_), .A2(new_n889_), .ZN(new_n892_));
  AOI22_X1  g691(.A1(new_n887_), .A2(new_n890_), .B1(new_n891_), .B2(new_n892_), .ZN(G1343gat));
  NOR4_X1   g692(.A1(new_n626_), .A2(new_n445_), .A3(new_n394_), .A4(new_n635_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n873_), .A2(new_n894_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n203_), .A3(new_n555_), .ZN(new_n897_));
  OAI21_X1  g696(.A(G141gat), .B1(new_n895_), .B2(new_n554_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n897_), .A2(new_n898_), .ZN(G1344gat));
  NAND3_X1  g698(.A1(new_n896_), .A2(new_n204_), .A3(new_n592_), .ZN(new_n900_));
  OAI21_X1  g699(.A(G148gat), .B1(new_n895_), .B2(new_n593_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1345gat));
  XNOR2_X1  g701(.A(KEYINPUT61), .B(G155gat), .ZN(new_n903_));
  OR3_X1    g702(.A1(new_n895_), .A2(new_n621_), .A3(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n895_), .B2(new_n621_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1346gat));
  OR3_X1    g705(.A1(new_n895_), .A2(G162gat), .A3(new_n518_), .ZN(new_n907_));
  OAI21_X1  g706(.A(G162gat), .B1(new_n895_), .B2(new_n618_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n907_), .A2(new_n908_), .ZN(G1347gat));
  NOR2_X1   g708(.A1(new_n447_), .A2(new_n451_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(new_n626_), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n448_), .B(new_n911_), .C1(new_n847_), .C2(new_n797_), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n267_), .B1(new_n912_), .B2(new_n555_), .ZN(new_n913_));
  OR2_X1    g712(.A1(new_n913_), .A2(KEYINPUT62), .ZN(new_n914_));
  NAND3_X1  g713(.A1(new_n912_), .A2(new_n301_), .A3(new_n555_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n913_), .A2(KEYINPUT62), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(G1348gat));
  AND2_X1   g716(.A1(new_n859_), .A2(new_n797_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n448_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n911_), .A2(new_n268_), .A3(new_n593_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n912_), .A2(new_n592_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n919_), .A2(new_n920_), .B1(new_n300_), .B2(new_n921_), .ZN(G1349gat));
  NAND2_X1  g721(.A1(new_n328_), .A2(new_n329_), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n912_), .A2(new_n923_), .A3(new_n610_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n911_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n919_), .A2(new_n620_), .A3(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(new_n303_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n924_), .B1(new_n926_), .B2(new_n927_), .ZN(G1350gat));
  NAND3_X1  g727(.A1(new_n912_), .A2(new_n289_), .A3(new_n798_), .ZN(new_n929_));
  AND2_X1   g728(.A1(new_n912_), .A2(new_n619_), .ZN(new_n930_));
  INV_X1    g729(.A(G190gat), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n929_), .B1(new_n930_), .B2(new_n931_), .ZN(G1351gat));
  NOR4_X1   g731(.A1(new_n445_), .A2(new_n258_), .A3(new_n394_), .A4(new_n451_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n918_), .A2(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(G197gat), .B1(new_n935_), .B2(new_n555_), .ZN(new_n936_));
  NOR4_X1   g735(.A1(new_n918_), .A2(new_n312_), .A3(new_n554_), .A4(new_n934_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n936_), .A2(new_n937_), .ZN(G1352gat));
  NAND2_X1  g737(.A1(new_n309_), .A2(new_n311_), .ZN(new_n939_));
  AND4_X1   g738(.A1(new_n939_), .A2(new_n873_), .A3(new_n592_), .A4(new_n933_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n935_), .A2(new_n592_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n941_), .B2(new_n308_), .ZN(G1353gat));
  XNOR2_X1  g741(.A(KEYINPUT63), .B(G211gat), .ZN(new_n943_));
  NOR4_X1   g742(.A1(new_n918_), .A2(new_n856_), .A3(new_n934_), .A4(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n935_), .A2(new_n610_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n944_), .B1(new_n945_), .B2(new_n946_), .ZN(G1354gat));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948_));
  NAND4_X1  g747(.A1(new_n873_), .A2(new_n948_), .A3(new_n798_), .A4(new_n933_), .ZN(new_n949_));
  INV_X1    g748(.A(G218gat), .ZN(new_n950_));
  AND2_X1   g749(.A1(new_n949_), .A2(new_n950_), .ZN(new_n951_));
  NAND3_X1  g750(.A1(new_n873_), .A2(new_n798_), .A3(new_n933_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n952_), .A2(KEYINPUT127), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n618_), .A2(new_n950_), .ZN(new_n954_));
  AOI22_X1  g753(.A1(new_n951_), .A2(new_n953_), .B1(new_n935_), .B2(new_n954_), .ZN(G1355gat));
endmodule


