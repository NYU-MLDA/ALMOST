//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 0 0 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n609_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n615_, new_n616_, new_n617_, new_n618_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n786_, new_n787_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n799_, new_n801_, new_n802_, new_n803_, new_n804_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n853_, new_n854_, new_n855_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(G141gat), .ZN(new_n203_));
  INV_X1    g002(.A(G148gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(KEYINPUT83), .A2(KEYINPUT3), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT85), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n208_), .B1(new_n209_), .B2(KEYINPUT84), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT2), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n212_), .B1(new_n209_), .B2(new_n208_), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n207_), .B(new_n211_), .C1(new_n213_), .C2(new_n210_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215_));
  OR2_X1    g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n214_), .A2(new_n215_), .A3(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(new_n215_), .A2(KEYINPUT1), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(KEYINPUT1), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(new_n216_), .A3(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(new_n205_), .A3(new_n209_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(G127gat), .B(G134gat), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G113gat), .B(G120gat), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n222_), .B(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT4), .ZN(new_n227_));
  INV_X1    g026(.A(new_n222_), .ZN(new_n228_));
  OR3_X1    g027(.A1(new_n228_), .A2(KEYINPUT4), .A3(new_n225_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n202_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(G57gat), .B(G85gat), .Z(new_n231_));
  XNOR2_X1  g030(.A(G1gat), .B(G29gat), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n202_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n226_), .A2(new_n236_), .ZN(new_n237_));
  OR3_X1    g036(.A1(new_n230_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n235_), .B1(new_n230_), .B2(new_n237_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n241_), .A2(G1gat), .ZN(new_n242_));
  INV_X1    g041(.A(G204gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(G197gat), .ZN(new_n244_));
  INV_X1    g043(.A(G197gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G204gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n244_), .A2(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(G211gat), .A2(G218gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G211gat), .A2(G218gat), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n247_), .A2(KEYINPUT21), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  AND2_X1   g049(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n251_));
  NOR2_X1   g050(.A1(KEYINPUT86), .A2(KEYINPUT21), .ZN(new_n252_));
  OAI211_X1 g051(.A(new_n244_), .B(new_n246_), .C1(new_n251_), .C2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT87), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT86), .B(KEYINPUT21), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n256_), .A2(KEYINPUT87), .A3(new_n244_), .A4(new_n246_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n250_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n247_), .A2(KEYINPUT21), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n248_), .A2(new_n249_), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT88), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n258_), .A2(new_n261_), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n250_), .A2(new_n255_), .A3(new_n257_), .A4(KEYINPUT88), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n265_), .B1(KEYINPUT29), .B2(new_n222_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G228gat), .A2(G233gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(G78gat), .B(G106gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n268_), .B(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT89), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n222_), .A2(KEYINPUT29), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT28), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G22gat), .B(G50gat), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n273_), .A2(new_n274_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n271_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n270_), .A2(new_n277_), .ZN(new_n278_));
  OR3_X1    g077(.A1(new_n275_), .A2(new_n276_), .A3(new_n271_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n279_), .A2(new_n277_), .A3(new_n270_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n278_), .A2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n283_));
  AND2_X1   g082(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n284_));
  AND2_X1   g083(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n285_));
  NOR2_X1   g084(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n286_));
  OAI22_X1  g085(.A1(new_n283_), .A2(new_n284_), .B1(new_n285_), .B2(new_n286_), .ZN(new_n287_));
  OR3_X1    g086(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n288_));
  INV_X1    g087(.A(G169gat), .ZN(new_n289_));
  INV_X1    g088(.A(G176gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G169gat), .A2(G176gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(KEYINPUT24), .A3(new_n292_), .ZN(new_n293_));
  AND3_X1   g092(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n287_), .A2(new_n288_), .A3(new_n293_), .A4(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G183gat), .A2(G190gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT23), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OR2_X1    g099(.A1(G183gat), .A2(G190gat), .ZN(new_n301_));
  NAND3_X1  g100(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  AND2_X1   g102(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n304_));
  NOR2_X1   g103(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n305_));
  OAI21_X1  g104(.A(new_n290_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n303_), .A2(new_n306_), .A3(new_n292_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n297_), .A2(new_n307_), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n262_), .A2(new_n263_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n309_), .A2(KEYINPUT20), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT90), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT91), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n292_), .A2(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n306_), .A2(new_n292_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n314_), .B(new_n303_), .C1(new_n315_), .C2(new_n313_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(new_n297_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n264_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n309_), .A2(KEYINPUT90), .A3(KEYINPUT20), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n312_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G226gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT19), .ZN(new_n322_));
  INV_X1    g121(.A(new_n317_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n265_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT20), .ZN(new_n325_));
  INV_X1    g124(.A(new_n308_), .ZN(new_n326_));
  AOI211_X1 g125(.A(new_n325_), .B(new_n322_), .C1(new_n264_), .C2(new_n326_), .ZN(new_n327_));
  AOI22_X1  g126(.A1(new_n320_), .A2(new_n322_), .B1(new_n324_), .B2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G8gat), .B(G36gat), .ZN(new_n329_));
  INV_X1    g128(.A(G92gat), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT18), .B(G64gat), .ZN(new_n332_));
  XOR2_X1   g131(.A(new_n331_), .B(new_n332_), .Z(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT92), .B1(new_n328_), .B2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n320_), .A2(new_n322_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n327_), .A2(new_n324_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n336_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT92), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n328_), .A2(new_n340_), .A3(new_n334_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  OR3_X1    g141(.A1(new_n339_), .A2(KEYINPUT27), .A3(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n264_), .B1(new_n323_), .B2(KEYINPUT98), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(KEYINPUT98), .B2(new_n323_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n345_), .B(KEYINPUT20), .C1(new_n265_), .C2(new_n308_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(new_n322_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n347_), .B1(new_n322_), .B2(new_n320_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(new_n333_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n336_), .A2(new_n334_), .A3(new_n337_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(KEYINPUT27), .A3(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n343_), .A2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n282_), .A2(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n225_), .B(G71gat), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G227gat), .A2(G233gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n354_), .B(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n357_));
  XOR2_X1   g156(.A(new_n357_), .B(KEYINPUT31), .Z(new_n358_));
  XNOR2_X1  g157(.A(new_n356_), .B(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G15gat), .B(G43gat), .ZN(new_n360_));
  INV_X1    g159(.A(G99gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n308_), .B(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n359_), .B(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n353_), .A2(new_n241_), .A3(new_n364_), .ZN(new_n365_));
  AND2_X1   g164(.A1(new_n226_), .A2(new_n236_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT95), .B1(new_n366_), .B2(new_n235_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n227_), .A2(new_n202_), .A3(new_n229_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n235_), .B1(new_n226_), .B2(new_n236_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT95), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n367_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT96), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT96), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n367_), .A2(new_n374_), .A3(new_n368_), .A4(new_n371_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n373_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n239_), .A2(KEYINPUT33), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT33), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n378_), .B(new_n235_), .C1(new_n230_), .C2(new_n237_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n309_), .A2(KEYINPUT90), .A3(KEYINPUT20), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT90), .B1(new_n309_), .B2(KEYINPUT20), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n264_), .A2(new_n317_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n381_), .A2(new_n382_), .A3(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n322_), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n337_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(new_n333_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n387_), .A2(KEYINPUT92), .A3(new_n350_), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n388_), .A2(KEYINPUT93), .A3(new_n341_), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT93), .B1(new_n388_), .B2(new_n341_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n376_), .B(new_n380_), .C1(new_n389_), .C2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT97), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n334_), .A2(KEYINPUT32), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n348_), .A2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n240_), .B(new_n394_), .C1(new_n393_), .C2(new_n386_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT93), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n396_), .B1(new_n339_), .B2(new_n342_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n388_), .A2(KEYINPUT93), .A3(new_n341_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT97), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n376_), .A4(new_n380_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n392_), .A2(new_n395_), .A3(new_n401_), .ZN(new_n402_));
  AND3_X1   g201(.A1(new_n402_), .A2(KEYINPUT99), .A3(new_n281_), .ZN(new_n403_));
  AOI21_X1  g202(.A(KEYINPUT99), .B1(new_n402_), .B2(new_n281_), .ZN(new_n404_));
  NOR3_X1   g203(.A1(new_n352_), .A2(new_n240_), .A3(new_n281_), .ZN(new_n405_));
  NOR3_X1   g204(.A1(new_n403_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n364_), .B(KEYINPUT82), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n365_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT100), .ZN(new_n409_));
  XOR2_X1   g208(.A(G29gat), .B(G36gat), .Z(new_n410_));
  XNOR2_X1  g209(.A(G43gat), .B(G50gat), .ZN(new_n411_));
  OR2_X1    g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n411_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT15), .ZN(new_n415_));
  XNOR2_X1  g214(.A(G15gat), .B(G22gat), .ZN(new_n416_));
  INV_X1    g215(.A(G1gat), .ZN(new_n417_));
  INV_X1    g216(.A(G8gat), .ZN(new_n418_));
  OAI21_X1  g217(.A(KEYINPUT14), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(G1gat), .B(G8gat), .ZN(new_n421_));
  XNOR2_X1  g220(.A(new_n420_), .B(new_n421_), .ZN(new_n422_));
  MUX2_X1   g221(.A(new_n414_), .B(new_n415_), .S(new_n422_), .Z(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n414_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT80), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G229gat), .A2(G233gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  MUX2_X1   g226(.A(new_n423_), .B(new_n425_), .S(new_n427_), .Z(new_n428_));
  XNOR2_X1  g227(.A(G113gat), .B(G141gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G169gat), .B(G197gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n429_), .B(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n428_), .B(new_n431_), .Z(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n408_), .A2(new_n409_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n365_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n402_), .A2(new_n281_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT99), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n402_), .A2(KEYINPUT99), .A3(new_n281_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n405_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n407_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n435_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT100), .B1(new_n443_), .B2(new_n432_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n434_), .A2(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(G85gat), .B(G92gat), .Z(new_n446_));
  NAND2_X1  g245(.A1(G99gat), .A2(G106gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT6), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT65), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT7), .ZN(new_n450_));
  INV_X1    g249(.A(G106gat), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n450_), .A2(new_n361_), .A3(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT66), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n446_), .B1(new_n449_), .B2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT8), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT67), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n456_), .A2(KEYINPUT67), .A3(KEYINPUT8), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT8), .ZN(new_n461_));
  INV_X1    g260(.A(new_n448_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n461_), .B(new_n446_), .C1(new_n462_), .C2(new_n454_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n459_), .A2(new_n460_), .A3(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n446_), .A2(KEYINPUT9), .ZN(new_n465_));
  XOR2_X1   g264(.A(KEYINPUT10), .B(G99gat), .Z(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n451_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT64), .ZN(new_n468_));
  NOR3_X1   g267(.A1(new_n468_), .A2(new_n330_), .A3(KEYINPUT9), .ZN(new_n469_));
  NOR2_X1   g268(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n470_));
  OAI21_X1  g269(.A(G85gat), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n465_), .A2(new_n467_), .A3(new_n471_), .A4(new_n448_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n464_), .A2(new_n472_), .ZN(new_n473_));
  XOR2_X1   g272(.A(G57gat), .B(G64gat), .Z(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT11), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT11), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G71gat), .B(G78gat), .ZN(new_n478_));
  MUX2_X1   g277(.A(new_n475_), .B(new_n477_), .S(new_n478_), .Z(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n473_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT12), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n482_), .A2(KEYINPUT68), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G230gat), .A2(G233gat), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n482_), .A2(KEYINPUT68), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n473_), .A2(new_n480_), .A3(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n486_), .B1(new_n473_), .B2(new_n480_), .ZN(new_n488_));
  OAI211_X1 g287(.A(new_n484_), .B(new_n485_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n464_), .A2(new_n472_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n490_), .A2(new_n479_), .ZN(new_n491_));
  OAI211_X1 g290(.A(G230gat), .B(G233gat), .C1(new_n491_), .C2(new_n481_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n489_), .A2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(KEYINPUT69), .B(KEYINPUT5), .Z(new_n494_));
  XNOR2_X1  g293(.A(G120gat), .B(G148gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G176gat), .B(G204gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n496_), .B(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n493_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n489_), .A2(new_n492_), .A3(new_n498_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(KEYINPUT70), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(KEYINPUT70), .B1(new_n500_), .B2(new_n501_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT13), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n504_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT13), .ZN(new_n507_));
  NAND3_X1  g306(.A1(new_n506_), .A2(new_n502_), .A3(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(KEYINPUT71), .B1(new_n505_), .B2(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n505_), .A2(new_n508_), .A3(KEYINPUT71), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(new_n511_), .A3(KEYINPUT72), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT72), .ZN(new_n513_));
  INV_X1    g312(.A(new_n511_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n513_), .B1(new_n514_), .B2(new_n509_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G231gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n422_), .B(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n480_), .B(new_n517_), .ZN(new_n518_));
  XOR2_X1   g317(.A(G127gat), .B(G155gat), .Z(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(G211gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(KEYINPUT16), .B(G183gat), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n520_), .B(new_n521_), .Z(new_n522_));
  AND2_X1   g321(.A1(new_n522_), .A2(KEYINPUT17), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n518_), .A2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n524_), .B(KEYINPUT78), .Z(new_n525_));
  NOR2_X1   g324(.A1(new_n518_), .A2(new_n523_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n526_), .B1(KEYINPUT17), .B2(new_n522_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n525_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G232gat), .A2(G233gat), .ZN(new_n529_));
  XOR2_X1   g328(.A(new_n529_), .B(KEYINPUT34), .Z(new_n530_));
  NAND4_X1  g329(.A1(new_n464_), .A2(new_n413_), .A3(new_n412_), .A4(new_n472_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n531_), .B1(new_n490_), .B2(new_n415_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n530_), .B1(new_n532_), .B2(KEYINPUT35), .ZN(new_n533_));
  OR2_X1    g332(.A1(new_n530_), .A2(KEYINPUT35), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n532_), .A2(KEYINPUT73), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n536_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n538_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n537_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G134gat), .B(G162gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(G218gat), .ZN(new_n542_));
  XOR2_X1   g341(.A(KEYINPUT74), .B(G190gat), .Z(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT36), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT75), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n540_), .A2(KEYINPUT76), .A3(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n537_), .A2(new_n539_), .A3(new_n545_), .A4(new_n544_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  AOI21_X1  g350(.A(KEYINPUT76), .B1(new_n540_), .B2(new_n548_), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT37), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n540_), .A2(KEYINPUT77), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT77), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n537_), .A2(new_n555_), .A3(new_n539_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(new_n556_), .A3(new_n548_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT37), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(new_n550_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n528_), .B1(new_n553_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT79), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  AOI211_X1 g361(.A(KEYINPUT79), .B(new_n528_), .C1(new_n553_), .C2(new_n559_), .ZN(new_n563_));
  OAI211_X1 g362(.A(new_n512_), .B(new_n515_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  AOI21_X1  g364(.A(KEYINPUT101), .B1(new_n445_), .B2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT101), .ZN(new_n567_));
  AOI211_X1 g366(.A(new_n567_), .B(new_n564_), .C1(new_n434_), .C2(new_n444_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT102), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n566_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n409_), .B1(new_n408_), .B2(new_n433_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n443_), .A2(KEYINPUT100), .A3(new_n432_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n565_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n567_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n445_), .A2(KEYINPUT101), .A3(new_n565_), .ZN(new_n575_));
  AOI21_X1  g374(.A(KEYINPUT102), .B1(new_n574_), .B2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n242_), .B1(new_n570_), .B2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT103), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n569_), .B1(new_n566_), .B2(new_n568_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n574_), .A2(KEYINPUT102), .A3(new_n575_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n582_), .A2(KEYINPUT103), .A3(new_n242_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n579_), .A2(KEYINPUT38), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT104), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n579_), .A2(new_n583_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT38), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n510_), .A2(new_n511_), .A3(new_n433_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT105), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n557_), .A2(new_n550_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n592_), .A2(new_n528_), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n591_), .A2(new_n408_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  OAI21_X1  g394(.A(G1gat), .B1(new_n595_), .B2(new_n241_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n579_), .A2(KEYINPUT104), .A3(KEYINPUT38), .A4(new_n583_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n586_), .A2(new_n589_), .A3(new_n596_), .A4(new_n597_), .ZN(G1324gat));
  AOI21_X1  g397(.A(new_n418_), .B1(new_n594_), .B2(new_n352_), .ZN(new_n599_));
  XOR2_X1   g398(.A(new_n599_), .B(KEYINPUT39), .Z(new_n600_));
  AND4_X1   g399(.A1(KEYINPUT106), .A2(new_n582_), .A3(new_n418_), .A4(new_n352_), .ZN(new_n601_));
  AOI21_X1  g400(.A(G8gat), .B1(new_n580_), .B2(new_n581_), .ZN(new_n602_));
  AOI21_X1  g401(.A(KEYINPUT106), .B1(new_n602_), .B2(new_n352_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n600_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT40), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  OAI211_X1 g405(.A(KEYINPUT40), .B(new_n600_), .C1(new_n601_), .C2(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(G1325gat));
  INV_X1    g407(.A(G15gat), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n609_), .B1(new_n594_), .B2(new_n407_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT41), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n566_), .A2(new_n568_), .ZN(new_n612_));
  NAND3_X1  g411(.A1(new_n612_), .A2(new_n609_), .A3(new_n407_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(G1326gat));
  INV_X1    g413(.A(G22gat), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n615_), .B1(new_n594_), .B2(new_n282_), .ZN(new_n616_));
  XOR2_X1   g415(.A(new_n616_), .B(KEYINPUT42), .Z(new_n617_));
  NAND3_X1  g416(.A1(new_n612_), .A2(new_n615_), .A3(new_n282_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(G1327gat));
  NOR2_X1   g418(.A1(new_n514_), .A2(new_n509_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n592_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n528_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AND3_X1   g422(.A1(new_n445_), .A2(new_n620_), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(G29gat), .B1(new_n624_), .B2(new_n240_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT43), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n553_), .A2(new_n559_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n626_), .B1(new_n443_), .B2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n627_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n408_), .A2(KEYINPUT43), .A3(new_n629_), .ZN(new_n630_));
  NAND4_X1  g429(.A1(new_n591_), .A2(new_n528_), .A3(new_n628_), .A4(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT44), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(G29gat), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n631_), .A2(new_n632_), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n635_), .A2(new_n241_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n625_), .B1(new_n634_), .B2(new_n636_), .ZN(G1328gat));
  INV_X1    g436(.A(G36gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n624_), .A2(new_n638_), .A3(new_n352_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n639_), .B(KEYINPUT45), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n633_), .A2(new_n352_), .ZN(new_n641_));
  OAI21_X1  g440(.A(G36gat), .B1(new_n641_), .B2(new_n635_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT46), .Z(G1329gat));
  INV_X1    g443(.A(G43gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n645_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n646_));
  OAI211_X1 g445(.A(new_n646_), .B(new_n364_), .C1(new_n632_), .C2(new_n631_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT107), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n647_), .A2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n647_), .A2(new_n648_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n624_), .A2(new_n407_), .ZN(new_n651_));
  OAI22_X1  g450(.A1(new_n649_), .A2(new_n650_), .B1(G43gat), .B2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g452(.A(G50gat), .B1(new_n624_), .B2(new_n282_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n633_), .A2(G50gat), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n635_), .A2(new_n281_), .ZN(new_n656_));
  AOI21_X1  g455(.A(new_n654_), .B1(new_n655_), .B2(new_n656_), .ZN(G1331gat));
  NOR2_X1   g456(.A1(new_n443_), .A2(new_n433_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n562_), .A2(new_n563_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(new_n620_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n658_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(G57gat), .B1(new_n663_), .B2(new_n240_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n512_), .A2(new_n515_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n658_), .A2(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n593_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n667_), .A2(new_n241_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n664_), .B1(new_n668_), .B2(G57gat), .ZN(G1332gat));
  INV_X1    g468(.A(new_n352_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G64gat), .B1(new_n667_), .B2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT48), .ZN(new_n672_));
  OR2_X1    g471(.A1(new_n670_), .A2(G64gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n662_), .B2(new_n673_), .ZN(G1333gat));
  OAI21_X1  g473(.A(G71gat), .B1(new_n667_), .B2(new_n442_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT49), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n442_), .A2(G71gat), .ZN(new_n677_));
  XOR2_X1   g476(.A(new_n677_), .B(KEYINPUT108), .Z(new_n678_));
  OAI21_X1  g477(.A(new_n676_), .B1(new_n662_), .B2(new_n678_), .ZN(G1334gat));
  OAI21_X1  g478(.A(G78gat), .B1(new_n667_), .B2(new_n281_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT50), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n662_), .A2(G78gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n681_), .B1(new_n281_), .B2(new_n682_), .ZN(G1335gat));
  AND2_X1   g482(.A1(new_n666_), .A2(new_n623_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G85gat), .B1(new_n684_), .B2(new_n240_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n630_), .A2(new_n628_), .ZN(new_n686_));
  NAND4_X1  g485(.A1(new_n686_), .A2(new_n432_), .A3(new_n528_), .A4(new_n661_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n687_), .A2(new_n241_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n685_), .B1(new_n688_), .B2(G85gat), .ZN(G1336gat));
  AOI21_X1  g488(.A(G92gat), .B1(new_n684_), .B2(new_n352_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n687_), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n468_), .A2(new_n330_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n352_), .B1(new_n470_), .B2(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT109), .Z(new_n694_));
  AOI21_X1  g493(.A(new_n690_), .B1(new_n691_), .B2(new_n694_), .ZN(G1337gat));
  OAI21_X1  g494(.A(G99gat), .B1(new_n687_), .B2(new_n442_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n684_), .A2(new_n364_), .A3(new_n466_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n698_), .B(new_n699_), .ZN(G1338gat));
  OAI21_X1  g499(.A(G106gat), .B1(new_n687_), .B2(new_n281_), .ZN(new_n701_));
  XOR2_X1   g500(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  OR2_X1    g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n684_), .A2(new_n451_), .A3(new_n282_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n701_), .A2(new_n703_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n704_), .A2(new_n705_), .A3(new_n706_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g507(.A(KEYINPUT117), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT55), .ZN(new_n710_));
  OR3_X1    g509(.A1(new_n489_), .A2(KEYINPUT113), .A3(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n484_), .B1(new_n488_), .B2(new_n487_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT112), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT112), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n484_), .B(new_n714_), .C1(new_n487_), .C2(new_n488_), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n713_), .A2(G230gat), .A3(G233gat), .A4(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n489_), .A2(new_n710_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT113), .B1(new_n489_), .B2(new_n710_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n711_), .A2(new_n716_), .A3(new_n717_), .A4(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n499_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT56), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n428_), .A2(new_n431_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n425_), .A2(new_n426_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n431_), .ZN(new_n725_));
  XOR2_X1   g524(.A(new_n725_), .B(KEYINPUT114), .Z(new_n726_));
  NAND2_X1  g525(.A1(new_n423_), .A2(new_n427_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n723_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n722_), .A2(new_n501_), .A3(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT58), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n722_), .A2(KEYINPUT58), .A3(new_n501_), .A4(new_n728_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n629_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT115), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT57), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n433_), .A2(new_n501_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n720_), .A2(new_n721_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT56), .B1(new_n719_), .B2(new_n499_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n736_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n506_), .A2(new_n502_), .A3(new_n728_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  OAI211_X1 g540(.A(new_n734_), .B(new_n735_), .C1(new_n741_), .C2(new_n592_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n592_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n743_));
  OAI21_X1  g542(.A(KEYINPUT57), .B1(new_n743_), .B2(KEYINPUT115), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n733_), .A2(new_n742_), .A3(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n528_), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n505_), .A2(new_n508_), .A3(new_n432_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n560_), .A2(new_n747_), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(KEYINPUT54), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(KEYINPUT54), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n746_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT116), .ZN(new_n754_));
  AOI21_X1  g553(.A(KEYINPUT59), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n240_), .A2(new_n364_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n753_), .A2(new_n353_), .A3(new_n757_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n755_), .A2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n751_), .B1(new_n745_), .B2(new_n528_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n353_), .ZN(new_n761_));
  NOR3_X1   g560(.A1(new_n760_), .A2(new_n761_), .A3(new_n756_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT59), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n763_), .B1(new_n760_), .B2(KEYINPUT116), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n762_), .A2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n433_), .B1(new_n759_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(G113gat), .ZN(new_n767_));
  INV_X1    g566(.A(G113gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n762_), .A2(new_n768_), .A3(new_n433_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n709_), .B1(new_n767_), .B2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n755_), .A2(new_n758_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n762_), .A2(new_n764_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n432_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n709_), .B(new_n769_), .C1(new_n773_), .C2(new_n768_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n770_), .A2(new_n775_), .ZN(G1340gat));
  INV_X1    g575(.A(G120gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n620_), .B2(KEYINPUT60), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT118), .ZN(new_n779_));
  OAI211_X1 g578(.A(new_n762_), .B(new_n779_), .C1(KEYINPUT60), .C2(new_n777_), .ZN(new_n780_));
  XOR2_X1   g579(.A(new_n780_), .B(KEYINPUT119), .Z(new_n781_));
  NOR2_X1   g580(.A1(new_n759_), .A2(new_n765_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n665_), .ZN(new_n783_));
  OAI21_X1  g582(.A(G120gat), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n781_), .A2(new_n784_), .ZN(G1341gat));
  AOI21_X1  g584(.A(G127gat), .B1(new_n762_), .B2(new_n622_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n782_), .A2(new_n528_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g587(.A(G134gat), .B1(new_n762_), .B2(new_n592_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n782_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n629_), .A2(G134gat), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT120), .Z(new_n792_));
  AOI21_X1  g591(.A(new_n789_), .B1(new_n790_), .B2(new_n792_), .ZN(G1343gat));
  NOR3_X1   g592(.A1(new_n760_), .A2(new_n241_), .A3(new_n352_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n407_), .A2(new_n281_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n796_), .A2(new_n432_), .ZN(new_n797_));
  XNOR2_X1  g596(.A(new_n797_), .B(new_n203_), .ZN(G1344gat));
  NOR2_X1   g597(.A1(new_n796_), .A2(new_n783_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(new_n204_), .ZN(G1345gat));
  OR3_X1    g599(.A1(new_n796_), .A2(KEYINPUT121), .A3(new_n528_), .ZN(new_n801_));
  OAI21_X1  g600(.A(KEYINPUT121), .B1(new_n796_), .B2(new_n528_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(KEYINPUT61), .B(G155gat), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n803_), .B(new_n804_), .ZN(G1346gat));
  INV_X1    g604(.A(new_n796_), .ZN(new_n806_));
  AOI21_X1  g605(.A(G162gat), .B1(new_n806_), .B2(new_n592_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n629_), .A2(G162gat), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT122), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n807_), .B1(new_n806_), .B2(new_n809_), .ZN(G1347gat));
  NOR3_X1   g609(.A1(new_n760_), .A2(new_n240_), .A3(new_n670_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(new_n281_), .A3(new_n407_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n812_), .A2(new_n432_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n813_), .A2(new_n289_), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n814_), .A2(KEYINPUT62), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n813_), .B1(new_n305_), .B2(new_n304_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n814_), .A2(KEYINPUT62), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n816_), .A3(new_n817_), .ZN(G1348gat));
  AND3_X1   g617(.A1(new_n811_), .A2(new_n281_), .A3(new_n407_), .ZN(new_n819_));
  AOI21_X1  g618(.A(G176gat), .B1(new_n819_), .B2(new_n661_), .ZN(new_n820_));
  NOR3_X1   g619(.A1(new_n812_), .A2(new_n290_), .A3(new_n783_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1349gat));
  INV_X1    g621(.A(new_n284_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT123), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n283_), .A2(new_n824_), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n819_), .A2(new_n823_), .A3(new_n622_), .A4(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(G183gat), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n824_), .B(new_n827_), .C1(new_n812_), .C2(new_n528_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT124), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(G1350gat));
  OAI21_X1  g630(.A(G190gat), .B1(new_n812_), .B2(new_n627_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n819_), .B1(new_n286_), .B2(new_n285_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n832_), .B1(new_n833_), .B2(new_n621_), .ZN(G1351gat));
  NAND2_X1  g633(.A1(new_n811_), .A2(new_n795_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n432_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n836_), .B(new_n245_), .ZN(G1352gat));
  NOR2_X1   g636(.A1(new_n835_), .A2(new_n783_), .ZN(new_n838_));
  XNOR2_X1  g637(.A(new_n838_), .B(new_n243_), .ZN(G1353gat));
  AND2_X1   g638(.A1(new_n811_), .A2(new_n795_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n528_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n840_), .B1(KEYINPUT125), .B2(new_n842_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n842_), .A2(KEYINPUT125), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT126), .ZN(new_n846_));
  NOR2_X1   g645(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n846_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n850_));
  OAI211_X1 g649(.A(new_n849_), .B(new_n850_), .C1(new_n843_), .C2(new_n844_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n848_), .A2(new_n851_), .ZN(G1354gat));
  NAND3_X1  g651(.A1(new_n840_), .A2(G218gat), .A3(new_n629_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n835_), .A2(new_n621_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(G218gat), .B2(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


