//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n829_, new_n830_, new_n831_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n840_, new_n841_, new_n843_, new_n844_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n872_, new_n873_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(G113gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(G127gat), .A2(G134gat), .ZN(new_n204_));
  INV_X1    g003(.A(G113gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G127gat), .A2(G134gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  AND3_X1   g006(.A1(new_n203_), .A2(G120gat), .A3(new_n207_), .ZN(new_n208_));
  AOI21_X1  g007(.A(G120gat), .B1(new_n203_), .B2(new_n207_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  NOR2_X1   g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT2), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n218_));
  NAND4_X1  g017(.A1(new_n213_), .A2(new_n216_), .A3(new_n217_), .A4(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT82), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  AND2_X1   g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT83), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G155gat), .ZN(new_n225_));
  INV_X1    g024(.A(G162gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT83), .ZN(new_n228_));
  NAND2_X1  g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  AND2_X1   g029(.A1(new_n224_), .A2(new_n230_), .ZN(new_n231_));
  AND3_X1   g030(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n234_), .A2(KEYINPUT82), .A3(new_n217_), .A4(new_n213_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n221_), .A2(new_n231_), .A3(new_n235_), .ZN(new_n236_));
  AOI22_X1  g035(.A1(new_n222_), .A2(KEYINPUT1), .B1(G141gat), .B2(G148gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n227_), .A2(new_n229_), .ZN(new_n238_));
  OAI221_X1 g037(.A(new_n237_), .B1(G141gat), .B2(G148gat), .C1(KEYINPUT1), .C2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n236_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n210_), .A2(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n208_), .A2(new_n209_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(new_n239_), .A3(new_n236_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n241_), .A2(KEYINPUT95), .A3(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT95), .ZN(new_n245_));
  NAND4_X1  g044(.A1(new_n242_), .A2(new_n245_), .A3(new_n239_), .A4(new_n236_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(KEYINPUT4), .A3(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248_));
  XOR2_X1   g047(.A(new_n248_), .B(KEYINPUT96), .Z(new_n249_));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n241_), .A2(new_n250_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n247_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n249_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n244_), .A2(new_n253_), .A3(new_n246_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT0), .B(G57gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(G85gat), .ZN(new_n257_));
  XOR2_X1   g056(.A(G1gat), .B(G29gat), .Z(new_n258_));
  XOR2_X1   g057(.A(new_n257_), .B(new_n258_), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n255_), .B(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT88), .ZN(new_n263_));
  INV_X1    g062(.A(G204gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n263_), .B1(new_n264_), .B2(G197gat), .ZN(new_n265_));
  INV_X1    g064(.A(G197gat), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(KEYINPUT88), .A3(G204gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT87), .B(G204gat), .ZN(new_n268_));
  OAI211_X1 g067(.A(new_n265_), .B(new_n267_), .C1(new_n268_), .C2(new_n266_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G211gat), .B(G218gat), .Z(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(KEYINPUT21), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT89), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n270_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G197gat), .A2(G204gat), .ZN(new_n275_));
  OAI211_X1 g074(.A(KEYINPUT21), .B(new_n275_), .C1(new_n268_), .C2(G197gat), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n274_), .B(new_n276_), .C1(new_n269_), .C2(KEYINPUT21), .ZN(new_n277_));
  NAND4_X1  g076(.A1(new_n269_), .A2(KEYINPUT89), .A3(KEYINPUT21), .A4(new_n270_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n273_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  AND3_X1   g078(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G169gat), .ZN(new_n283_));
  INV_X1    g082(.A(G176gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(KEYINPUT24), .A3(new_n286_), .ZN(new_n287_));
  OR3_X1    g086(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n288_));
  AND3_X1   g087(.A1(new_n282_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT25), .B(G183gat), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT78), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n292_), .A2(new_n293_), .A3(KEYINPUT78), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n289_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  OR2_X1    g097(.A1(G183gat), .A2(G190gat), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n282_), .A2(new_n299_), .B1(G169gat), .B2(G176gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(G169gat), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n283_), .A2(KEYINPUT79), .A3(KEYINPUT22), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n302_), .A2(new_n303_), .A3(new_n284_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT80), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT80), .ZN(new_n306_));
  NAND4_X1  g105(.A1(new_n302_), .A2(new_n303_), .A3(new_n306_), .A4(new_n284_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n300_), .A2(new_n305_), .A3(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n298_), .A2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT20), .B1(new_n279_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT91), .ZN(new_n311_));
  AND3_X1   g110(.A1(new_n290_), .A2(KEYINPUT92), .A3(new_n291_), .ZN(new_n312_));
  AOI21_X1  g111(.A(KEYINPUT92), .B1(new_n290_), .B2(new_n291_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n293_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT22), .B(G169gat), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n284_), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n314_), .A2(new_n289_), .B1(new_n300_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n279_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT91), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n320_), .B(KEYINPUT20), .C1(new_n279_), .C2(new_n309_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n311_), .A2(new_n319_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(KEYINPUT19), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n324_), .ZN(new_n325_));
  XOR2_X1   g124(.A(G8gat), .B(G36gat), .Z(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT94), .B(KEYINPUT18), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G64gat), .B(G92gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n317_), .A2(new_n273_), .A3(new_n277_), .A4(new_n278_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT93), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT20), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n335_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n324_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n279_), .A2(new_n309_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n334_), .A2(new_n336_), .A3(new_n337_), .A4(new_n338_), .ZN(new_n339_));
  AND3_X1   g138(.A1(new_n325_), .A2(new_n331_), .A3(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n331_), .B1(new_n325_), .B2(new_n339_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n342_), .A2(KEYINPUT27), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n322_), .A2(new_n324_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n332_), .A2(KEYINPUT20), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n345_), .A2(KEYINPUT98), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n345_), .A2(KEYINPUT98), .B1(new_n309_), .B2(new_n279_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n337_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n330_), .B1(new_n344_), .B2(new_n348_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n325_), .A2(new_n331_), .A3(new_n339_), .ZN(new_n350_));
  AND3_X1   g149(.A1(new_n349_), .A2(KEYINPUT27), .A3(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n343_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n240_), .A2(KEYINPUT29), .ZN(new_n353_));
  AND2_X1   g152(.A1(new_n353_), .A2(new_n279_), .ZN(new_n354_));
  INV_X1    g153(.A(G233gat), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n355_), .A2(KEYINPUT86), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n355_), .A2(KEYINPUT86), .ZN(new_n357_));
  OAI21_X1  g156(.A(G228gat), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  OR2_X1    g157(.A1(new_n354_), .A2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n279_), .A2(new_n358_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT85), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n361_), .B1(new_n240_), .B2(KEYINPUT29), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n363_));
  AOI211_X1 g162(.A(KEYINPUT85), .B(new_n363_), .C1(new_n236_), .C2(new_n239_), .ZN(new_n364_));
  NOR4_X1   g163(.A1(new_n360_), .A2(new_n362_), .A3(new_n364_), .A4(KEYINPUT90), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT90), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n362_), .A2(new_n364_), .ZN(new_n367_));
  AND2_X1   g166(.A1(new_n279_), .A2(new_n358_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n359_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G78gat), .B(G106gat), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  OAI211_X1 g172(.A(new_n359_), .B(new_n371_), .C1(new_n365_), .C2(new_n369_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(KEYINPUT84), .A3(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n236_), .A2(new_n363_), .A3(new_n239_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G22gat), .B(G50gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n377_), .B(KEYINPUT28), .ZN(new_n378_));
  XOR2_X1   g177(.A(new_n376_), .B(new_n378_), .Z(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n375_), .A2(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(G71gat), .B(G99gat), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT30), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n298_), .A2(new_n308_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n384_), .B1(new_n298_), .B2(new_n308_), .ZN(new_n387_));
  OAI21_X1  g186(.A(G43gat), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n309_), .A2(KEYINPUT30), .ZN(new_n389_));
  INV_X1    g188(.A(G43gat), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n389_), .A2(new_n390_), .A3(new_n385_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G227gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(G15gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n388_), .A2(new_n391_), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n394_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n210_), .B(KEYINPUT31), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n398_), .A2(KEYINPUT81), .ZN(new_n399_));
  NOR3_X1   g198(.A1(new_n396_), .A2(new_n397_), .A3(new_n399_), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n398_), .A2(KEYINPUT81), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n388_), .A2(new_n391_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n394_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n401_), .B1(new_n404_), .B2(new_n395_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n383_), .B1(new_n400_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n399_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n404_), .A2(new_n401_), .A3(new_n395_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n382_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n406_), .A2(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n373_), .A2(KEYINPUT84), .A3(new_n374_), .A4(new_n379_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n381_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n410_), .B1(new_n381_), .B2(new_n411_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n262_), .B(new_n352_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n259_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT33), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(KEYINPUT97), .A3(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n249_), .B1(new_n247_), .B2(new_n251_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n253_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n420_));
  OR3_X1    g219(.A1(new_n419_), .A2(new_n260_), .A3(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT97), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT33), .B1(new_n415_), .B2(new_n422_), .ZN(new_n423_));
  NAND4_X1  g222(.A1(new_n342_), .A2(new_n418_), .A3(new_n421_), .A4(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n331_), .A2(KEYINPUT32), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(new_n426_), .B1(new_n344_), .B2(new_n348_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n325_), .A2(new_n425_), .A3(new_n339_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n255_), .A2(new_n260_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n427_), .B(new_n428_), .C1(new_n429_), .C2(new_n415_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(KEYINPUT99), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT99), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n261_), .A2(new_n432_), .A3(new_n428_), .A4(new_n427_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n424_), .A2(new_n431_), .A3(new_n433_), .ZN(new_n434_));
  AND2_X1   g233(.A1(new_n406_), .A2(new_n409_), .ZN(new_n435_));
  AND3_X1   g234(.A1(new_n435_), .A2(new_n411_), .A3(new_n381_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n434_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n414_), .A2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G29gat), .B(G36gat), .Z(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n390_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G29gat), .B(G36gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(G43gat), .ZN(new_n442_));
  AND3_X1   g241(.A1(new_n440_), .A2(G50gat), .A3(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(G50gat), .B1(new_n440_), .B2(new_n442_), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G15gat), .B(G22gat), .ZN(new_n446_));
  INV_X1    g245(.A(G1gat), .ZN(new_n447_));
  INV_X1    g246(.A(G8gat), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT14), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G1gat), .B(G8gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n450_), .B(new_n451_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n445_), .A2(new_n452_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n443_), .A2(new_n444_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT15), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT15), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n456_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(new_n453_), .B1(new_n458_), .B2(new_n452_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G229gat), .A2(G233gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n445_), .B(new_n452_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n460_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AND2_X1   g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G113gat), .B(G141gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(new_n283_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(new_n266_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT77), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n465_), .A2(KEYINPUT77), .A3(new_n469_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n468_), .B(KEYINPUT76), .ZN(new_n475_));
  OR2_X1    g274(.A1(new_n465_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n438_), .A2(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n478_), .B(KEYINPUT100), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G190gat), .B(G218gat), .ZN(new_n480_));
  XNOR2_X1  g279(.A(new_n480_), .B(G134gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n481_), .B(new_n226_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT36), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n483_), .A2(KEYINPUT36), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(KEYINPUT66), .A3(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT66), .ZN(new_n491_));
  INV_X1    g290(.A(new_n489_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n491_), .B1(new_n492_), .B2(new_n487_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT67), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT7), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n494_), .B(new_n495_), .C1(G99gat), .C2(G106gat), .ZN(new_n496_));
  INV_X1    g295(.A(G99gat), .ZN(new_n497_));
  INV_X1    g296(.A(G106gat), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n497_), .B(new_n498_), .C1(KEYINPUT67), .C2(KEYINPUT7), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n490_), .A2(new_n493_), .B1(new_n496_), .B2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G85gat), .B(G92gat), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT8), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n496_), .A2(new_n499_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n492_), .A2(new_n487_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n501_), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  OAI22_X1  g306(.A1(new_n500_), .A2(new_n504_), .B1(new_n507_), .B2(new_n503_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT70), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n490_), .A2(new_n493_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n511_));
  NOR2_X1   g310(.A1(new_n511_), .A2(KEYINPUT9), .ZN(new_n512_));
  NOR2_X1   g311(.A1(KEYINPUT65), .A2(G85gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(G92gat), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n502_), .A2(KEYINPUT9), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT10), .B(G99gat), .Z(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n498_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n510_), .A2(new_n514_), .A3(new_n515_), .A4(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n508_), .A2(new_n509_), .A3(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n509_), .B1(new_n508_), .B2(new_n518_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n458_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n454_), .A2(new_n508_), .A3(new_n518_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(G232gat), .A2(G233gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT34), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n525_), .A2(KEYINPUT35), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n522_), .A2(new_n523_), .A3(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(KEYINPUT35), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT72), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n508_), .A2(new_n518_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT70), .ZN(new_n533_));
  AOI22_X1  g332(.A1(new_n533_), .A2(new_n519_), .B1(new_n455_), .B2(new_n457_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n531_), .B1(new_n534_), .B2(KEYINPUT73), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n528_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT73), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n530_), .B1(new_n522_), .B2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n522_), .A2(new_n523_), .A3(new_n527_), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n484_), .B(new_n486_), .C1(new_n536_), .C2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n528_), .A2(new_n535_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n538_), .A2(new_n539_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n542_), .A2(new_n543_), .A3(new_n485_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n541_), .A2(KEYINPUT37), .A3(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n541_), .A2(KEYINPUT74), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n485_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT74), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n549_), .A3(new_n484_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n547_), .A2(new_n550_), .A3(new_n544_), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT37), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n546_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(KEYINPUT11), .ZN(new_n557_));
  XOR2_X1   g356(.A(G71gat), .B(G78gat), .Z(new_n558_));
  NAND3_X1  g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n557_), .A2(new_n558_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n561_), .B1(new_n508_), .B2(new_n518_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n562_), .A2(KEYINPUT12), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n533_), .A2(new_n519_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT71), .ZN(new_n565_));
  OAI21_X1  g364(.A(KEYINPUT12), .B1(new_n561_), .B2(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n566_), .B1(new_n565_), .B2(new_n561_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n563_), .B1(new_n564_), .B2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n508_), .A2(new_n561_), .A3(new_n518_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G230gat), .A2(G233gat), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n570_), .B(KEYINPUT64), .ZN(new_n571_));
  INV_X1    g370(.A(new_n571_), .ZN(new_n572_));
  AND2_X1   g371(.A1(new_n569_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n568_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G120gat), .B(G148gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(new_n264_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT5), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(new_n284_), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n569_), .B(KEYINPUT68), .Z(new_n579_));
  OR2_X1    g378(.A1(new_n579_), .A2(KEYINPUT69), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n562_), .B1(new_n579_), .B2(KEYINPUT69), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n574_), .B(new_n578_), .C1(new_n582_), .C2(new_n572_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT13), .ZN(new_n584_));
  INV_X1    g383(.A(new_n578_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n572_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n574_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  AND3_X1   g387(.A1(new_n583_), .A2(new_n584_), .A3(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n584_), .B1(new_n583_), .B2(new_n588_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(G231gat), .A2(G233gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT75), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n452_), .B(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(new_n561_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(KEYINPUT16), .B(G183gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(G211gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(G127gat), .B(G155gat), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n597_), .B(new_n598_), .Z(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n595_), .B1(KEYINPUT17), .B2(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n565_), .A3(KEYINPUT17), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n601_), .B(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n554_), .A2(new_n591_), .A3(new_n604_), .ZN(new_n605_));
  AND2_X1   g404(.A1(new_n479_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n447_), .A3(new_n261_), .ZN(new_n607_));
  INV_X1    g406(.A(KEYINPUT38), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n606_), .A2(KEYINPUT38), .A3(new_n447_), .A4(new_n261_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n551_), .B(KEYINPUT102), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n603_), .B(new_n477_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT101), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n611_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n612_), .A2(new_n613_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(new_n438_), .A3(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(G1gat), .B1(new_n617_), .B2(new_n262_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(KEYINPUT103), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n609_), .A2(new_n610_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT104), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(G1324gat));
  INV_X1    g421(.A(new_n352_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n615_), .A2(new_n623_), .A3(new_n438_), .A4(new_n616_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(G8gat), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT105), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n479_), .A2(new_n448_), .A3(new_n605_), .A4(new_n623_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n626_), .A2(new_n627_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(KEYINPUT105), .A2(KEYINPUT39), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n624_), .A2(G8gat), .A3(new_n630_), .A4(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n628_), .A2(new_n629_), .A3(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT106), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT106), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n628_), .A2(new_n629_), .A3(new_n635_), .A4(new_n632_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT40), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n637_), .B(new_n638_), .ZN(G1325gat));
  NAND3_X1  g438(.A1(new_n606_), .A2(new_n393_), .A3(new_n410_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G15gat), .B1(new_n617_), .B2(new_n435_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n641_), .A2(KEYINPUT107), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(KEYINPUT107), .ZN(new_n643_));
  AND3_X1   g442(.A1(new_n642_), .A2(KEYINPUT41), .A3(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(KEYINPUT41), .B1(new_n642_), .B2(new_n643_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n640_), .B1(new_n644_), .B2(new_n645_), .ZN(G1326gat));
  NAND2_X1  g445(.A1(new_n381_), .A2(new_n411_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  OAI21_X1  g447(.A(G22gat), .B1(new_n617_), .B2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT42), .ZN(new_n650_));
  INV_X1    g449(.A(G22gat), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n606_), .A2(new_n651_), .A3(new_n647_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(G1327gat));
  INV_X1    g452(.A(new_n591_), .ZN(new_n654_));
  NOR2_X1   g453(.A1(new_n611_), .A2(new_n603_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n479_), .A2(new_n654_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  AOI21_X1  g456(.A(G29gat), .B1(new_n657_), .B2(new_n261_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n438_), .A2(new_n554_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT43), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT43), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n438_), .A2(new_n661_), .A3(new_n554_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n477_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n591_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n663_), .A2(new_n604_), .A3(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND4_X1  g467(.A1(new_n663_), .A2(KEYINPUT44), .A3(new_n604_), .A4(new_n665_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(new_n262_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n658_), .B1(new_n671_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g471(.A(KEYINPUT45), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n352_), .A2(G36gat), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n673_), .B1(new_n656_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT100), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n478_), .B(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n678_), .A2(new_n591_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n679_), .A2(KEYINPUT45), .A3(new_n655_), .A4(new_n674_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n676_), .A2(new_n680_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G36gat), .B1(new_n670_), .B2(new_n352_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT46), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n681_), .A2(new_n682_), .A3(KEYINPUT46), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1329gat));
  AND4_X1   g486(.A1(G43gat), .A2(new_n668_), .A3(new_n410_), .A4(new_n669_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n657_), .A2(new_n410_), .ZN(new_n689_));
  XNOR2_X1  g488(.A(KEYINPUT108), .B(G43gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n688_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT47), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n689_), .A2(new_n690_), .ZN(new_n694_));
  OAI21_X1  g493(.A(KEYINPUT47), .B1(new_n694_), .B2(new_n688_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n693_), .A2(new_n695_), .ZN(G1330gat));
  OR3_X1    g495(.A1(new_n656_), .A2(G50gat), .A3(new_n648_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n668_), .A2(new_n647_), .A3(new_n669_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n698_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(KEYINPUT109), .B1(new_n698_), .B2(G50gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n697_), .B1(new_n699_), .B2(new_n700_), .ZN(G1331gat));
  INV_X1    g500(.A(G57gat), .ZN(new_n702_));
  AND3_X1   g501(.A1(new_n438_), .A2(new_n591_), .A3(new_n664_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n554_), .A2(new_n604_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n702_), .B1(new_n705_), .B2(new_n262_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT110), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n703_), .A2(new_n603_), .A3(new_n611_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(G57gat), .A3(new_n261_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n707_), .A2(new_n709_), .ZN(new_n710_));
  XOR2_X1   g509(.A(new_n710_), .B(KEYINPUT111), .Z(G1332gat));
  INV_X1    g510(.A(G64gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n708_), .B2(new_n623_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT48), .Z(new_n714_));
  INV_X1    g513(.A(new_n705_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n712_), .A3(new_n623_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1333gat));
  INV_X1    g516(.A(G71gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n708_), .B2(new_n410_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT49), .Z(new_n720_));
  NAND2_X1  g519(.A1(new_n410_), .A2(new_n718_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT112), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n705_), .B2(new_n722_), .ZN(G1334gat));
  INV_X1    g522(.A(G78gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n715_), .A2(new_n724_), .A3(new_n647_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT50), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n708_), .A2(new_n647_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(G78gat), .ZN(new_n728_));
  AOI211_X1 g527(.A(KEYINPUT50), .B(new_n724_), .C1(new_n708_), .C2(new_n647_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT113), .ZN(G1335gat));
  NAND2_X1  g530(.A1(new_n703_), .A2(new_n655_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n261_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n654_), .A2(new_n603_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n661_), .B1(new_n438_), .B2(new_n554_), .ZN(new_n736_));
  AOI211_X1 g535(.A(KEYINPUT43), .B(new_n553_), .C1(new_n414_), .C2(new_n437_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n664_), .B(new_n735_), .C1(new_n736_), .C2(new_n737_), .ZN(new_n738_));
  OR2_X1    g537(.A1(new_n738_), .A2(KEYINPUT114), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(KEYINPUT114), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n513_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n262_), .B1(new_n743_), .B2(new_n511_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n734_), .B1(new_n742_), .B2(new_n744_), .ZN(G1336gat));
  AOI21_X1  g544(.A(G92gat), .B1(new_n733_), .B2(new_n623_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n623_), .A2(G92gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n742_), .B2(new_n747_), .ZN(G1337gat));
  OAI21_X1  g547(.A(G99gat), .B1(new_n741_), .B2(new_n435_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n733_), .A2(new_n516_), .A3(new_n410_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g551(.A(new_n735_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT115), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n754_), .A2(new_n755_), .A3(new_n647_), .A4(new_n664_), .ZN(new_n756_));
  OAI21_X1  g555(.A(KEYINPUT115), .B1(new_n738_), .B2(new_n648_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n757_), .A3(G106gat), .ZN(new_n758_));
  XNOR2_X1  g557(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n759_));
  INV_X1    g558(.A(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  NAND4_X1  g560(.A1(new_n756_), .A2(new_n757_), .A3(G106gat), .A4(new_n759_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n761_), .A2(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n733_), .A2(new_n498_), .A3(new_n647_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT53), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT53), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n763_), .A2(new_n767_), .A3(new_n764_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1339gat));
  NOR2_X1   g568(.A1(new_n623_), .A2(new_n262_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n412_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n462_), .A2(new_n460_), .ZN(new_n774_));
  AOI211_X1 g573(.A(new_n469_), .B(new_n774_), .C1(new_n463_), .C2(new_n459_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  OAI21_X1  g576(.A(KEYINPUT119), .B1(new_n574_), .B2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n568_), .A2(new_n579_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(new_n571_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n574_), .A2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT119), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n568_), .A2(new_n783_), .A3(KEYINPUT55), .A4(new_n573_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n778_), .A2(new_n780_), .A3(new_n782_), .A4(new_n784_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(KEYINPUT56), .A3(new_n585_), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT56), .B1(new_n785_), .B2(new_n585_), .ZN(new_n788_));
  OAI211_X1 g587(.A(new_n583_), .B(new_n776_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT58), .ZN(new_n790_));
  OR2_X1    g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n790_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n554_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n583_), .A2(new_n588_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n794_), .A2(new_n776_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n787_), .A2(new_n788_), .A3(KEYINPUT120), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n785_), .A2(KEYINPUT120), .A3(KEYINPUT56), .A4(new_n585_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n477_), .A2(new_n583_), .A3(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n795_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n800_), .A3(new_n611_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n800_), .B1(new_n799_), .B2(new_n611_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n793_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(new_n603_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n605_), .A2(new_n664_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT117), .B(KEYINPUT54), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n807_), .B(new_n808_), .ZN(new_n809_));
  OAI211_X1 g608(.A(new_n772_), .B(new_n773_), .C1(new_n806_), .C2(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n664_), .A2(new_n205_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n804_), .A2(KEYINPUT121), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT121), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n813_), .B(new_n793_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n812_), .A2(new_n604_), .A3(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n809_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n771_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT59), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n810_), .B(new_n811_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(G113gat), .B1(new_n817_), .B2(new_n477_), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n820_), .A2(new_n821_), .ZN(G1340gat));
  INV_X1    g621(.A(G120gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n823_), .B1(new_n654_), .B2(KEYINPUT60), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n817_), .B(new_n824_), .C1(KEYINPUT60), .C2(new_n823_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n810_), .B(new_n591_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n827_), .B2(new_n823_), .ZN(G1341gat));
  AOI21_X1  g627(.A(G127gat), .B1(new_n817_), .B2(new_n603_), .ZN(new_n829_));
  OAI211_X1 g628(.A(new_n810_), .B(G127gat), .C1(new_n817_), .C2(new_n818_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n829_), .B1(new_n831_), .B2(new_n603_), .ZN(G1342gat));
  AND2_X1   g631(.A1(new_n554_), .A2(G134gat), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n810_), .B(new_n833_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT102), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n551_), .B(new_n836_), .ZN(new_n837_));
  AOI21_X1  g636(.A(G134gat), .B1(new_n817_), .B2(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n835_), .A2(new_n838_), .ZN(G1343gat));
  NAND2_X1  g638(.A1(new_n815_), .A2(new_n816_), .ZN(new_n840_));
  NAND4_X1  g639(.A1(new_n840_), .A2(new_n413_), .A3(new_n477_), .A4(new_n770_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n841_), .B(G141gat), .ZN(G1344gat));
  NAND4_X1  g641(.A1(new_n840_), .A2(new_n591_), .A3(new_n413_), .A4(new_n770_), .ZN(new_n843_));
  XNOR2_X1  g642(.A(KEYINPUT123), .B(G148gat), .ZN(new_n844_));
  XNOR2_X1  g643(.A(new_n843_), .B(new_n844_), .ZN(G1345gat));
  NAND4_X1  g644(.A1(new_n840_), .A2(new_n603_), .A3(new_n413_), .A4(new_n770_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(KEYINPUT61), .B(G155gat), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1346gat));
  AND2_X1   g647(.A1(new_n840_), .A2(new_n413_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n849_), .A2(G162gat), .A3(new_n554_), .A4(new_n770_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n840_), .A2(new_n413_), .A3(new_n837_), .A4(new_n770_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n226_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1347gat));
  OAI21_X1  g652(.A(new_n816_), .B1(new_n603_), .B2(new_n805_), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n854_), .A2(new_n648_), .ZN(new_n855_));
  NOR3_X1   g654(.A1(new_n352_), .A2(new_n261_), .A3(new_n435_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT124), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n855_), .A2(new_n315_), .A3(new_n477_), .A4(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n477_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(KEYINPUT125), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n854_), .A2(new_n648_), .A3(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT62), .ZN(new_n862_));
  AND3_X1   g661(.A1(new_n861_), .A2(new_n862_), .A3(G169gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n861_), .B2(G169gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n858_), .B1(new_n863_), .B2(new_n864_), .ZN(G1348gat));
  AOI21_X1  g664(.A(new_n647_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n866_));
  AND4_X1   g665(.A1(G176gat), .A2(new_n866_), .A3(new_n591_), .A4(new_n857_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n855_), .A2(new_n591_), .A3(new_n857_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n284_), .B2(new_n868_), .ZN(G1349gat));
  NAND4_X1  g668(.A1(new_n854_), .A2(new_n603_), .A3(new_n648_), .A4(new_n857_), .ZN(new_n870_));
  MUX2_X1   g669(.A(new_n293_), .B(G183gat), .S(new_n870_), .Z(G1350gat));
  NAND4_X1  g670(.A1(new_n854_), .A2(new_n554_), .A3(new_n648_), .A4(new_n857_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G190gat), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n855_), .A2(new_n857_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n837_), .B1(new_n313_), .B2(new_n312_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n873_), .B1(new_n874_), .B2(new_n875_), .ZN(G1351gat));
  INV_X1    g675(.A(KEYINPUT126), .ZN(new_n877_));
  INV_X1    g676(.A(new_n413_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n878_), .B2(new_n261_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n413_), .A2(KEYINPUT126), .A3(new_n262_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n352_), .B1(new_n879_), .B2(new_n880_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n840_), .A2(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(new_n266_), .A3(new_n477_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n840_), .A2(new_n881_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G197gat), .B1(new_n884_), .B2(new_n664_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n883_), .A2(new_n885_), .ZN(G1352gat));
  INV_X1    g685(.A(new_n268_), .ZN(new_n887_));
  NAND4_X1  g686(.A1(new_n882_), .A2(KEYINPUT127), .A3(new_n591_), .A4(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT127), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n840_), .A2(new_n591_), .A3(new_n881_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(G204gat), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n268_), .ZN(new_n892_));
  OAI21_X1  g691(.A(new_n888_), .B1(new_n891_), .B2(new_n892_), .ZN(G1353gat));
  NOR2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  AND2_X1   g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  NOR4_X1   g694(.A1(new_n884_), .A2(new_n604_), .A3(new_n894_), .A4(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n894_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n882_), .B2(new_n603_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n896_), .A2(new_n898_), .ZN(G1354gat));
  AOI21_X1  g698(.A(G218gat), .B1(new_n882_), .B2(new_n837_), .ZN(new_n900_));
  INV_X1    g699(.A(G218gat), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n884_), .A2(new_n901_), .A3(new_n553_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n900_), .A2(new_n902_), .ZN(G1355gat));
endmodule


