//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 0 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n601_, new_n602_, new_n603_, new_n604_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n813_, new_n814_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n848_, new_n850_, new_n851_, new_n852_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT76), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT1), .ZN(new_n205_));
  NAND3_X1  g004(.A1(KEYINPUT76), .A2(G155gat), .A3(G162gat), .ZN(new_n206_));
  NAND3_X1  g005(.A1(new_n204_), .A2(new_n205_), .A3(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT77), .ZN(new_n208_));
  OR2_X1    g007(.A1(G155gat), .A2(G162gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n206_), .ZN(new_n210_));
  AOI21_X1  g009(.A(KEYINPUT76), .B1(G155gat), .B2(G162gat), .ZN(new_n211_));
  OAI21_X1  g010(.A(KEYINPUT1), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT77), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n204_), .A2(new_n213_), .A3(new_n205_), .A4(new_n206_), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n208_), .A2(new_n209_), .A3(new_n212_), .A4(new_n214_), .ZN(new_n215_));
  XOR2_X1   g014(.A(G141gat), .B(G148gat), .Z(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT3), .ZN(new_n218_));
  INV_X1    g017(.A(G141gat), .ZN(new_n219_));
  INV_X1    g018(.A(G148gat), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n218_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT2), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n221_), .A2(new_n224_), .A3(new_n225_), .A4(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n204_), .A2(new_n206_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n209_), .A3(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n217_), .A2(new_n229_), .ZN(new_n230_));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(G113gat), .ZN(new_n232_));
  INV_X1    g031(.A(G113gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n233_), .A2(KEYINPUT74), .ZN(new_n234_));
  OAI21_X1  g033(.A(G120gat), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  XOR2_X1   g034(.A(G127gat), .B(G134gat), .Z(new_n236_));
  NAND2_X1  g035(.A1(new_n233_), .A2(KEYINPUT74), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n231_), .A2(G113gat), .ZN(new_n238_));
  INV_X1    g037(.A(G120gat), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n237_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n235_), .A2(new_n236_), .A3(new_n240_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n236_), .B1(new_n235_), .B2(new_n240_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n230_), .A2(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n229_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n246_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(new_n243_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n245_), .A2(KEYINPUT4), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G225gat), .A2(G233gat), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT86), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n243_), .B1(new_n217_), .B2(new_n229_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NOR4_X1   g054(.A1(new_n247_), .A2(new_n243_), .A3(KEYINPUT86), .A4(KEYINPUT4), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n249_), .B(new_n251_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT87), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n230_), .A2(new_n254_), .A3(new_n244_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT86), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n253_), .A2(new_n252_), .A3(new_n254_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT87), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n262_), .A2(new_n263_), .A3(new_n251_), .A4(new_n249_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n245_), .A2(new_n250_), .A3(new_n248_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n258_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT0), .B(G57gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(G85gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(G1gat), .B(G29gat), .Z(new_n269_));
  XOR2_X1   g068(.A(new_n268_), .B(new_n269_), .Z(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n270_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n258_), .A2(new_n264_), .A3(new_n272_), .A4(new_n265_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n271_), .A2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT90), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n271_), .A2(KEYINPUT90), .A3(new_n273_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT22), .B(G169gat), .Z(new_n280_));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281_));
  INV_X1    g080(.A(KEYINPUT23), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284_));
  OAI221_X1 g083(.A(new_n279_), .B1(new_n280_), .B2(G176gat), .C1(new_n283_), .C2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(G169gat), .ZN(new_n286_));
  INV_X1    g085(.A(G176gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(KEYINPUT73), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n289_), .B1(G169gat), .B2(G176gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(KEYINPUT24), .A3(new_n279_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n283_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT24), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n288_), .A2(new_n290_), .A3(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT26), .ZN(new_n296_));
  INV_X1    g095(.A(G190gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT25), .B(G183gat), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n292_), .A2(new_n293_), .A3(new_n295_), .A4(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n285_), .A2(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT30), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(new_n244_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G15gat), .B(G43gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT31), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n306_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G71gat), .B(G99gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(G227gat), .A2(G233gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  OR2_X1    g111(.A1(new_n309_), .A2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n309_), .A2(new_n312_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(G204gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(G197gat), .ZN(new_n317_));
  INV_X1    g116(.A(G197gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(G204gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT21), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G211gat), .B(G218gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT21), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n317_), .A2(new_n319_), .A3(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n321_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT80), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n321_), .A2(new_n322_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n321_), .A2(KEYINPUT80), .A3(new_n322_), .A4(new_n324_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n327_), .A2(new_n328_), .A3(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n331_), .B1(KEYINPUT29), .B2(new_n230_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT78), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(G233gat), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT79), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n336_), .A2(G228gat), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(G228gat), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n335_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n230_), .A2(KEYINPUT29), .A3(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G22gat), .B(G50gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n340_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n344_), .B1(new_n247_), .B2(new_n345_), .ZN(new_n346_));
  OR3_X1    g145(.A1(new_n341_), .A2(new_n343_), .A3(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n343_), .B1(new_n341_), .B2(new_n346_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n334_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n347_), .A2(new_n348_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n332_), .B(KEYINPUT78), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  XOR2_X1   g151(.A(G78gat), .B(G106gat), .Z(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT81), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT28), .ZN(new_n355_));
  AND3_X1   g154(.A1(new_n349_), .A2(new_n352_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n355_), .B1(new_n349_), .B2(new_n352_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G8gat), .B(G36gat), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G64gat), .B(G92gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT84), .B(KEYINPUT18), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G226gat), .A2(G233gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT19), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT82), .ZN(new_n368_));
  AND3_X1   g167(.A1(new_n298_), .A2(new_n368_), .A3(new_n299_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n368_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n301_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n294_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n292_), .A3(new_n372_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n285_), .B1(new_n373_), .B2(new_n283_), .ZN(new_n374_));
  OAI211_X1 g173(.A(KEYINPUT20), .B(new_n367_), .C1(new_n374_), .C2(new_n330_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n330_), .A2(new_n304_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT83), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT83), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n330_), .A2(new_n304_), .A3(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n375_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(KEYINPUT20), .B1(new_n330_), .B2(new_n304_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n374_), .A2(new_n330_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n367_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n364_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n386_));
  AND2_X1   g185(.A1(new_n374_), .A2(new_n330_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n366_), .B1(new_n387_), .B2(new_n381_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n364_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n377_), .A2(new_n379_), .ZN(new_n390_));
  OAI211_X1 g189(.A(new_n388_), .B(new_n389_), .C1(new_n390_), .C2(new_n375_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n385_), .A2(new_n386_), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT27), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n380_), .A2(new_n384_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(KEYINPUT85), .A3(new_n389_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n392_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n397_));
  AOI21_X1  g196(.A(new_n397_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n374_), .A2(new_n330_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n367_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n387_), .A2(new_n366_), .A3(new_n381_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n364_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT91), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n391_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n375_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n377_), .A2(new_n379_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n407_), .A2(KEYINPUT91), .A3(new_n389_), .A4(new_n388_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n402_), .A2(new_n404_), .A3(KEYINPUT27), .A4(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n396_), .A2(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n278_), .A2(new_n315_), .A3(new_n359_), .A4(new_n410_), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n271_), .A2(KEYINPUT90), .A3(new_n273_), .ZN(new_n412_));
  AOI21_X1  g211(.A(KEYINPUT90), .B1(new_n271_), .B2(new_n273_), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n410_), .B(new_n358_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT92), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n262_), .A2(new_n250_), .A3(new_n249_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n245_), .A2(new_n251_), .A3(new_n248_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n417_), .A2(new_n270_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n392_), .A2(new_n395_), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n273_), .A2(KEYINPUT33), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n273_), .A2(KEYINPUT33), .ZN(new_n422_));
  OAI211_X1 g221(.A(new_n419_), .B(new_n420_), .C1(new_n421_), .C2(new_n422_), .ZN(new_n423_));
  OAI211_X1 g222(.A(KEYINPUT32), .B(new_n389_), .C1(new_n400_), .C2(new_n401_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT88), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n389_), .A2(KEYINPUT32), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n394_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n425_), .B1(new_n394_), .B2(new_n426_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n274_), .A2(new_n424_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n423_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n359_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n278_), .A2(KEYINPUT92), .A3(new_n358_), .A4(new_n410_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n416_), .A2(new_n432_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT93), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n315_), .B(KEYINPUT75), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n434_), .A2(new_n435_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n411_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT67), .B(G8gat), .ZN(new_n440_));
  INV_X1    g239(.A(G1gat), .ZN(new_n441_));
  OAI21_X1  g240(.A(KEYINPUT14), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT66), .B(G22gat), .ZN(new_n444_));
  INV_X1    g243(.A(G15gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  OR2_X1    g245(.A1(KEYINPUT66), .A2(G22gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(KEYINPUT66), .A2(G22gat), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(G15gat), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n446_), .A2(new_n449_), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT68), .B1(new_n443_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT68), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n442_), .A2(new_n452_), .A3(new_n449_), .A4(new_n446_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n451_), .A2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(G1gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n451_), .A2(new_n441_), .A3(new_n453_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(G8gat), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(G8gat), .B1(new_n455_), .B2(new_n456_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(G57gat), .B(G64gat), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n461_), .A2(KEYINPUT11), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(KEYINPUT11), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G71gat), .B(G78gat), .ZN(new_n464_));
  OR3_X1    g263(.A1(new_n462_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n461_), .A2(new_n464_), .A3(KEYINPUT11), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G231gat), .A2(G233gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n460_), .B(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT17), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT16), .B(G183gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(G211gat), .ZN(new_n474_));
  XOR2_X1   g273(.A(G127gat), .B(G155gat), .Z(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  OR3_X1    g275(.A1(new_n471_), .A2(new_n472_), .A3(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(KEYINPUT17), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n471_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G29gat), .B(G36gat), .ZN(new_n482_));
  INV_X1    g281(.A(G43gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n482_), .B(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(G50gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT15), .ZN(new_n487_));
  NAND2_X1  g286(.A1(G99gat), .A2(G106gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT6), .ZN(new_n489_));
  OAI21_X1  g288(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n490_));
  OR3_X1    g289(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  XOR2_X1   g291(.A(G85gat), .B(G92gat), .Z(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT8), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(KEYINPUT9), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n496_), .A2(new_n489_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G85gat), .A2(G92gat), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT10), .B(G99gat), .ZN(new_n499_));
  OAI221_X1 g298(.A(new_n497_), .B1(KEYINPUT9), .B2(new_n498_), .C1(G106gat), .C2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n495_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n487_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G232gat), .A2(G233gat), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT34), .ZN(new_n504_));
  INV_X1    g303(.A(new_n486_), .ZN(new_n505_));
  OAI221_X1 g304(.A(new_n502_), .B1(KEYINPUT35), .B2(new_n504_), .C1(new_n505_), .C2(new_n501_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(KEYINPUT35), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT64), .B(G134gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n509_), .B(G162gat), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G190gat), .B(G218gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(new_n510_), .B(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n512_), .A2(KEYINPUT36), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n508_), .B(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n512_), .A2(KEYINPUT36), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT37), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n508_), .A2(new_n513_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n517_), .B1(new_n518_), .B2(KEYINPUT65), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n516_), .B(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n439_), .A2(new_n481_), .A3(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT69), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n505_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n455_), .A2(new_n456_), .ZN(new_n525_));
  INV_X1    g324(.A(G8gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n527_), .A2(new_n457_), .A3(new_n486_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n524_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n523_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  AOI211_X1 g331(.A(KEYINPUT69), .B(new_n530_), .C1(new_n524_), .C2(new_n528_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT71), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n487_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n536_), .A2(new_n530_), .A3(new_n528_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G169gat), .B(G197gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT70), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(G113gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(new_n219_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n534_), .A2(new_n535_), .A3(new_n537_), .A4(new_n542_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n458_), .A2(new_n459_), .A3(new_n505_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n486_), .B1(new_n527_), .B2(new_n457_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n531_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT69), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n529_), .A2(new_n523_), .A3(new_n531_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n547_), .A2(new_n537_), .A3(new_n548_), .A4(new_n542_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT71), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n543_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n534_), .A2(new_n537_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n552_), .A2(new_n541_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n551_), .A2(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT72), .ZN(new_n555_));
  INV_X1    g354(.A(G230gat), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(new_n335_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n467_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n501_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n495_), .A2(new_n467_), .A3(new_n500_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(KEYINPUT12), .A3(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT12), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n501_), .A2(new_n562_), .A3(new_n558_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n557_), .B1(new_n561_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n559_), .A2(new_n560_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n564_), .B1(new_n557_), .B2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G120gat), .B(G148gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n567_), .B(new_n316_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT5), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(new_n287_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(new_n566_), .B(new_n570_), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT13), .Z(new_n572_));
  NOR2_X1   g371(.A1(new_n555_), .A2(new_n572_), .ZN(new_n573_));
  AND2_X1   g372(.A1(new_n522_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n278_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n574_), .A2(new_n441_), .A3(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT38), .ZN(new_n577_));
  INV_X1    g376(.A(new_n516_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n439_), .A2(new_n578_), .A3(new_n481_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n551_), .A2(new_n553_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n572_), .A2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n582_), .A2(new_n575_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n577_), .B1(new_n441_), .B2(new_n583_), .ZN(G1324gat));
  INV_X1    g383(.A(KEYINPUT39), .ZN(new_n585_));
  INV_X1    g384(.A(new_n410_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n526_), .B1(new_n582_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT94), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n587_), .A2(new_n588_), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n585_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n591_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(KEYINPUT39), .A3(new_n589_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n574_), .A2(new_n440_), .A3(new_n586_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n592_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT40), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n592_), .A2(new_n594_), .A3(KEYINPUT40), .A4(new_n595_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(G1325gat));
  INV_X1    g399(.A(new_n436_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n445_), .B1(new_n582_), .B2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT41), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n574_), .A2(new_n445_), .A3(new_n601_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(G1326gat));
  INV_X1    g404(.A(G22gat), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n606_), .B1(new_n582_), .B2(new_n358_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT42), .ZN(new_n608_));
  AND3_X1   g407(.A1(new_n574_), .A2(new_n606_), .A3(new_n358_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(KEYINPUT95), .ZN(G1327gat));
  NAND2_X1  g410(.A1(new_n439_), .A2(new_n516_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n612_), .A2(new_n572_), .A3(new_n555_), .ZN(new_n613_));
  INV_X1    g412(.A(G29gat), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n613_), .A2(new_n614_), .A3(new_n575_), .A4(new_n480_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n581_), .A2(new_n480_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT43), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n439_), .A2(new_n618_), .A3(new_n520_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n618_), .B1(new_n439_), .B2(new_n520_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n617_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT96), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  XOR2_X1   g422(.A(KEYINPUT97), .B(KEYINPUT44), .Z(new_n624_));
  OAI211_X1 g423(.A(KEYINPUT96), .B(new_n617_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n620_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n439_), .A2(new_n618_), .A3(new_n520_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n616_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n278_), .B1(new_n629_), .B2(KEYINPUT44), .ZN(new_n630_));
  AND3_X1   g429(.A1(new_n626_), .A2(KEYINPUT98), .A3(new_n630_), .ZN(new_n631_));
  AOI21_X1  g430(.A(KEYINPUT98), .B1(new_n626_), .B2(new_n630_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT99), .B1(new_n633_), .B2(G29gat), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n635_));
  NOR4_X1   g434(.A1(new_n631_), .A2(new_n632_), .A3(new_n635_), .A4(new_n614_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n615_), .B1(new_n634_), .B2(new_n636_), .ZN(G1328gat));
  NAND2_X1  g436(.A1(new_n613_), .A2(new_n480_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(G36gat), .A3(new_n410_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT45), .Z(new_n640_));
  NAND2_X1  g439(.A1(new_n629_), .A2(KEYINPUT44), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n626_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G36gat), .B1(new_n642_), .B2(new_n410_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT46), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n640_), .A2(KEYINPUT46), .A3(new_n643_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1329gat));
  OAI21_X1  g447(.A(new_n483_), .B1(new_n638_), .B2(new_n436_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT100), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n626_), .A2(G43gat), .A3(new_n315_), .A4(new_n641_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g452(.A(G50gat), .B1(new_n642_), .B2(new_n359_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n613_), .A2(new_n485_), .A3(new_n480_), .ZN(new_n655_));
  OAI21_X1  g454(.A(new_n654_), .B1(new_n359_), .B2(new_n655_), .ZN(G1331gat));
  INV_X1    g455(.A(new_n572_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(new_n554_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n522_), .A2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(G57gat), .B1(new_n659_), .B2(new_n575_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n579_), .A2(new_n572_), .A3(new_n555_), .ZN(new_n661_));
  INV_X1    g460(.A(G57gat), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n661_), .A2(new_n662_), .A3(new_n278_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n660_), .A2(new_n663_), .ZN(G1332gat));
  OAI21_X1  g463(.A(G64gat), .B1(new_n661_), .B2(new_n410_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT48), .ZN(new_n666_));
  INV_X1    g465(.A(G64gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n659_), .A2(new_n667_), .A3(new_n586_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1333gat));
  OAI21_X1  g468(.A(G71gat), .B1(new_n661_), .B2(new_n436_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n670_), .B(KEYINPUT101), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT49), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n436_), .A2(G71gat), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT102), .Z(new_n674_));
  NAND2_X1  g473(.A1(new_n659_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(new_n675_), .ZN(G1334gat));
  OAI21_X1  g475(.A(G78gat), .B1(new_n661_), .B2(new_n359_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT50), .ZN(new_n678_));
  INV_X1    g477(.A(G78gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n659_), .A2(new_n679_), .A3(new_n358_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1335gat));
  NAND2_X1  g480(.A1(new_n658_), .A2(new_n480_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n612_), .A2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(G85gat), .B1(new_n683_), .B2(new_n575_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n682_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n685_), .A2(KEYINPUT103), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(KEYINPUT103), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n575_), .A2(G85gat), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT104), .Z(new_n690_));
  AOI21_X1  g489(.A(new_n684_), .B1(new_n688_), .B2(new_n690_), .ZN(G1336gat));
  INV_X1    g490(.A(G92gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n683_), .A2(new_n692_), .A3(new_n586_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n410_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(new_n692_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT105), .ZN(G1337gat));
  NAND2_X1  g495(.A1(new_n685_), .A2(new_n601_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n315_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n698_), .A2(new_n499_), .ZN(new_n699_));
  AOI22_X1  g498(.A1(new_n697_), .A2(G99gat), .B1(new_n683_), .B2(new_n699_), .ZN(new_n700_));
  XOR2_X1   g499(.A(new_n700_), .B(KEYINPUT51), .Z(G1338gat));
  INV_X1    g500(.A(new_n685_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G106gat), .B1(new_n702_), .B2(new_n359_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT52), .ZN(new_n704_));
  OR2_X1    g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n704_), .ZN(new_n706_));
  NOR4_X1   g505(.A1(new_n612_), .A2(G106gat), .A3(new_n359_), .A4(new_n682_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT106), .Z(new_n708_));
  NAND3_X1  g507(.A1(new_n705_), .A2(new_n706_), .A3(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g509(.A1(new_n278_), .A2(new_n586_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n561_), .A2(new_n557_), .A3(new_n563_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n712_), .A2(KEYINPUT55), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT110), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT110), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n712_), .A2(new_n715_), .A3(KEYINPUT55), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n564_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n570_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n714_), .A2(new_n564_), .A3(new_n716_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n719_), .A2(new_n720_), .A3(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT56), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n719_), .A2(KEYINPUT56), .A3(new_n720_), .A4(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n566_), .A2(new_n570_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n536_), .A2(new_n528_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n536_), .A2(KEYINPUT111), .A3(new_n528_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n730_), .A2(new_n531_), .A3(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n529_), .A2(new_n530_), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(new_n541_), .A3(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  AND4_X1   g534(.A1(KEYINPUT112), .A2(new_n551_), .A3(new_n727_), .A4(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n734_), .B1(new_n543_), .B2(new_n550_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT112), .B1(new_n737_), .B2(new_n727_), .ZN(new_n738_));
  OAI211_X1 g537(.A(KEYINPUT113), .B(new_n726_), .C1(new_n736_), .C2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT58), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n551_), .A2(new_n727_), .A3(new_n735_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT112), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n737_), .A2(KEYINPUT112), .A3(new_n727_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(KEYINPUT113), .B1(new_n746_), .B2(new_n726_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n520_), .B1(new_n741_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n746_), .A2(KEYINPUT58), .A3(new_n726_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT114), .B(new_n520_), .C1(new_n741_), .C2(new_n747_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n750_), .A2(new_n751_), .A3(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n554_), .A2(new_n727_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT109), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n554_), .A2(KEYINPUT109), .A3(new_n727_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n756_), .A2(new_n726_), .A3(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n737_), .A2(new_n571_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n516_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT57), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n760_), .B(new_n761_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n481_), .B1(new_n753_), .B2(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n554_), .A2(KEYINPUT72), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n554_), .A2(KEYINPUT72), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n481_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT107), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n555_), .A2(KEYINPUT107), .A3(new_n481_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n520_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT108), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(KEYINPUT54), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n572_), .B1(new_n771_), .B2(KEYINPUT54), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n770_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n772_), .B1(new_n770_), .B2(new_n773_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n359_), .B(new_n711_), .C1(new_n763_), .C2(new_n776_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n777_), .A2(new_n580_), .A3(new_n698_), .ZN(new_n778_));
  OAI21_X1  g577(.A(KEYINPUT115), .B1(new_n778_), .B2(G113gat), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT115), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n753_), .A2(new_n762_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n480_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n776_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n784_), .A2(new_n315_), .A3(new_n359_), .A4(new_n711_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n780_), .B(new_n233_), .C1(new_n785_), .C2(new_n580_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n779_), .A2(new_n786_), .ZN(new_n787_));
  XNOR2_X1  g586(.A(KEYINPUT116), .B(G113gat), .ZN(new_n788_));
  INV_X1    g587(.A(new_n711_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n790_));
  NAND4_X1  g589(.A1(new_n790_), .A2(KEYINPUT59), .A3(new_n315_), .A4(new_n359_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT59), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n792_), .B1(new_n777_), .B2(new_n698_), .ZN(new_n793_));
  AOI211_X1 g592(.A(new_n555_), .B(new_n788_), .C1(new_n791_), .C2(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n787_), .A2(new_n794_), .ZN(G1340gat));
  INV_X1    g594(.A(new_n785_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n239_), .B1(new_n657_), .B2(KEYINPUT60), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n796_), .B(new_n797_), .C1(KEYINPUT60), .C2(new_n239_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n657_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n239_), .ZN(G1341gat));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801_));
  NOR3_X1   g600(.A1(new_n777_), .A2(new_n698_), .A3(new_n480_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(G127gat), .ZN(new_n803_));
  INV_X1    g602(.A(G127gat), .ZN(new_n804_));
  OAI211_X1 g603(.A(KEYINPUT117), .B(new_n804_), .C1(new_n785_), .C2(new_n480_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n804_), .B(new_n480_), .C1(new_n791_), .C2(new_n793_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(G1342gat));
  AOI21_X1  g607(.A(G134gat), .B1(new_n796_), .B2(new_n516_), .ZN(new_n809_));
  INV_X1    g608(.A(G134gat), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n810_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n809_), .B1(new_n811_), .B2(new_n520_), .ZN(G1343gat));
  NAND2_X1  g611(.A1(new_n790_), .A2(new_n436_), .ZN(new_n813_));
  NOR3_X1   g612(.A1(new_n813_), .A2(new_n580_), .A3(new_n359_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(new_n219_), .ZN(G1344gat));
  NOR3_X1   g614(.A1(new_n813_), .A2(new_n657_), .A3(new_n359_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(KEYINPUT118), .B(G148gat), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n816_), .B(new_n817_), .ZN(G1345gat));
  NOR3_X1   g617(.A1(new_n813_), .A2(new_n359_), .A3(new_n480_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(KEYINPUT119), .B(KEYINPUT61), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n820_), .B(G155gat), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n819_), .B(new_n822_), .ZN(G1346gat));
  NOR2_X1   g622(.A1(new_n813_), .A2(new_n359_), .ZN(new_n824_));
  AND3_X1   g623(.A1(new_n824_), .A2(G162gat), .A3(new_n520_), .ZN(new_n825_));
  AOI21_X1  g624(.A(G162gat), .B1(new_n824_), .B2(new_n516_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(G1347gat));
  INV_X1    g626(.A(KEYINPUT62), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n601_), .A2(new_n278_), .A3(new_n359_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n784_), .A2(new_n554_), .A3(new_n586_), .A4(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n829_), .B1(new_n832_), .B2(G169gat), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n586_), .B(new_n831_), .C1(new_n763_), .C2(new_n776_), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n829_), .B(G169gat), .C1(new_n834_), .C2(new_n580_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n828_), .B1(new_n833_), .B2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n834_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n580_), .A2(new_n280_), .ZN(new_n839_));
  XOR2_X1   g638(.A(new_n839_), .B(KEYINPUT121), .Z(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(G169gat), .B1(new_n834_), .B2(new_n580_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(KEYINPUT120), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n843_), .A2(KEYINPUT62), .A3(new_n835_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n837_), .A2(new_n841_), .A3(new_n844_), .ZN(G1348gat));
  NOR2_X1   g644(.A1(new_n834_), .A2(new_n657_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(new_n287_), .ZN(G1349gat));
  NOR2_X1   g646(.A1(new_n834_), .A2(new_n480_), .ZN(new_n848_));
  MUX2_X1   g647(.A(G183gat), .B(new_n301_), .S(new_n848_), .Z(G1350gat));
  OAI211_X1 g648(.A(new_n838_), .B(new_n516_), .C1(new_n370_), .C2(new_n369_), .ZN(new_n850_));
  OAI21_X1  g649(.A(G190gat), .B1(new_n834_), .B2(new_n521_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(KEYINPUT122), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT122), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n850_), .A2(new_n854_), .A3(new_n851_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n853_), .A2(new_n855_), .ZN(G1351gat));
  NOR2_X1   g655(.A1(KEYINPUT123), .A2(G197gat), .ZN(new_n857_));
  XOR2_X1   g656(.A(KEYINPUT123), .B(G197gat), .Z(new_n858_));
  OAI211_X1 g657(.A(new_n436_), .B(new_n586_), .C1(new_n763_), .C2(new_n776_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n278_), .A2(new_n358_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n861_), .A2(new_n554_), .ZN(new_n862_));
  MUX2_X1   g661(.A(new_n857_), .B(new_n858_), .S(new_n862_), .Z(G1352gat));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n572_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT124), .B(G204gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1353gat));
  OAI21_X1  g665(.A(KEYINPUT126), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR3_X1   g667(.A1(KEYINPUT126), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n480_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT125), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n861_), .A2(new_n872_), .ZN(new_n873_));
  MUX2_X1   g672(.A(new_n870_), .B(new_n868_), .S(new_n873_), .Z(G1354gat));
  INV_X1    g673(.A(G218gat), .ZN(new_n875_));
  NOR4_X1   g674(.A1(new_n859_), .A2(new_n875_), .A3(new_n860_), .A4(new_n521_), .ZN(new_n876_));
  INV_X1    g675(.A(KEYINPUT127), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n877_), .B1(new_n861_), .B2(new_n516_), .ZN(new_n878_));
  NOR4_X1   g677(.A1(new_n859_), .A2(KEYINPUT127), .A3(new_n860_), .A4(new_n578_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n876_), .B1(new_n880_), .B2(new_n875_), .ZN(G1355gat));
endmodule


