//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n716_, new_n717_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n869_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n908_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  INV_X1    g001(.A(G92gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT18), .B(G64gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  NAND2_X1  g005(.A1(G226gat), .A2(G233gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT19), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n210_));
  INV_X1    g009(.A(G169gat), .ZN(new_n211_));
  INV_X1    g010(.A(G176gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G183gat), .A2(G190gat), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n217_));
  AND2_X1   g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n211_), .A2(new_n212_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G169gat), .A2(G176gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n213_), .B(new_n218_), .C1(new_n221_), .C2(new_n210_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT26), .B(G190gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n225_));
  NAND2_X1  g024(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT87), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT87), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n225_), .A2(new_n229_), .A3(new_n226_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n224_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n220_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(KEYINPUT22), .B(G169gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n232_), .B1(new_n233_), .B2(new_n212_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n234_), .A2(KEYINPUT89), .ZN(new_n235_));
  OAI211_X1 g034(.A(new_n216_), .B(new_n217_), .C1(G183gat), .C2(G190gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT89), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n236_), .B1(new_n237_), .B2(new_n232_), .ZN(new_n238_));
  OAI22_X1  g037(.A1(new_n222_), .A2(new_n231_), .B1(new_n235_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G197gat), .B(G204gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G211gat), .B(G218gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT21), .ZN(new_n242_));
  OR3_X1    g041(.A1(new_n240_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n241_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n244_));
  AND2_X1   g043(.A1(new_n240_), .A2(new_n242_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n239_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT90), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n239_), .A2(KEYINPUT90), .A3(new_n246_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT86), .ZN(new_n252_));
  INV_X1    g051(.A(new_n246_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n227_), .A2(new_n223_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n219_), .A2(KEYINPUT24), .A3(new_n220_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n254_), .A2(new_n218_), .A3(new_n255_), .A4(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n234_), .A2(new_n236_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n259_), .A2(KEYINPUT79), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT79), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n257_), .A2(new_n258_), .A3(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n253_), .A2(new_n260_), .A3(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n252_), .B1(new_n263_), .B2(KEYINPUT20), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n251_), .A2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n252_), .A3(KEYINPUT20), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n209_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n239_), .A2(new_n246_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n260_), .A2(new_n262_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n268_), .B(KEYINPUT20), .C1(new_n269_), .C2(new_n253_), .ZN(new_n270_));
  NOR2_X1   g069(.A1(new_n270_), .A2(new_n208_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n206_), .B1(new_n267_), .B2(new_n271_), .ZN(new_n272_));
  OR2_X1    g071(.A1(new_n270_), .A2(new_n208_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n206_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n266_), .ZN(new_n275_));
  NOR3_X1   g074(.A1(new_n275_), .A2(new_n251_), .A3(new_n264_), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n273_), .B(new_n274_), .C1(new_n276_), .C2(new_n209_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n272_), .A2(KEYINPUT91), .A3(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n267_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT91), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n279_), .A2(new_n280_), .A3(new_n274_), .A4(new_n273_), .ZN(new_n281_));
  XOR2_X1   g080(.A(KEYINPUT96), .B(KEYINPUT27), .Z(new_n282_));
  NAND3_X1  g081(.A1(new_n278_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT95), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(new_n270_), .B2(new_n208_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n265_), .A2(new_n266_), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n285_), .B1(new_n286_), .B2(new_n208_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n270_), .A2(new_n284_), .A3(new_n208_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(new_n206_), .A3(new_n288_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(KEYINPUT27), .A3(new_n277_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n283_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n291_), .A2(KEYINPUT98), .ZN(new_n292_));
  INV_X1    g091(.A(KEYINPUT98), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n283_), .A2(new_n290_), .A3(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(KEYINPUT30), .B(G15gat), .Z(new_n295_));
  XNOR2_X1  g094(.A(new_n269_), .B(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G227gat), .A2(G233gat), .ZN(new_n297_));
  XOR2_X1   g096(.A(new_n297_), .B(KEYINPUT82), .Z(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT31), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n296_), .A2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G127gat), .B(G134gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G113gat), .B(G120gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(KEYINPUT80), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G127gat), .B(G134gat), .Z(new_n306_));
  XOR2_X1   g105(.A(G113gat), .B(G120gat), .Z(new_n307_));
  NAND2_X1  g106(.A1(new_n306_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(KEYINPUT81), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n302_), .A2(new_n303_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT81), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n305_), .B1(new_n309_), .B2(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n308_), .A2(KEYINPUT81), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n310_), .A2(new_n311_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(new_n315_), .A3(new_n304_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n313_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G71gat), .B(G99gat), .ZN(new_n318_));
  INV_X1    g117(.A(G43gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n317_), .B(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n296_), .A2(new_n299_), .ZN(new_n323_));
  OR3_X1    g122(.A1(new_n301_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n322_), .B1(new_n301_), .B2(new_n323_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT2), .ZN(new_n328_));
  OR4_X1    g127(.A1(KEYINPUT83), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n329_));
  OR2_X1    g128(.A1(G141gat), .A2(G148gat), .ZN(new_n330_));
  OAI21_X1  g129(.A(KEYINPUT3), .B1(new_n330_), .B2(KEYINPUT83), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n328_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n332_));
  OR2_X1    g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G155gat), .A2(G162gat), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n332_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  AND3_X1   g134(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n336_));
  AOI21_X1  g135(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n337_));
  OAI21_X1  g136(.A(new_n333_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n338_), .A2(new_n327_), .A3(new_n330_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n317_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n302_), .A2(new_n303_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n308_), .A2(new_n342_), .ZN(new_n343_));
  AND3_X1   g142(.A1(new_n335_), .A2(new_n339_), .A3(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n341_), .A2(new_n345_), .A3(KEYINPUT92), .A4(KEYINPUT4), .ZN(new_n346_));
  AOI22_X1  g145(.A1(new_n313_), .A2(new_n316_), .B1(new_n339_), .B2(new_n335_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT4), .ZN(new_n348_));
  NOR3_X1   g147(.A1(new_n347_), .A2(new_n348_), .A3(new_n344_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n316_), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n304_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n348_), .B(new_n340_), .C1(new_n350_), .C2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT92), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n346_), .B1(new_n349_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G225gat), .A2(G233gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n356_), .B(KEYINPUT93), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  OR3_X1    g157(.A1(new_n347_), .A2(new_n357_), .A3(new_n344_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G1gat), .B(G29gat), .Z(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(G85gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT0), .B(G57gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n364_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n358_), .A2(new_n359_), .A3(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n335_), .A2(new_n339_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(KEYINPUT84), .B(KEYINPUT29), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n246_), .B1(new_n369_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n371_), .A2(G228gat), .A3(G233gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G228gat), .A2(G233gat), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n373_), .B(new_n246_), .C1(new_n369_), .C2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n372_), .A2(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G78gat), .B(G106gat), .Z(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n372_), .A2(new_n375_), .A3(new_n377_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n340_), .A2(KEYINPUT29), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G22gat), .B(G50gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n383_), .B(KEYINPUT28), .Z(new_n384_));
  XNOR2_X1  g183(.A(new_n382_), .B(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n377_), .B1(new_n372_), .B2(new_n375_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT85), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n385_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n381_), .A2(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n379_), .A2(new_n387_), .A3(new_n380_), .A4(new_n385_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n326_), .A2(new_n368_), .A3(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n292_), .A2(new_n294_), .A3(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(KEYINPUT99), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT99), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n292_), .A2(new_n392_), .A3(new_n395_), .A4(new_n294_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n389_), .A2(new_n390_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT33), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n367_), .A2(new_n398_), .ZN(new_n399_));
  NAND4_X1  g198(.A1(new_n358_), .A2(KEYINPUT33), .A3(new_n359_), .A4(new_n366_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n347_), .A2(new_n344_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n366_), .B1(new_n401_), .B2(new_n357_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n355_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n402_), .B1(new_n403_), .B2(new_n357_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n399_), .A2(new_n400_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(new_n281_), .B2(new_n278_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n287_), .A2(KEYINPUT32), .A3(new_n274_), .A4(new_n288_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n274_), .A2(KEYINPUT32), .ZN(new_n408_));
  OAI211_X1 g207(.A(new_n273_), .B(new_n408_), .C1(new_n276_), .C2(new_n209_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT94), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n279_), .A2(KEYINPUT94), .A3(new_n273_), .A4(new_n408_), .ZN(new_n412_));
  AND4_X1   g211(.A1(new_n368_), .A2(new_n407_), .A3(new_n411_), .A4(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n397_), .B1(new_n406_), .B2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n397_), .A2(new_n368_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(new_n283_), .A3(new_n290_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n416_), .A2(KEYINPUT97), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT97), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n415_), .A2(new_n283_), .A3(new_n290_), .A4(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n414_), .A2(new_n417_), .A3(new_n419_), .ZN(new_n420_));
  AOI22_X1  g219(.A1(new_n394_), .A2(new_n396_), .B1(new_n420_), .B2(new_n326_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(G71gat), .B(G78gat), .ZN(new_n422_));
  INV_X1    g221(.A(G57gat), .ZN(new_n423_));
  INV_X1    g222(.A(G64gat), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G57gat), .A2(G64gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n422_), .B1(KEYINPUT11), .B2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT11), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n425_), .A2(new_n429_), .A3(new_n426_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n427_), .A2(new_n422_), .A3(KEYINPUT11), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G99gat), .A2(G106gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT6), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT10), .B(G99gat), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n436_), .B(new_n437_), .C1(new_n438_), .C2(G106gat), .ZN(new_n439_));
  NAND3_X1  g238(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(G85gat), .B2(G92gat), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT64), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(new_n203_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n443_), .A2(G85gat), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT9), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n441_), .B1(new_n447_), .B2(KEYINPUT65), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT65), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n445_), .A2(new_n449_), .A3(new_n446_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n439_), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT7), .ZN(new_n452_));
  INV_X1    g251(.A(G99gat), .ZN(new_n453_));
  INV_X1    g252(.A(G106gat), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n452_), .A2(new_n453_), .A3(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n456_));
  NAND4_X1  g255(.A1(new_n455_), .A2(new_n436_), .A3(new_n437_), .A4(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT8), .ZN(new_n458_));
  XOR2_X1   g257(.A(G85gat), .B(G92gat), .Z(new_n459_));
  AND3_X1   g258(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n458_), .B1(new_n457_), .B2(new_n459_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n433_), .B1(new_n451_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n457_), .A2(new_n459_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT8), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n457_), .A2(new_n458_), .A3(new_n459_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n431_), .A2(new_n432_), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n445_), .A2(new_n449_), .A3(new_n446_), .ZN(new_n469_));
  AOI21_X1  g268(.A(new_n449_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n470_));
  NOR3_X1   g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n441_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n467_), .B(new_n468_), .C1(new_n471_), .C2(new_n439_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n463_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(G230gat), .ZN(new_n474_));
  INV_X1    g273(.A(G233gat), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n477_), .A2(KEYINPUT66), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT66), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n473_), .A2(new_n479_), .A3(new_n476_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n478_), .A2(new_n480_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n463_), .A2(new_n472_), .A3(KEYINPUT12), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT12), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n483_), .B(new_n433_), .C1(new_n451_), .C2(new_n462_), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n476_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT69), .B1(new_n481_), .B2(new_n485_), .ZN(new_n486_));
  XOR2_X1   g285(.A(G176gat), .B(G204gat), .Z(new_n487_));
  XNOR2_X1  g286(.A(G120gat), .B(G148gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  INV_X1    g290(.A(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT67), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n482_), .A2(new_n484_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n476_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT69), .ZN(new_n498_));
  NAND4_X1  g297(.A1(new_n497_), .A2(new_n478_), .A3(new_n498_), .A4(new_n480_), .ZN(new_n499_));
  AND3_X1   g298(.A1(new_n486_), .A2(new_n494_), .A3(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n494_), .B1(new_n486_), .B2(new_n499_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  OR2_X1    g301(.A1(new_n502_), .A2(KEYINPUT13), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(KEYINPUT13), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G169gat), .B(G197gat), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n507_), .B(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G229gat), .A2(G233gat), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(KEYINPUT72), .A2(G15gat), .ZN(new_n512_));
  NOR2_X1   g311(.A1(KEYINPUT72), .A2(G15gat), .ZN(new_n513_));
  OAI21_X1  g312(.A(G22gat), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(KEYINPUT73), .A2(G8gat), .ZN(new_n515_));
  NOR2_X1   g314(.A1(KEYINPUT73), .A2(G8gat), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT14), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT72), .ZN(new_n518_));
  INV_X1    g317(.A(G15gat), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(G22gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(KEYINPUT72), .A2(G15gat), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n520_), .A2(new_n521_), .A3(new_n522_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n514_), .A2(new_n517_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(G1gat), .ZN(new_n525_));
  INV_X1    g324(.A(G8gat), .ZN(new_n526_));
  NOR2_X1   g325(.A1(KEYINPUT14), .A2(G1gat), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n514_), .A2(new_n523_), .A3(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n525_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G43gat), .B(G50gat), .Z(new_n531_));
  INV_X1    g330(.A(KEYINPUT70), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(G43gat), .B(G50gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT70), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G29gat), .B(G36gat), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n533_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n526_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n542_));
  NOR3_X1   g341(.A1(new_n530_), .A2(new_n541_), .A3(new_n542_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n533_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n537_), .B1(new_n533_), .B2(new_n535_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n525_), .A2(new_n528_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(G8gat), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n546_), .B1(new_n548_), .B2(new_n529_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n511_), .B1(new_n543_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT76), .ZN(new_n551_));
  INV_X1    g350(.A(new_n543_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n541_), .B(KEYINPUT15), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n530_), .A2(new_n542_), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n552_), .B(new_n510_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT76), .ZN(new_n557_));
  OAI211_X1 g356(.A(new_n557_), .B(new_n511_), .C1(new_n543_), .C2(new_n549_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n509_), .B1(new_n556_), .B2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n509_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n551_), .A2(new_n555_), .A3(new_n558_), .A4(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n560_), .A2(KEYINPUT77), .A3(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT77), .ZN(new_n564_));
  OAI211_X1 g363(.A(new_n564_), .B(new_n509_), .C1(new_n556_), .C2(new_n559_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  XOR2_X1   g365(.A(new_n566_), .B(KEYINPUT78), .Z(new_n567_));
  NOR3_X1   g366(.A1(new_n421_), .A2(new_n506_), .A3(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n451_), .A2(new_n462_), .ZN(new_n569_));
  OR2_X1    g368(.A1(new_n553_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G232gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT34), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT35), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n569_), .A2(new_n546_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n572_), .A2(KEYINPUT35), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n570_), .A2(new_n573_), .A3(new_n574_), .A4(new_n575_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n553_), .A2(new_n569_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n574_), .ZN(new_n578_));
  OAI211_X1 g377(.A(KEYINPUT35), .B(new_n572_), .C1(new_n577_), .C2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(G190gat), .B(G218gat), .Z(new_n581_));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT36), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  OR2_X1    g384(.A1(new_n580_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n580_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n583_), .B(new_n584_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n586_), .B(KEYINPUT37), .C1(new_n587_), .C2(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n580_), .A2(new_n585_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n587_), .A2(KEYINPUT71), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT71), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n588_), .B1(new_n580_), .B2(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n590_), .B1(new_n591_), .B2(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n589_), .B1(new_n594_), .B2(KEYINPUT37), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n554_), .B(new_n596_), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(new_n433_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G127gat), .B(G155gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(G211gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT16), .B(G183gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n602_), .B(KEYINPUT17), .Z(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n604_), .A2(KEYINPUT75), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n604_), .A2(KEYINPUT75), .ZN(new_n606_));
  XOR2_X1   g405(.A(KEYINPUT74), .B(KEYINPUT17), .Z(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  OAI22_X1  g407(.A1(new_n605_), .A2(new_n606_), .B1(new_n598_), .B2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n595_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n568_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n368_), .ZN(new_n612_));
  NOR3_X1   g411(.A1(new_n611_), .A2(G1gat), .A3(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT38), .Z(new_n614_));
  XOR2_X1   g413(.A(new_n594_), .B(KEYINPUT101), .Z(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n421_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n566_), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT100), .B1(new_n505_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT100), .ZN(new_n621_));
  AOI211_X1 g420(.A(new_n621_), .B(new_n566_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n620_), .A2(new_n622_), .A3(new_n609_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n618_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n626_), .B2(new_n612_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT102), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n627_), .A2(new_n628_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n614_), .A2(new_n629_), .A3(new_n630_), .ZN(G1324gat));
  NAND2_X1  g430(.A1(new_n292_), .A2(new_n294_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n632_), .B1(new_n516_), .B2(new_n515_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n611_), .A2(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n394_), .A2(new_n396_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n420_), .A2(new_n326_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n637_), .A2(new_n623_), .A3(new_n632_), .A4(new_n615_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT103), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n617_), .A2(KEYINPUT103), .A3(new_n632_), .A4(new_n623_), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(G8gat), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n642_), .A2(KEYINPUT39), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n640_), .A2(new_n641_), .A3(new_n644_), .A4(G8gat), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n634_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n647_));
  INV_X1    g446(.A(new_n647_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n646_), .B(new_n648_), .ZN(G1325gat));
  NOR2_X1   g448(.A1(new_n626_), .A2(new_n326_), .ZN(new_n650_));
  OR3_X1    g449(.A1(new_n650_), .A2(KEYINPUT41), .A3(new_n519_), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT41), .B1(new_n650_), .B2(new_n519_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n611_), .A2(G15gat), .A3(new_n326_), .ZN(new_n653_));
  OR2_X1    g452(.A1(new_n653_), .A2(KEYINPUT105), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(KEYINPUT105), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n651_), .A2(new_n652_), .A3(new_n654_), .A4(new_n655_), .ZN(G1326gat));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n397_), .B(KEYINPUT106), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n625_), .A2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n657_), .B1(new_n660_), .B2(G22gat), .ZN(new_n661_));
  AOI211_X1 g460(.A(KEYINPUT42), .B(new_n521_), .C1(new_n625_), .C2(new_n659_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n659_), .A2(new_n521_), .ZN(new_n663_));
  OAI22_X1  g462(.A1(new_n661_), .A2(new_n662_), .B1(new_n611_), .B2(new_n663_), .ZN(G1327gat));
  INV_X1    g463(.A(G29gat), .ZN(new_n665_));
  INV_X1    g464(.A(new_n609_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n594_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n568_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n669_), .B2(new_n612_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n595_), .B(KEYINPUT107), .Z(new_n671_));
  OAI21_X1  g470(.A(KEYINPUT43), .B1(new_n421_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n595_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(KEYINPUT43), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n637_), .A2(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n672_), .A2(new_n675_), .ZN(new_n676_));
  NOR3_X1   g475(.A1(new_n620_), .A2(new_n622_), .A3(new_n666_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n680_), .A2(G29gat), .A3(new_n368_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n677_), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n679_), .B(new_n682_), .C1(new_n672_), .C2(new_n675_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n670_), .B1(new_n681_), .B2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(KEYINPUT108), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n686_), .B(new_n670_), .C1(new_n681_), .C2(new_n683_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(G1328gat));
  INV_X1    g487(.A(G36gat), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n568_), .A2(new_n689_), .A3(new_n632_), .A4(new_n668_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT45), .ZN(new_n691_));
  INV_X1    g490(.A(new_n632_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n682_), .B1(new_n672_), .B2(new_n675_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT44), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n693_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(KEYINPUT46), .B(new_n691_), .C1(new_n696_), .C2(new_n689_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  INV_X1    g497(.A(new_n691_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n689_), .B1(new_n693_), .B2(new_n695_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n697_), .A2(new_n701_), .ZN(G1329gat));
  NOR2_X1   g501(.A1(new_n326_), .A2(new_n319_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n703_), .B1(new_n694_), .B2(KEYINPUT44), .ZN(new_n704_));
  OAI21_X1  g503(.A(KEYINPUT109), .B1(new_n704_), .B2(new_n683_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n680_), .A2(new_n706_), .A3(new_n695_), .A4(new_n703_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n319_), .B1(new_n669_), .B2(new_n326_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n705_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT47), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT47), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n705_), .A2(new_n707_), .A3(new_n711_), .A4(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(G1330gat));
  NAND3_X1  g512(.A1(new_n680_), .A2(new_n391_), .A3(new_n695_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n714_), .A2(G50gat), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n658_), .A2(G50gat), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT110), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n715_), .B1(new_n669_), .B2(new_n717_), .ZN(G1331gat));
  NAND4_X1  g517(.A1(new_n617_), .A2(new_n666_), .A3(new_n506_), .A4(new_n567_), .ZN(new_n719_));
  NOR3_X1   g518(.A1(new_n719_), .A2(new_n423_), .A3(new_n612_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n505_), .A2(new_n619_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n421_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n610_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT111), .Z(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n368_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n720_), .B1(new_n726_), .B2(new_n423_), .ZN(G1332gat));
  OAI21_X1  g526(.A(G64gat), .B1(new_n719_), .B2(new_n692_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT48), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n725_), .A2(new_n424_), .A3(new_n632_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1333gat));
  INV_X1    g530(.A(G71gat), .ZN(new_n732_));
  INV_X1    g531(.A(new_n326_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n725_), .A2(new_n732_), .A3(new_n733_), .ZN(new_n734_));
  OAI21_X1  g533(.A(G71gat), .B1(new_n719_), .B2(new_n326_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(KEYINPUT49), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(KEYINPUT49), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n734_), .B1(new_n736_), .B2(new_n737_), .ZN(G1334gat));
  OAI21_X1  g537(.A(G78gat), .B1(new_n719_), .B2(new_n658_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT50), .ZN(new_n740_));
  INV_X1    g539(.A(G78gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n725_), .A2(new_n741_), .A3(new_n659_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n740_), .A2(new_n742_), .ZN(G1335gat));
  INV_X1    g542(.A(KEYINPUT113), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n721_), .A2(new_n609_), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n676_), .B2(new_n746_), .ZN(new_n747_));
  AOI211_X1 g546(.A(KEYINPUT113), .B(new_n745_), .C1(new_n672_), .C2(new_n675_), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT114), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n751_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n750_), .A2(G85gat), .A3(new_n368_), .A4(new_n752_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n723_), .A2(new_n668_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(G85gat), .B1(new_n755_), .B2(new_n368_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT112), .Z(new_n757_));
  AND2_X1   g556(.A1(new_n753_), .A2(new_n757_), .ZN(G1336gat));
  AND3_X1   g557(.A1(new_n632_), .A2(new_n443_), .A3(new_n444_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n750_), .A2(new_n752_), .A3(new_n759_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n203_), .B1(new_n754_), .B2(new_n692_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1337gat));
  OR3_X1    g561(.A1(new_n754_), .A2(new_n326_), .A3(new_n438_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n747_), .A2(new_n748_), .A3(new_n326_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n763_), .B1(new_n764_), .B2(new_n453_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(KEYINPUT51), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT51), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n767_), .B(new_n763_), .C1(new_n764_), .C2(new_n453_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(G1338gat));
  NAND3_X1  g568(.A1(new_n755_), .A2(new_n454_), .A3(new_n391_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n676_), .A2(new_n391_), .A3(new_n746_), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772_));
  AND3_X1   g571(.A1(new_n771_), .A2(new_n772_), .A3(G106gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n772_), .B1(new_n771_), .B2(G106gat), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n770_), .B1(new_n773_), .B2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT53), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n770_), .B(new_n777_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1339gat));
  NAND3_X1  g578(.A1(new_n610_), .A2(new_n505_), .A3(new_n567_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n780_), .B(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT58), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT55), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n497_), .A2(KEYINPUT116), .A3(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n482_), .A2(new_n476_), .A3(new_n484_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789_));
  OAI21_X1  g588(.A(KEYINPUT55), .B1(new_n485_), .B2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n791_), .A2(KEYINPUT56), .A3(new_n492_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT56), .B1(new_n791_), .B2(new_n492_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n497_), .A2(new_n478_), .A3(new_n491_), .A4(new_n480_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n510_), .B1(new_n543_), .B2(new_n549_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n552_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n798_));
  OAI211_X1 g597(.A(new_n509_), .B(new_n797_), .C1(new_n798_), .C2(new_n510_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n562_), .A2(new_n796_), .A3(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n785_), .B1(new_n795_), .B2(new_n802_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n800_), .B(KEYINPUT119), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n804_), .B(KEYINPUT58), .C1(new_n793_), .C2(new_n794_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n803_), .A2(new_n805_), .A3(new_n595_), .ZN(new_n806_));
  OR2_X1    g605(.A1(new_n806_), .A2(KEYINPUT120), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT57), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n792_), .A2(KEYINPUT118), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT118), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n790_), .A2(new_n788_), .ZN(new_n811_));
  NOR3_X1   g610(.A1(new_n485_), .A2(new_n789_), .A3(KEYINPUT55), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n810_), .B(new_n492_), .C1(new_n811_), .C2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n814_), .A2(KEYINPUT56), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n813_), .A2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n815_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n791_), .A2(new_n810_), .A3(new_n492_), .A4(new_n817_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n809_), .A2(new_n816_), .A3(new_n818_), .ZN(new_n819_));
  AND3_X1   g618(.A1(new_n563_), .A2(new_n565_), .A3(new_n796_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n562_), .A2(new_n799_), .ZN(new_n821_));
  AOI22_X1  g620(.A1(new_n819_), .A2(new_n820_), .B1(new_n502_), .B2(new_n821_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n808_), .B1(new_n822_), .B2(new_n594_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n819_), .A2(new_n820_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n502_), .A2(new_n821_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n594_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT57), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n806_), .A2(KEYINPUT120), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n807_), .A2(new_n823_), .A3(new_n827_), .A4(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n609_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n784_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n692_), .A2(new_n368_), .ZN(new_n832_));
  NOR3_X1   g631(.A1(new_n832_), .A2(new_n326_), .A3(new_n391_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(G113gat), .B1(new_n835_), .B2(new_n619_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n837_), .B(new_n806_), .C1(new_n826_), .C2(KEYINPUT57), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n827_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n837_), .B1(new_n823_), .B2(new_n806_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n609_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT122), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n843_), .B(new_n609_), .C1(new_n839_), .C2(new_n840_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n842_), .A2(new_n784_), .A3(new_n844_), .ZN(new_n845_));
  NOR4_X1   g644(.A1(new_n832_), .A2(KEYINPUT59), .A3(new_n326_), .A4(new_n391_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n845_), .A2(new_n846_), .B1(new_n834_), .B2(KEYINPUT59), .ZN(new_n847_));
  INV_X1    g646(.A(G113gat), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n567_), .A2(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n836_), .B1(new_n847_), .B2(new_n849_), .ZN(G1340gat));
  INV_X1    g649(.A(KEYINPUT60), .ZN(new_n851_));
  AOI21_X1  g650(.A(G120gat), .B1(new_n506_), .B2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n851_), .B2(G120gat), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n835_), .A2(new_n853_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(new_n854_), .B(KEYINPUT123), .ZN(new_n855_));
  INV_X1    g654(.A(G120gat), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n847_), .A2(new_n506_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(G1341gat));
  AOI21_X1  g657(.A(G127gat), .B1(new_n835_), .B2(new_n666_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n666_), .A2(G127gat), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n859_), .B1(new_n847_), .B2(new_n860_), .ZN(G1342gat));
  AOI21_X1  g660(.A(G134gat), .B1(new_n835_), .B2(new_n616_), .ZN(new_n862_));
  AND2_X1   g661(.A1(new_n595_), .A2(G134gat), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n847_), .B2(new_n863_), .ZN(G1343gat));
  AOI21_X1  g663(.A(new_n733_), .B1(new_n784_), .B2(new_n830_), .ZN(new_n865_));
  AND4_X1   g664(.A1(new_n368_), .A2(new_n865_), .A3(new_n391_), .A4(new_n692_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n619_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n506_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g669(.A1(new_n866_), .A2(new_n666_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(KEYINPUT61), .B(G155gat), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n871_), .B(new_n872_), .ZN(G1346gat));
  AOI21_X1  g672(.A(G162gat), .B1(new_n866_), .B2(new_n616_), .ZN(new_n874_));
  INV_X1    g673(.A(G162gat), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n671_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n866_), .B2(new_n876_), .ZN(G1347gat));
  NOR2_X1   g676(.A1(new_n326_), .A2(new_n368_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n632_), .A2(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n659_), .A2(new_n566_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n783_), .B1(new_n841_), .B2(KEYINPUT122), .ZN(new_n882_));
  AOI211_X1 g681(.A(new_n879_), .B(new_n881_), .C1(new_n882_), .C2(new_n844_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n233_), .ZN(new_n884_));
  OAI21_X1  g683(.A(KEYINPUT62), .B1(new_n883_), .B2(new_n211_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n879_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n845_), .A2(new_n886_), .A3(new_n880_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT124), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .A4(G169gat), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n885_), .A2(new_n890_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n879_), .B1(new_n882_), .B2(new_n844_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n211_), .B1(new_n892_), .B2(new_n880_), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n888_), .B1(new_n893_), .B2(new_n889_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n884_), .B1(new_n891_), .B2(new_n894_), .ZN(G1348gat));
  NAND3_X1  g694(.A1(new_n831_), .A2(new_n397_), .A3(new_n886_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n896_), .A2(new_n212_), .A3(new_n505_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n892_), .A2(new_n658_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n506_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n899_), .B2(new_n212_), .ZN(G1349gat));
  AND3_X1   g699(.A1(new_n666_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n892_), .A2(new_n658_), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(G183gat), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n903_), .B1(new_n896_), .B2(new_n609_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(new_n905_));
  XNOR2_X1  g704(.A(new_n905_), .B(KEYINPUT125), .ZN(G1350gat));
  NAND2_X1  g705(.A1(new_n898_), .A2(new_n595_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G190gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n898_), .A2(new_n223_), .A3(new_n616_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1351gat));
  AND4_X1   g709(.A1(new_n326_), .A2(new_n831_), .A3(new_n415_), .A4(new_n632_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(new_n619_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT126), .A2(G197gat), .ZN(new_n915_));
  XNOR2_X1  g714(.A(new_n914_), .B(new_n915_), .ZN(G1352gat));
  NAND2_X1  g715(.A1(new_n911_), .A2(new_n506_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g717(.A1(new_n911_), .A2(new_n666_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  AND2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  NOR3_X1   g720(.A1(new_n919_), .A2(new_n920_), .A3(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n922_), .B1(new_n919_), .B2(new_n920_), .ZN(G1354gat));
  NAND2_X1  g722(.A1(new_n911_), .A2(new_n616_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(KEYINPUT127), .B(G218gat), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n673_), .A2(new_n925_), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n924_), .A2(new_n925_), .B1(new_n911_), .B2(new_n926_), .ZN(G1355gat));
endmodule


