//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n837_, new_n839_,
    new_n840_, new_n841_, new_n842_, new_n843_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_;
  XNOR2_X1  g000(.A(KEYINPUT74), .B(G15gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G22gat), .ZN(new_n203_));
  INV_X1    g002(.A(G1gat), .ZN(new_n204_));
  INV_X1    g003(.A(G8gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  XOR2_X1   g006(.A(G1gat), .B(G8gat), .Z(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G231gat), .A2(G233gat), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n209_), .B(new_n210_), .Z(new_n211_));
  XNOR2_X1  g010(.A(KEYINPUT67), .B(G71gat), .ZN(new_n212_));
  INV_X1    g011(.A(G78gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G57gat), .B(G64gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n215_), .B(KEYINPUT11), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n215_), .A2(KEYINPUT11), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n217_), .B1(new_n219_), .B2(new_n214_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n211_), .B(new_n220_), .ZN(new_n221_));
  XNOR2_X1  g020(.A(G127gat), .B(G155gat), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n222_), .B(KEYINPUT16), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n223_), .B(G183gat), .ZN(new_n224_));
  INV_X1    g023(.A(G211gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(new_n224_), .B(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT17), .ZN(new_n227_));
  NOR2_X1   g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n221_), .A2(KEYINPUT75), .A3(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT75), .B1(new_n221_), .B2(new_n228_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n226_), .B(new_n227_), .ZN(new_n231_));
  OAI22_X1  g030(.A1(new_n229_), .A2(new_n230_), .B1(new_n221_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  AOI211_X1 g032(.A(G99gat), .B(G106gat), .C1(KEYINPUT65), .C2(KEYINPUT7), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n234_), .B1(KEYINPUT65), .B2(KEYINPUT7), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT64), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G99gat), .A2(G106gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT6), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n235_), .A2(new_n238_), .A3(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G85gat), .B(G92gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n241_), .A2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT8), .ZN(new_n246_));
  INV_X1    g045(.A(new_n242_), .ZN(new_n247_));
  XOR2_X1   g046(.A(KEYINPUT10), .B(G99gat), .Z(new_n248_));
  INV_X1    g047(.A(G106gat), .ZN(new_n249_));
  AOI22_X1  g048(.A1(new_n247_), .A2(KEYINPUT9), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G85gat), .A2(G92gat), .ZN(new_n251_));
  OAI211_X1 g050(.A(new_n250_), .B(new_n240_), .C1(KEYINPUT9), .C2(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n246_), .A2(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n253_), .A2(new_n220_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n220_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n254_), .A2(KEYINPUT68), .A3(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n255_), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT68), .B1(new_n253_), .B2(new_n220_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AND2_X1   g058(.A1(G230gat), .A2(G233gat), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n256_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT12), .B1(new_n253_), .B2(new_n220_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(new_n262_), .B(new_n255_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n261_), .B1(new_n263_), .B2(new_n260_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G120gat), .B(G148gat), .ZN(new_n265_));
  INV_X1    g064(.A(G204gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT5), .B(G176gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(new_n268_), .Z(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n264_), .A2(new_n270_), .ZN(new_n271_));
  OAI211_X1 g070(.A(new_n261_), .B(new_n269_), .C1(new_n263_), .C2(new_n260_), .ZN(new_n272_));
  AND3_X1   g071(.A1(new_n271_), .A2(KEYINPUT13), .A3(new_n272_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT13), .B1(new_n271_), .B2(new_n272_), .ZN(new_n274_));
  NOR2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT76), .ZN(new_n277_));
  INV_X1    g076(.A(new_n209_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G43gat), .B(G50gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G29gat), .B(G36gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n277_), .B1(new_n278_), .B2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n209_), .A2(KEYINPUT76), .A3(new_n283_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n283_), .B(KEYINPUT15), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n278_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(G229gat), .A2(G233gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n287_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G113gat), .B(G141gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(G197gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT77), .B(G169gat), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n293_), .B(new_n294_), .Z(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AOI22_X1  g095(.A1(new_n285_), .A2(new_n286_), .B1(new_n278_), .B2(new_n284_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n291_), .B(new_n296_), .C1(new_n297_), .C2(new_n290_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT78), .ZN(new_n299_));
  OR2_X1    g098(.A1(new_n297_), .A2(new_n290_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT78), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n300_), .A2(new_n301_), .A3(new_n291_), .A4(new_n296_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n299_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n291_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n295_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n303_), .A2(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n276_), .A2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G225gat), .A2(G233gat), .ZN(new_n309_));
  XOR2_X1   g108(.A(G141gat), .B(G148gat), .Z(new_n310_));
  NAND2_X1  g109(.A1(G155gat), .A2(G162gat), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT83), .ZN(new_n312_));
  AND3_X1   g111(.A1(new_n311_), .A2(new_n312_), .A3(KEYINPUT1), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n312_), .B1(new_n311_), .B2(KEYINPUT1), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT84), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n316_), .B1(new_n311_), .B2(KEYINPUT1), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT82), .ZN(new_n318_));
  INV_X1    g117(.A(G155gat), .ZN(new_n319_));
  INV_X1    g118(.A(G162gat), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n318_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT1), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n323_), .A2(KEYINPUT84), .A3(G155gat), .A4(G162gat), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n317_), .A2(new_n321_), .A3(new_n322_), .A4(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n310_), .B1(new_n315_), .B2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G141gat), .A2(G148gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT85), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(KEYINPUT2), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT2), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n327_), .A2(KEYINPUT85), .A3(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n332_));
  OR3_X1    g131(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n329_), .A2(new_n331_), .A3(new_n332_), .A4(new_n333_), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n321_), .A2(new_n311_), .A3(new_n322_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n326_), .A2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G127gat), .B(G134gat), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G113gat), .B(G120gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n337_), .B(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n341_), .A2(KEYINPUT4), .ZN(new_n342_));
  INV_X1    g141(.A(new_n337_), .ZN(new_n343_));
  OR3_X1    g142(.A1(new_n343_), .A2(KEYINPUT4), .A3(new_n340_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n309_), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT0), .ZN(new_n347_));
  INV_X1    g146(.A(G57gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(G85gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n349_), .B(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n309_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n341_), .A2(new_n353_), .ZN(new_n354_));
  OR3_X1    g153(.A1(new_n345_), .A2(new_n352_), .A3(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n352_), .B1(new_n345_), .B2(new_n354_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT87), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT29), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n326_), .A2(new_n360_), .A3(new_n336_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n361_), .A2(KEYINPUT86), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G22gat), .B(G50gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n363_), .B(KEYINPUT28), .Z(new_n364_));
  INV_X1    g163(.A(KEYINPUT86), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n326_), .A2(new_n336_), .A3(new_n365_), .A4(new_n360_), .ZN(new_n366_));
  AND3_X1   g165(.A1(new_n362_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n364_), .B1(new_n362_), .B2(new_n366_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n359_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n362_), .A2(new_n366_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n364_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n362_), .A2(new_n364_), .A3(new_n366_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n372_), .A2(KEYINPUT87), .A3(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G78gat), .B(G106gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(G228gat), .A2(G233gat), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n376_), .A2(KEYINPUT91), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n375_), .B(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(G218gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G211gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n225_), .A2(G218gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT21), .ZN(new_n383_));
  AND2_X1   g182(.A1(G197gat), .A2(G204gat), .ZN(new_n384_));
  NOR2_X1   g183(.A1(G197gat), .A2(G204gat), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n386_), .A2(KEYINPUT90), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n386_), .A2(KEYINPUT90), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n383_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT88), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n386_), .B2(KEYINPUT21), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT21), .ZN(new_n393_));
  OAI211_X1 g192(.A(KEYINPUT88), .B(new_n393_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n382_), .B1(KEYINPUT21), .B2(new_n386_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n395_), .A2(KEYINPUT89), .A3(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT89), .B1(new_n395_), .B2(new_n396_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n390_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n360_), .B1(new_n326_), .B2(new_n336_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n399_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n376_), .A2(KEYINPUT91), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n378_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G197gat), .B(G204gat), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT88), .B1(new_n405_), .B2(new_n393_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n394_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n396_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT89), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n395_), .A2(KEYINPUT89), .A3(new_n396_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n389_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n403_), .B(new_n378_), .C1(new_n412_), .C2(new_n400_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n369_), .B(new_n374_), .C1(new_n404_), .C2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT92), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n403_), .B1(new_n412_), .B2(new_n400_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n378_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n413_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n421_), .A2(KEYINPUT92), .A3(new_n374_), .A4(new_n369_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n372_), .A2(new_n373_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n423_), .A2(new_n420_), .A3(new_n413_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  AND4_X1   g224(.A1(KEYINPUT93), .A2(new_n417_), .A3(new_n422_), .A4(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n424_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n427_));
  AOI21_X1  g226(.A(KEYINPUT93), .B1(new_n427_), .B2(new_n422_), .ZN(new_n428_));
  OAI21_X1  g227(.A(new_n358_), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G8gat), .B(G36gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(KEYINPUT18), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(G64gat), .ZN(new_n432_));
  INV_X1    g231(.A(G92gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G169gat), .A2(G176gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n436_), .B(KEYINPUT79), .ZN(new_n437_));
  NOR2_X1   g236(.A1(G169gat), .A2(G176gat), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n437_), .A2(KEYINPUT24), .A3(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(KEYINPUT25), .B(G183gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(KEYINPUT26), .B(G190gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(G183gat), .A2(G190gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(KEYINPUT23), .ZN(new_n445_));
  INV_X1    g244(.A(KEYINPUT23), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(G183gat), .A3(G190gat), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT24), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n445_), .A2(new_n447_), .B1(new_n448_), .B2(new_n438_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n443_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(G169gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(KEYINPUT22), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT22), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(G169gat), .ZN(new_n454_));
  INV_X1    g253(.A(G176gat), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n452_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n437_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT80), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n445_), .A2(new_n447_), .A3(new_n458_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n446_), .A2(KEYINPUT80), .A3(G183gat), .A4(G190gat), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n459_), .B(new_n460_), .C1(G183gat), .C2(G190gat), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n440_), .A2(new_n450_), .B1(new_n457_), .B2(new_n461_), .ZN(new_n462_));
  OAI211_X1 g261(.A(new_n462_), .B(new_n390_), .C1(new_n397_), .C2(new_n398_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n448_), .A2(KEYINPUT94), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n448_), .A2(KEYINPUT94), .ZN(new_n465_));
  OR3_X1    g264(.A1(new_n464_), .A2(new_n439_), .A3(new_n465_), .ZN(new_n466_));
  OAI211_X1 g265(.A(new_n436_), .B(new_n439_), .C1(new_n464_), .C2(new_n465_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n466_), .A2(new_n443_), .A3(new_n467_), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n459_), .A2(new_n460_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n445_), .A2(new_n447_), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n470_), .B1(G183gat), .B2(G190gat), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n468_), .A2(new_n469_), .B1(new_n457_), .B2(new_n471_), .ZN(new_n472_));
  OAI211_X1 g271(.A(new_n463_), .B(KEYINPUT20), .C1(new_n412_), .C2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G226gat), .A2(G233gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n474_), .B(KEYINPUT19), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n475_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n478_), .B1(new_n412_), .B2(new_n472_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n462_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n399_), .A2(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n477_), .B1(new_n479_), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n435_), .B1(new_n476_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n473_), .A2(new_n475_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT95), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n479_), .A2(new_n477_), .A3(new_n481_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n484_), .A2(new_n485_), .A3(new_n434_), .A4(new_n486_), .ZN(new_n487_));
  AND3_X1   g286(.A1(new_n483_), .A2(KEYINPUT27), .A3(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n484_), .A2(new_n434_), .A3(new_n486_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT95), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT96), .ZN(new_n492_));
  INV_X1    g291(.A(new_n486_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n468_), .A2(new_n469_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n457_), .A2(new_n471_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  AOI21_X1  g295(.A(new_n478_), .B1(new_n399_), .B2(new_n496_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n477_), .B1(new_n497_), .B2(new_n463_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n435_), .B1(new_n493_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n489_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT27), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n492_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  AOI211_X1 g301(.A(KEYINPUT96), .B(KEYINPUT27), .C1(new_n499_), .C2(new_n489_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n491_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT97), .B1(new_n429_), .B2(new_n504_), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n484_), .A2(new_n434_), .A3(new_n486_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n434_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n501_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT96), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n500_), .A2(new_n492_), .A3(new_n501_), .ZN(new_n510_));
  AOI22_X1  g309(.A1(new_n509_), .A2(new_n510_), .B1(new_n490_), .B2(new_n488_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n417_), .A2(new_n422_), .A3(new_n425_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT93), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n427_), .A2(KEYINPUT93), .A3(new_n422_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT97), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n511_), .A2(new_n516_), .A3(new_n517_), .A4(new_n358_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n516_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT33), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n356_), .B(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n342_), .A2(new_n309_), .A3(new_n344_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n341_), .A2(new_n353_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n351_), .A3(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n499_), .A2(new_n489_), .A3(new_n524_), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n434_), .A2(KEYINPUT32), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n526_), .B1(new_n476_), .B2(new_n482_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n484_), .A2(new_n486_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n527_), .B1(new_n528_), .B2(new_n526_), .ZN(new_n529_));
  OAI22_X1  g328(.A1(new_n521_), .A2(new_n525_), .B1(new_n358_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n519_), .A2(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n505_), .A2(new_n518_), .A3(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT98), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n462_), .B(KEYINPUT30), .ZN(new_n534_));
  XOR2_X1   g333(.A(G71gat), .B(G99gat), .Z(new_n535_));
  NAND2_X1  g334(.A1(G227gat), .A2(G233gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n535_), .B(new_n536_), .Z(new_n537_));
  XNOR2_X1  g336(.A(new_n534_), .B(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT81), .B(KEYINPUT31), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(new_n539_), .ZN(new_n540_));
  XOR2_X1   g339(.A(G15gat), .B(G43gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n340_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n540_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n540_), .A2(new_n543_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  AND3_X1   g346(.A1(new_n532_), .A2(new_n533_), .A3(new_n547_), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n533_), .B1(new_n532_), .B2(new_n547_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n519_), .A2(new_n511_), .ZN(new_n550_));
  NOR3_X1   g349(.A1(new_n550_), .A2(new_n547_), .A3(new_n357_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n548_), .A2(new_n549_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n288_), .A2(new_n253_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT71), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n288_), .A2(KEYINPUT71), .A3(new_n253_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT34), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT35), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n246_), .A2(new_n252_), .ZN(new_n564_));
  AOI22_X1  g363(.A1(new_n564_), .A2(new_n283_), .B1(new_n561_), .B2(new_n560_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n557_), .A2(new_n563_), .A3(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(new_n563_), .B1(new_n557_), .B2(new_n565_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT73), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n568_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT73), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n570_), .A2(new_n571_), .A3(new_n566_), .ZN(new_n572_));
  XOR2_X1   g371(.A(G190gat), .B(G218gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(G134gat), .B(G162gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT36), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n569_), .A2(new_n572_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT36), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n575_), .A2(new_n578_), .ZN(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT72), .Z(new_n580_));
  OR3_X1    g379(.A1(new_n567_), .A2(new_n568_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n577_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NOR3_X1   g382(.A1(new_n552_), .A2(KEYINPUT102), .A3(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT102), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n532_), .A2(new_n547_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT98), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n532_), .A2(new_n533_), .A3(new_n547_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n551_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n585_), .B1(new_n590_), .B2(new_n582_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n233_), .B(new_n308_), .C1(new_n584_), .C2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT103), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n593_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n357_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(G1gat), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT99), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n590_), .A2(new_n598_), .A3(new_n306_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n598_), .B1(new_n590_), .B2(new_n306_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT37), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n582_), .A2(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n576_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n581_), .A2(KEYINPUT37), .A3(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n604_), .A2(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n273_), .A2(new_n274_), .A3(new_n232_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n602_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT100), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT100), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n602_), .B2(new_n609_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n358_), .A2(G1gat), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n611_), .A2(new_n613_), .A3(new_n614_), .ZN(new_n615_));
  NAND4_X1  g414(.A1(new_n611_), .A2(KEYINPUT38), .A3(new_n613_), .A4(new_n614_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n616_), .A2(new_n617_), .ZN(new_n619_));
  OAI221_X1 g418(.A(new_n597_), .B1(KEYINPUT38), .B2(new_n615_), .C1(new_n618_), .C2(new_n619_), .ZN(G1324gat));
  NAND4_X1  g419(.A1(new_n611_), .A2(new_n205_), .A3(new_n504_), .A4(new_n613_), .ZN(new_n621_));
  OAI21_X1  g420(.A(G8gat), .B1(new_n592_), .B2(new_n511_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n622_), .A2(KEYINPUT39), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n622_), .A2(KEYINPUT39), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n621_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT40), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  OAI211_X1 g426(.A(new_n621_), .B(KEYINPUT40), .C1(new_n623_), .C2(new_n624_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1325gat));
  NAND3_X1  g428(.A1(new_n594_), .A2(new_n546_), .A3(new_n595_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(G15gat), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n631_), .A2(KEYINPUT41), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(KEYINPUT41), .ZN(new_n633_));
  NOR4_X1   g432(.A1(new_n602_), .A2(G15gat), .A3(new_n547_), .A4(new_n609_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT104), .Z(new_n635_));
  NAND3_X1  g434(.A1(new_n632_), .A2(new_n633_), .A3(new_n635_), .ZN(G1326gat));
  INV_X1    g435(.A(G22gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n610_), .A2(new_n637_), .A3(new_n516_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n594_), .A2(new_n516_), .A3(new_n595_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT42), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n639_), .A2(new_n640_), .A3(G22gat), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n639_), .B2(G22gat), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n638_), .B1(new_n641_), .B2(new_n642_), .ZN(G1327gat));
  NOR3_X1   g442(.A1(new_n276_), .A2(new_n582_), .A3(new_n233_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(KEYINPUT99), .B1(new_n552_), .B2(new_n307_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n645_), .B1(new_n646_), .B2(new_n599_), .ZN(new_n647_));
  AOI21_X1  g446(.A(G29gat), .B1(new_n647_), .B2(new_n357_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n551_), .B1(new_n586_), .B2(KEYINPUT98), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n607_), .B1(new_n649_), .B2(new_n588_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT43), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT105), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT105), .ZN(new_n653_));
  OAI211_X1 g452(.A(new_n653_), .B(KEYINPUT43), .C1(new_n552_), .C2(new_n607_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n607_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n590_), .A2(new_n651_), .A3(new_n655_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n652_), .A2(new_n654_), .A3(new_n656_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n276_), .A2(new_n307_), .A3(new_n233_), .ZN(new_n658_));
  AOI21_X1  g457(.A(KEYINPUT44), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(G29gat), .A3(new_n357_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n651_), .B1(new_n590_), .B2(new_n655_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n656_), .B1(new_n662_), .B2(new_n653_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n650_), .A2(KEYINPUT105), .A3(new_n651_), .ZN(new_n664_));
  OAI211_X1 g463(.A(KEYINPUT44), .B(new_n658_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT106), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n657_), .A2(new_n667_), .A3(KEYINPUT44), .A4(new_n658_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n648_), .B1(new_n661_), .B2(new_n669_), .ZN(G1328gat));
  INV_X1    g469(.A(KEYINPUT108), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n671_), .A2(KEYINPUT46), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n511_), .A2(G36gat), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n644_), .B(new_n674_), .C1(new_n600_), .C2(new_n601_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(KEYINPUT107), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n647_), .A2(new_n677_), .A3(new_n674_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n676_), .A2(KEYINPUT45), .A3(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  AOI21_X1  g479(.A(KEYINPUT45), .B1(new_n676_), .B2(new_n678_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  AOI211_X1 g481(.A(new_n511_), .B(new_n659_), .C1(new_n666_), .C2(new_n668_), .ZN(new_n683_));
  INV_X1    g482(.A(G36gat), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n673_), .B(new_n682_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n659_), .A2(new_n511_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n684_), .B1(new_n669_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n676_), .A2(new_n678_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT45), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n690_), .A2(new_n679_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n672_), .B1(new_n687_), .B2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n685_), .A2(new_n692_), .ZN(G1329gat));
  NAND2_X1  g492(.A1(new_n546_), .A2(G43gat), .ZN(new_n694_));
  AOI211_X1 g493(.A(new_n659_), .B(new_n694_), .C1(new_n666_), .C2(new_n668_), .ZN(new_n695_));
  AOI21_X1  g494(.A(G43gat), .B1(new_n647_), .B2(new_n546_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT47), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NAND4_X1  g496(.A1(new_n669_), .A2(G43gat), .A3(new_n546_), .A4(new_n660_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT47), .ZN(new_n699_));
  INV_X1    g498(.A(new_n696_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n697_), .A2(new_n701_), .ZN(G1330gat));
  AOI21_X1  g501(.A(G50gat), .B1(new_n647_), .B2(new_n516_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n660_), .A2(G50gat), .A3(new_n516_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n704_), .B2(new_n669_), .ZN(G1331gat));
  NOR2_X1   g504(.A1(new_n584_), .A2(new_n591_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n275_), .A2(new_n306_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n233_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n358_), .A2(new_n348_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(KEYINPUT109), .B2(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(G57gat), .B1(new_n711_), .B2(KEYINPUT109), .ZN(new_n712_));
  NOR3_X1   g511(.A1(new_n552_), .A2(new_n655_), .A3(new_n708_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n711_), .A2(new_n357_), .A3(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT110), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n715_), .B(new_n716_), .ZN(G1332gat));
  INV_X1    g516(.A(G64gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n709_), .B2(new_n504_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT48), .Z(new_n720_));
  NAND3_X1  g519(.A1(new_n713_), .A2(new_n718_), .A3(new_n504_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1333gat));
  INV_X1    g521(.A(G71gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n709_), .B2(new_n546_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT49), .Z(new_n725_));
  NAND2_X1  g524(.A1(new_n546_), .A2(new_n723_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT111), .Z(new_n727_));
  NAND2_X1  g526(.A1(new_n713_), .A2(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n725_), .A2(new_n728_), .ZN(G1334gat));
  NAND3_X1  g528(.A1(new_n713_), .A2(new_n213_), .A3(new_n516_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n708_), .ZN(new_n731_));
  OAI211_X1 g530(.A(new_n516_), .B(new_n731_), .C1(new_n584_), .C2(new_n591_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n733_));
  AND3_X1   g532(.A1(new_n732_), .A2(new_n733_), .A3(G78gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n732_), .B2(G78gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n730_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT112), .ZN(G1335gat));
  NAND2_X1  g536(.A1(new_n707_), .A2(new_n232_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n657_), .A2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G85gat), .B1(new_n740_), .B2(new_n358_), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n552_), .A2(new_n582_), .A3(new_n738_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(new_n350_), .A3(new_n357_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1336gat));
  OAI21_X1  g543(.A(G92gat), .B1(new_n740_), .B2(new_n511_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n742_), .A2(new_n433_), .A3(new_n504_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1337gat));
  OAI21_X1  g546(.A(G99gat), .B1(new_n740_), .B2(new_n547_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n742_), .A2(new_n546_), .A3(new_n248_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT113), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g551(.A1(new_n742_), .A2(new_n249_), .A3(new_n516_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n657_), .A2(new_n516_), .A3(new_n739_), .ZN(new_n754_));
  XOR2_X1   g553(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n755_));
  AND3_X1   g554(.A1(new_n754_), .A2(G106gat), .A3(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n755_), .B1(new_n754_), .B2(G106gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  XOR2_X1   g557(.A(KEYINPUT115), .B(KEYINPUT53), .Z(new_n759_));
  XNOR2_X1  g558(.A(new_n758_), .B(new_n759_), .ZN(G1339gat));
  NAND4_X1  g559(.A1(new_n604_), .A2(new_n608_), .A3(new_n307_), .A4(new_n606_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT116), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n761_), .A2(new_n762_), .A3(KEYINPUT54), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n761_), .B2(KEYINPUT54), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n761_), .A2(KEYINPUT54), .ZN(new_n765_));
  NOR3_X1   g564(.A1(new_n763_), .A2(new_n764_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT120), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n254_), .A2(KEYINPUT12), .A3(new_n255_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n257_), .A2(new_n262_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n260_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n770_));
  OAI21_X1  g569(.A(KEYINPUT55), .B1(new_n770_), .B2(KEYINPUT117), .ZN(new_n771_));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772_));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n772_), .B(new_n773_), .C1(new_n263_), .C2(new_n260_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n263_), .A2(new_n260_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n771_), .A2(new_n774_), .A3(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(new_n270_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT56), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n776_), .A2(KEYINPUT56), .A3(new_n270_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(KEYINPUT119), .A3(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT119), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n776_), .A2(new_n782_), .A3(KEYINPUT56), .A4(new_n270_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n290_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n287_), .A2(new_n289_), .A3(new_n784_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n295_), .C1(new_n297_), .C2(new_n784_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n303_), .A2(new_n272_), .A3(new_n786_), .ZN(new_n787_));
  AND2_X1   g586(.A1(new_n783_), .A2(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT58), .B1(new_n781_), .B2(new_n788_), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n789_), .A2(new_n607_), .ZN(new_n790_));
  AND3_X1   g589(.A1(new_n781_), .A2(new_n788_), .A3(KEYINPUT58), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n767_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n791_), .A2(new_n789_), .A3(new_n607_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(KEYINPUT120), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n306_), .A2(new_n272_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n795_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n303_), .A2(new_n786_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n797_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n582_), .B1(new_n796_), .B2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(KEYINPUT118), .A2(KEYINPUT57), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI221_X1 g600(.A(new_n582_), .B1(KEYINPUT118), .B2(KEYINPUT57), .C1(new_n796_), .C2(new_n798_), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n792_), .A2(new_n794_), .A3(new_n801_), .A4(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n766_), .B1(new_n803_), .B2(new_n232_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n550_), .A2(new_n547_), .A3(new_n358_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT59), .B1(new_n804_), .B2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n801_), .A2(new_n802_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n232_), .B1(new_n809_), .B2(new_n793_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT122), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n766_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT122), .B(new_n232_), .C1(new_n809_), .C2(new_n793_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n805_), .B(new_n808_), .C1(new_n814_), .C2(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n807_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n306_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n819_), .A2(G113gat), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n804_), .A2(new_n806_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  OR3_X1    g621(.A1(new_n822_), .A2(G113gat), .A3(new_n307_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n823_), .ZN(G1340gat));
  INV_X1    g623(.A(KEYINPUT60), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n275_), .B2(G120gat), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n821_), .A2(new_n826_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n827_), .A2(new_n807_), .A3(new_n276_), .A4(new_n817_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(G120gat), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n829_), .B1(KEYINPUT60), .B2(new_n827_), .ZN(G1341gat));
  NAND2_X1  g629(.A1(new_n818_), .A2(new_n233_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(G127gat), .ZN(new_n832_));
  OR3_X1    g631(.A1(new_n822_), .A2(G127gat), .A3(new_n232_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1342gat));
  NAND2_X1  g633(.A1(new_n818_), .A2(new_n655_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G134gat), .ZN(new_n836_));
  OR3_X1    g635(.A1(new_n822_), .A2(G134gat), .A3(new_n582_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(G1343gat));
  INV_X1    g637(.A(new_n804_), .ZN(new_n839_));
  NOR4_X1   g638(.A1(new_n519_), .A2(new_n546_), .A3(new_n504_), .A4(new_n358_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n841_), .A2(new_n307_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(KEYINPUT123), .B(G141gat), .ZN(new_n843_));
  XNOR2_X1  g642(.A(new_n842_), .B(new_n843_), .ZN(G1344gat));
  NAND3_X1  g643(.A1(new_n839_), .A2(new_n276_), .A3(new_n840_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g645(.A1(new_n841_), .A2(new_n232_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(KEYINPUT61), .B(G155gat), .ZN(new_n848_));
  XNOR2_X1  g647(.A(new_n848_), .B(KEYINPUT124), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n847_), .B(new_n849_), .ZN(G1346gat));
  NOR3_X1   g649(.A1(new_n841_), .A2(new_n320_), .A3(new_n607_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n320_), .B1(new_n841_), .B2(new_n582_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT125), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT125), .B(new_n320_), .C1(new_n841_), .C2(new_n582_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n851_), .B1(new_n854_), .B2(new_n855_), .ZN(G1347gat));
  NOR2_X1   g655(.A1(new_n547_), .A2(new_n357_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n504_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n519_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n766_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n861_), .B2(new_n815_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n451_), .B1(new_n862_), .B2(new_n306_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n306_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n452_), .A2(new_n454_), .ZN(new_n865_));
  OAI22_X1  g664(.A1(new_n863_), .A2(KEYINPUT62), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  AOI211_X1 g666(.A(new_n867_), .B(new_n451_), .C1(new_n862_), .C2(new_n306_), .ZN(new_n868_));
  OAI21_X1  g667(.A(KEYINPUT126), .B1(new_n866_), .B2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n864_), .A2(G169gat), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n867_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n864_), .A2(new_n865_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT126), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n863_), .A2(KEYINPUT62), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .A4(new_n874_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n869_), .A2(new_n875_), .ZN(G1348gat));
  AOI21_X1  g675(.A(G176gat), .B1(new_n862_), .B2(new_n276_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n804_), .A2(new_n516_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n858_), .A2(new_n455_), .A3(new_n275_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n877_), .B1(new_n878_), .B2(new_n879_), .ZN(G1349gat));
  NAND3_X1  g679(.A1(new_n878_), .A2(new_n233_), .A3(new_n859_), .ZN(new_n881_));
  INV_X1    g680(.A(G183gat), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n232_), .A2(new_n441_), .ZN(new_n883_));
  AOI22_X1  g682(.A1(new_n881_), .A2(new_n882_), .B1(new_n862_), .B2(new_n883_), .ZN(G1350gat));
  INV_X1    g683(.A(new_n862_), .ZN(new_n885_));
  OAI21_X1  g684(.A(G190gat), .B1(new_n885_), .B2(new_n607_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n862_), .A2(new_n442_), .A3(new_n583_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1351gat));
  INV_X1    g687(.A(KEYINPUT127), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n547_), .A2(new_n504_), .A3(new_n358_), .A4(new_n516_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n889_), .B1(new_n804_), .B2(new_n890_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n891_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n804_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n306_), .B1(new_n892_), .B2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(G197gat), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n804_), .A2(new_n890_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(KEYINPUT127), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n891_), .ZN(new_n898_));
  INV_X1    g697(.A(G197gat), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n898_), .A2(new_n899_), .A3(new_n306_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n895_), .A2(new_n900_), .ZN(G1352gat));
  AOI21_X1  g700(.A(G204gat), .B1(new_n898_), .B2(new_n276_), .ZN(new_n902_));
  AOI211_X1 g701(.A(new_n266_), .B(new_n275_), .C1(new_n897_), .C2(new_n891_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(G1353gat));
  OR2_X1    g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(new_n898_), .B2(new_n233_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT63), .B(G211gat), .ZN(new_n907_));
  AOI211_X1 g706(.A(new_n232_), .B(new_n907_), .C1(new_n897_), .C2(new_n891_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1354gat));
  NAND3_X1  g708(.A1(new_n898_), .A2(new_n379_), .A3(new_n583_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n607_), .B1(new_n897_), .B2(new_n891_), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n910_), .B1(new_n379_), .B2(new_n911_), .ZN(G1355gat));
endmodule


