//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n747_, new_n748_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n758_, new_n759_, new_n760_, new_n761_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n785_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n890_, new_n891_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n898_, new_n899_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n205_), .A3(KEYINPUT85), .ZN(new_n206_));
  OR3_X1    g005(.A1(new_n202_), .A2(KEYINPUT85), .A3(KEYINPUT23), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n206_), .A2(new_n207_), .A3(new_n209_), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(KEYINPUT86), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(KEYINPUT86), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(KEYINPUT84), .A2(G169gat), .ZN(new_n215_));
  AOI21_X1  g014(.A(G176gat), .B1(new_n215_), .B2(KEYINPUT22), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT22), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(KEYINPUT84), .A3(G169gat), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n214_), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n211_), .A2(new_n212_), .A3(new_n219_), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT25), .B(G183gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT83), .ZN(new_n222_));
  INV_X1    g021(.A(G190gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT26), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n223_), .A2(KEYINPUT26), .ZN(new_n225_));
  OAI211_X1 g024(.A(new_n221_), .B(new_n224_), .C1(new_n225_), .C2(new_n222_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n203_), .A2(new_n205_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(G169gat), .B2(G176gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n228_), .ZN(new_n233_));
  NAND4_X1  g032(.A1(new_n226_), .A2(new_n227_), .A3(new_n232_), .A4(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n220_), .A2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n235_), .B(KEYINPUT30), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT88), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(G227gat), .A2(G233gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n239_), .B(KEYINPUT87), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G15gat), .B(G43gat), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n240_), .B(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G71gat), .B(G99gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n238_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT31), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT31), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n238_), .A2(new_n247_), .A3(new_n244_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(G113gat), .B(G120gat), .Z(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT89), .ZN(new_n251_));
  XNOR2_X1  g050(.A(G113gat), .B(G120gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT89), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G127gat), .B(G134gat), .Z(new_n256_));
  OR2_X1    g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n251_), .A2(new_n254_), .A3(new_n256_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT90), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT91), .ZN(new_n260_));
  AND3_X1   g059(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n260_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n257_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n258_), .A2(new_n259_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(KEYINPUT91), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n255_), .A2(new_n256_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n258_), .A2(new_n259_), .A3(new_n260_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n265_), .A2(new_n266_), .A3(new_n267_), .ZN(new_n268_));
  AND2_X1   g067(.A1(new_n263_), .A2(new_n268_), .ZN(new_n269_));
  OR3_X1    g068(.A1(new_n236_), .A2(new_n237_), .A3(new_n269_), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n269_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n249_), .A2(new_n272_), .ZN(new_n273_));
  NAND4_X1  g072(.A1(new_n246_), .A2(new_n248_), .A3(new_n270_), .A4(new_n271_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  XOR2_X1   g074(.A(G1gat), .B(G29gat), .Z(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT101), .B(G85gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT0), .B(G57gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G155gat), .A2(G162gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n282_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT2), .ZN(new_n285_));
  INV_X1    g084(.A(G141gat), .ZN(new_n286_));
  INV_X1    g085(.A(G148gat), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n285_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT3), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n293_));
  NAND4_X1  g092(.A1(new_n288_), .A2(new_n291_), .A3(new_n292_), .A4(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n284_), .A2(KEYINPUT94), .A3(new_n294_), .A4(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n282_), .A2(new_n283_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT93), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(KEYINPUT92), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT92), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(KEYINPUT93), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n299_), .A2(new_n301_), .A3(new_n283_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n294_), .B(new_n295_), .C1(new_n297_), .C2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT94), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n296_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n295_), .B(KEYINPUT1), .Z(new_n307_));
  NAND2_X1  g106(.A1(new_n284_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(G141gat), .B(G148gat), .Z(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n306_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n263_), .A2(new_n311_), .A3(new_n268_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT4), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n257_), .A2(new_n258_), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n296_), .A2(new_n305_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n313_), .B1(new_n312_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G225gat), .A2(G233gat), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n315_), .A2(new_n319_), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n312_), .A2(new_n318_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n320_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n281_), .B1(new_n321_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT102), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n322_), .A2(KEYINPUT4), .ZN(new_n327_));
  INV_X1    g126(.A(new_n320_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n328_), .A3(new_n314_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(new_n280_), .A3(new_n323_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n325_), .A2(new_n326_), .A3(new_n330_), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n329_), .A2(KEYINPUT102), .A3(new_n280_), .A4(new_n323_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n275_), .A2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G197gat), .B(G204gat), .Z(new_n335_));
  NAND2_X1  g134(.A1(new_n335_), .A2(KEYINPUT21), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G211gat), .B(G218gat), .ZN(new_n337_));
  OR2_X1    g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G197gat), .B(G204gat), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT21), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n336_), .A2(new_n341_), .A3(new_n337_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n343_), .B1(new_n220_), .B2(new_n234_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n338_), .A2(new_n342_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(KEYINPUT22), .B(G169gat), .ZN(new_n347_));
  INV_X1    g146(.A(G176gat), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n214_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n227_), .A2(new_n209_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT26), .B(G190gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n221_), .A2(new_n352_), .ZN(new_n353_));
  NAND4_X1  g152(.A1(new_n353_), .A2(new_n206_), .A3(new_n207_), .A4(new_n233_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT98), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n231_), .B1(new_n229_), .B2(new_n355_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n214_), .A2(KEYINPUT98), .A3(new_n228_), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n351_), .B1(new_n354_), .B2(new_n358_), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT20), .B1(new_n346_), .B2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G226gat), .A2(G233gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n345_), .A2(new_n361_), .A3(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n220_), .A2(new_n343_), .A3(new_n234_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT20), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n346_), .B2(new_n359_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n364_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G8gat), .B(G36gat), .Z(new_n372_));
  XNOR2_X1  g171(.A(new_n372_), .B(KEYINPUT18), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G64gat), .B(G92gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n373_), .B(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n366_), .A2(new_n371_), .A3(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT99), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n366_), .A2(new_n371_), .A3(KEYINPUT99), .A4(new_n375_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT100), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n366_), .A2(new_n371_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n375_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n344_), .A2(new_n364_), .A3(new_n360_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n365_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n385_));
  OAI211_X1 g184(.A(new_n380_), .B(new_n382_), .C1(new_n384_), .C2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n378_), .B(new_n379_), .C1(new_n383_), .C2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT27), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n364_), .B1(new_n344_), .B2(new_n360_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n391_), .B1(new_n364_), .B2(new_n370_), .ZN(new_n392_));
  XOR2_X1   g191(.A(new_n375_), .B(KEYINPUT103), .Z(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(KEYINPUT27), .A3(new_n376_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT104), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n394_), .A2(KEYINPUT104), .A3(KEYINPUT27), .A4(new_n376_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n390_), .A2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G78gat), .B(G106gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT29), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n346_), .B1(new_n317_), .B2(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(G228gat), .A3(G233gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G228gat), .A2(G233gat), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n406_), .B(new_n346_), .C1(new_n317_), .C2(new_n403_), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n402_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n405_), .A2(new_n407_), .A3(new_n402_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G22gat), .B(G50gat), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n317_), .A2(new_n403_), .A3(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n414_), .B1(new_n317_), .B2(new_n403_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n413_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n417_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT96), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n421_), .B1(new_n408_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n411_), .A2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n409_), .A2(new_n421_), .A3(new_n422_), .A4(new_n410_), .ZN(new_n425_));
  AND2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT105), .B1(new_n400_), .B2(new_n426_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n388_), .A2(new_n389_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT105), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n424_), .A2(new_n425_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n428_), .A2(new_n429_), .A3(new_n430_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n334_), .B1(new_n427_), .B2(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n375_), .A2(KEYINPUT32), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n381_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(new_n434_), .B1(new_n433_), .B2(new_n392_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n331_), .A2(new_n332_), .A3(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n280_), .B1(new_n329_), .B2(new_n323_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n280_), .B1(new_n322_), .B2(new_n320_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n327_), .A2(new_n314_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n438_), .B1(new_n439_), .B2(new_n320_), .ZN(new_n440_));
  OAI21_X1  g239(.A(KEYINPUT33), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n388_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n325_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n441_), .A2(new_n442_), .A3(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n436_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n430_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n430_), .B1(new_n332_), .B2(new_n331_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n428_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n273_), .A2(new_n274_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n432_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G57gat), .B(G64gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT68), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n454_), .A2(KEYINPUT11), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G71gat), .B(G78gat), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  OR2_X1    g256(.A1(new_n453_), .A2(KEYINPUT68), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT11), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n453_), .A2(KEYINPUT68), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n455_), .A2(new_n457_), .A3(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n454_), .A2(KEYINPUT11), .A3(new_n456_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G15gat), .B(G22gat), .ZN(new_n466_));
  INV_X1    g265(.A(G1gat), .ZN(new_n467_));
  INV_X1    g266(.A(G8gat), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT14), .B1(new_n467_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n466_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G1gat), .B(G8gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G231gat), .A2(G233gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n465_), .B(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT79), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G127gat), .B(G155gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT16), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G183gat), .B(G211gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT17), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n476_), .B(new_n481_), .ZN(new_n482_));
  OR3_X1    g281(.A1(new_n475_), .A2(KEYINPUT17), .A3(new_n480_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT78), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT6), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(G99gat), .A3(G106gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  XOR2_X1   g290(.A(KEYINPUT10), .B(G99gat), .Z(new_n492_));
  INV_X1    g291(.A(G106gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT64), .B(G92gat), .Z(new_n495_));
  AOI21_X1  g294(.A(KEYINPUT9), .B1(new_n495_), .B2(G85gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(G85gat), .A2(G92gat), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n497_), .B1(new_n498_), .B2(KEYINPUT65), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n499_), .B1(KEYINPUT65), .B2(new_n497_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n491_), .B(new_n494_), .C1(new_n496_), .C2(new_n500_), .ZN(new_n501_));
  OR3_X1    g300(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n502_));
  OAI21_X1  g301(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT66), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT66), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n505_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n491_), .A2(new_n502_), .A3(new_n504_), .A4(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT8), .ZN(new_n508_));
  XOR2_X1   g307(.A(G85gat), .B(G92gat), .Z(new_n509_));
  AND3_X1   g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n508_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n501_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT71), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n507_), .A2(new_n509_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(KEYINPUT8), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT71), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n517_), .A2(new_n518_), .A3(new_n501_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n513_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G29gat), .B(G36gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(G43gat), .B(G50gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT15), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n520_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n512_), .A2(KEYINPUT67), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT67), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n501_), .B(new_n527_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n523_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G232gat), .A2(G233gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT34), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT35), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n532_), .B(KEYINPUT75), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n531_), .A2(KEYINPUT35), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n525_), .A2(new_n529_), .A3(KEYINPUT76), .A4(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n513_), .A2(new_n519_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n524_), .ZN(new_n538_));
  OAI211_X1 g337(.A(new_n529_), .B(new_n535_), .C1(new_n537_), .C2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT76), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n525_), .A2(new_n529_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n532_), .ZN(new_n543_));
  AOI22_X1  g342(.A1(new_n536_), .A2(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G190gat), .B(G218gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT74), .ZN(new_n546_));
  XOR2_X1   g345(.A(G134gat), .B(G162gat), .Z(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT36), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n544_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n536_), .A2(new_n541_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n548_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(KEYINPUT36), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n542_), .A2(new_n543_), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n552_), .A2(new_n554_), .A3(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT77), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(KEYINPUT77), .B1(new_n544_), .B2(new_n554_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n486_), .B(new_n551_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT37), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n556_), .A2(new_n557_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n544_), .A2(KEYINPUT77), .A3(new_n554_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n565_), .A2(new_n486_), .A3(KEYINPUT37), .A4(new_n551_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n562_), .A2(new_n566_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n452_), .A2(new_n485_), .A3(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(G230gat), .ZN(new_n569_));
  INV_X1    g368(.A(G233gat), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n526_), .A2(new_n528_), .A3(new_n464_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT69), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT69), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n526_), .A2(new_n574_), .A3(new_n464_), .A4(new_n528_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(KEYINPUT70), .A3(new_n575_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n527_), .B1(new_n517_), .B2(new_n501_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n528_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n465_), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n576_), .A2(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(KEYINPUT70), .B1(new_n573_), .B2(new_n575_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n571_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n465_), .A2(new_n513_), .A3(new_n519_), .A4(KEYINPUT12), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n464_), .B1(new_n526_), .B2(new_n528_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n583_), .B1(new_n584_), .B2(KEYINPUT12), .ZN(new_n585_));
  INV_X1    g384(.A(new_n571_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n572_), .A2(new_n586_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G120gat), .B(G148gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT5), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G176gat), .B(G204gat), .ZN(new_n592_));
  XOR2_X1   g391(.A(new_n591_), .B(new_n592_), .Z(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n582_), .A2(new_n589_), .A3(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT72), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT72), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n582_), .A2(new_n597_), .A3(new_n589_), .A4(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n596_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n582_), .A2(new_n589_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(new_n593_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n599_), .B(new_n601_), .C1(KEYINPUT73), .C2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n573_), .A2(new_n575_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT70), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n606_), .A2(new_n579_), .A3(new_n576_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n588_), .B1(new_n607_), .B2(new_n571_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n597_), .B1(new_n608_), .B2(new_n594_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n598_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n601_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT73), .B(KEYINPUT13), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n603_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT80), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n523_), .B(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n472_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT81), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n524_), .A2(new_n472_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(G229gat), .A2(G233gat), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n617_), .A2(new_n618_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT82), .Z(new_n626_));
  AND2_X1   g425(.A1(new_n626_), .A2(new_n620_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n624_), .B1(new_n627_), .B2(new_n623_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G113gat), .B(G141gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(G169gat), .B(G197gat), .ZN(new_n630_));
  XOR2_X1   g429(.A(new_n629_), .B(new_n630_), .Z(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n628_), .A2(new_n632_), .ZN(new_n633_));
  OAI211_X1 g432(.A(new_n624_), .B(new_n631_), .C1(new_n627_), .C2(new_n623_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n615_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n568_), .A2(new_n637_), .ZN(new_n638_));
  NOR3_X1   g437(.A1(new_n638_), .A2(G1gat), .A3(new_n333_), .ZN(new_n639_));
  XNOR2_X1  g438(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n331_), .A2(new_n332_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n642_), .A2(new_n451_), .ZN(new_n643_));
  NOR3_X1   g442(.A1(new_n400_), .A2(new_n426_), .A3(KEYINPUT105), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n429_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n643_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  AOI22_X1  g445(.A1(new_n446_), .A2(new_n430_), .B1(new_n448_), .B2(new_n428_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n646_), .B1(new_n647_), .B2(new_n275_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n565_), .A2(new_n551_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n614_), .A2(new_n484_), .A3(new_n635_), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n651_), .A2(KEYINPUT107), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT107), .ZN(new_n655_));
  INV_X1    g454(.A(new_n652_), .ZN(new_n656_));
  NOR3_X1   g455(.A1(new_n642_), .A2(new_n430_), .A3(new_n400_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n426_), .B1(new_n436_), .B2(new_n445_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n451_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n649_), .B1(new_n659_), .B2(new_n646_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n655_), .B1(new_n656_), .B2(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n333_), .B1(new_n654_), .B2(new_n662_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n641_), .B1(new_n663_), .B2(new_n467_), .ZN(G1324gat));
  NAND3_X1  g463(.A1(new_n656_), .A2(new_n400_), .A3(new_n660_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(G8gat), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n666_), .B(KEYINPUT39), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n568_), .A2(new_n468_), .A3(new_n400_), .A4(new_n637_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(G1325gat));
  OR3_X1    g470(.A1(new_n638_), .A2(G15gat), .A3(new_n451_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n275_), .B1(new_n653_), .B2(new_n661_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n673_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n674_));
  AOI21_X1  g473(.A(KEYINPUT41), .B1(new_n673_), .B2(G15gat), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n672_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT109), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n678_));
  OAI211_X1 g477(.A(new_n678_), .B(new_n672_), .C1(new_n674_), .C2(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1326gat));
  AOI21_X1  g479(.A(new_n430_), .B1(new_n654_), .B2(new_n662_), .ZN(new_n681_));
  INV_X1    g480(.A(G22gat), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT42), .ZN(new_n684_));
  NOR2_X1   g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  NOR3_X1   g484(.A1(new_n681_), .A2(KEYINPUT42), .A3(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n426_), .A2(new_n682_), .ZN(new_n687_));
  OAI22_X1  g486(.A1(new_n685_), .A2(new_n686_), .B1(new_n638_), .B2(new_n687_), .ZN(G1327gat));
  NAND2_X1  g487(.A1(new_n649_), .A2(new_n485_), .ZN(new_n689_));
  XOR2_X1   g488(.A(new_n689_), .B(KEYINPUT113), .Z(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n452_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(new_n637_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G29gat), .B1(new_n693_), .B2(new_n642_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n614_), .A2(new_n485_), .A3(new_n635_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n562_), .A2(new_n698_), .A3(new_n566_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n698_), .B1(new_n562_), .B2(new_n566_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n697_), .B1(new_n701_), .B2(new_n648_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n567_), .A2(new_n697_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n703_), .B1(new_n659_), .B2(new_n646_), .ZN(new_n704_));
  OAI211_X1 g503(.A(KEYINPUT44), .B(new_n696_), .C1(new_n702_), .C2(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(KEYINPUT112), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n567_), .A2(KEYINPUT110), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n562_), .A2(new_n698_), .A3(new_n566_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(KEYINPUT43), .B1(new_n452_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n704_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT112), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n712_), .A2(new_n713_), .A3(KEYINPUT44), .A4(new_n696_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n706_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n712_), .A2(new_n696_), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n716_), .A2(new_n718_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n715_), .A2(new_n719_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n642_), .A2(G29gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n694_), .B1(new_n720_), .B2(new_n721_), .ZN(G1328gat));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723_));
  INV_X1    g522(.A(G36gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n428_), .B1(new_n716_), .B2(new_n718_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n715_), .B2(new_n725_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n691_), .A2(new_n724_), .A3(new_n400_), .A4(new_n637_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT45), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n723_), .B1(new_n726_), .B2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n695_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n400_), .B1(new_n731_), .B2(new_n717_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n706_), .B2(new_n714_), .ZN(new_n733_));
  OAI211_X1 g532(.A(KEYINPUT46), .B(new_n728_), .C1(new_n733_), .C2(new_n724_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(G1329gat));
  INV_X1    g534(.A(G43gat), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n451_), .A2(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n713_), .B1(new_n731_), .B2(KEYINPUT44), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n705_), .A2(KEYINPUT112), .ZN(new_n739_));
  OAI211_X1 g538(.A(new_n719_), .B(new_n737_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n692_), .B2(new_n451_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT47), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n740_), .A2(new_n744_), .A3(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1330gat));
  AOI21_X1  g545(.A(G50gat), .B1(new_n693_), .B2(new_n426_), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n426_), .A2(G50gat), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n747_), .B1(new_n720_), .B2(new_n748_), .ZN(G1331gat));
  NOR2_X1   g548(.A1(new_n614_), .A2(new_n635_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n568_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(G57gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n752_), .A3(new_n642_), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n660_), .A2(new_n484_), .A3(new_n750_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G57gat), .B1(new_n755_), .B2(new_n333_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n756_), .ZN(G1332gat));
  INV_X1    g556(.A(G64gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(new_n754_), .B2(new_n400_), .ZN(new_n759_));
  XOR2_X1   g558(.A(new_n759_), .B(KEYINPUT48), .Z(new_n760_));
  NAND3_X1  g559(.A1(new_n751_), .A2(new_n758_), .A3(new_n400_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(G1333gat));
  INV_X1    g561(.A(G71gat), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n763_), .B1(new_n754_), .B2(new_n275_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT49), .Z(new_n765_));
  NAND3_X1  g564(.A1(new_n751_), .A2(new_n763_), .A3(new_n275_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1334gat));
  INV_X1    g566(.A(G78gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n754_), .B2(new_n426_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT50), .Z(new_n770_));
  NAND2_X1  g569(.A1(new_n426_), .A2(new_n768_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT114), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n751_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n770_), .A2(new_n773_), .ZN(G1335gat));
  AND2_X1   g573(.A1(new_n691_), .A2(new_n750_), .ZN(new_n775_));
  INV_X1    g574(.A(G85gat), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(new_n642_), .ZN(new_n777_));
  AND3_X1   g576(.A1(new_n712_), .A2(new_n485_), .A3(new_n750_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n642_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n777_), .B1(new_n780_), .B2(new_n776_), .ZN(G1336gat));
  AOI21_X1  g580(.A(G92gat), .B1(new_n775_), .B2(new_n400_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n400_), .A2(new_n495_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n778_), .B2(new_n783_), .ZN(G1337gat));
  INV_X1    g583(.A(G99gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n778_), .B2(new_n275_), .ZN(new_n786_));
  AND2_X1   g585(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n775_), .A2(new_n275_), .A3(new_n492_), .ZN(new_n788_));
  OR3_X1    g587(.A1(new_n786_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n787_), .B1(new_n786_), .B2(new_n788_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1338gat));
  NAND4_X1  g590(.A1(new_n691_), .A2(new_n493_), .A3(new_n426_), .A4(new_n750_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n792_), .B(new_n793_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n712_), .A2(new_n426_), .A3(new_n485_), .A4(new_n750_), .ZN(new_n795_));
  XOR2_X1   g594(.A(KEYINPUT117), .B(KEYINPUT52), .Z(new_n796_));
  AND3_X1   g595(.A1(new_n795_), .A2(G106gat), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(new_n795_), .B2(G106gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT53), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n794_), .B(new_n801_), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1339gat));
  NOR2_X1   g602(.A1(new_n644_), .A2(new_n645_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n642_), .A2(new_n275_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT121), .ZN(new_n808_));
  INV_X1    g607(.A(new_n623_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n622_), .A2(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n810_), .B(new_n632_), .C1(new_n627_), .C2(new_n809_), .ZN(new_n811_));
  AND2_X1   g610(.A1(new_n634_), .A2(new_n811_), .ZN(new_n812_));
  AND2_X1   g611(.A1(new_n572_), .A2(new_n586_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT12), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n579_), .A2(new_n814_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n813_), .A2(new_n815_), .A3(KEYINPUT55), .A4(new_n583_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT120), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n464_), .A2(new_n814_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n814_), .A2(new_n579_), .B1(new_n520_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT120), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n819_), .A2(new_n820_), .A3(KEYINPUT55), .A4(new_n813_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT55), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n585_), .B2(new_n587_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n571_), .B1(new_n585_), .B2(new_n604_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n817_), .A2(new_n821_), .A3(new_n823_), .A4(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n593_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(KEYINPUT56), .ZN(new_n827_));
  INV_X1    g626(.A(KEYINPUT56), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n825_), .A2(new_n828_), .A3(new_n593_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n599_), .A2(new_n812_), .A3(new_n827_), .A4(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n825_), .A2(new_n828_), .A3(new_n593_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n828_), .B1(new_n825_), .B2(new_n593_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n835_), .A2(KEYINPUT58), .A3(new_n599_), .A4(new_n812_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n832_), .A2(new_n567_), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n611_), .A2(new_n812_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n599_), .A2(new_n635_), .A3(new_n827_), .A4(new_n829_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n649_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n837_), .B1(KEYINPUT57), .B2(new_n840_), .ZN(new_n841_));
  AND2_X1   g640(.A1(new_n840_), .A2(KEYINPUT57), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n808_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  OR2_X1    g642(.A1(new_n840_), .A2(KEYINPUT57), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n840_), .A2(KEYINPUT57), .ZN(new_n845_));
  NAND4_X1  g644(.A1(new_n844_), .A2(KEYINPUT121), .A3(new_n845_), .A4(new_n837_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n843_), .A2(new_n846_), .A3(new_n485_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT118), .B(KEYINPUT54), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n484_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n850_), .A2(new_n635_), .ZN(new_n851_));
  AND3_X1   g650(.A1(new_n562_), .A2(new_n851_), .A3(new_n566_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n848_), .ZN(new_n853_));
  AND3_X1   g652(.A1(new_n614_), .A2(new_n852_), .A3(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n614_), .B2(new_n852_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n807_), .B1(new_n847_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n485_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(new_n856_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n806_), .A2(new_n858_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n859_), .B1(new_n861_), .B2(new_n863_), .ZN(new_n864_));
  AOI211_X1 g663(.A(KEYINPUT122), .B(new_n862_), .C1(new_n860_), .C2(new_n856_), .ZN(new_n865_));
  OAI22_X1  g664(.A1(new_n857_), .A2(new_n858_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  OAI21_X1  g665(.A(G113gat), .B1(new_n866_), .B2(new_n636_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n857_), .ZN(new_n868_));
  OR3_X1    g667(.A1(new_n868_), .A2(G113gat), .A3(new_n636_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n867_), .A2(new_n869_), .ZN(G1340gat));
  OAI21_X1  g669(.A(G120gat), .B1(new_n866_), .B2(new_n614_), .ZN(new_n871_));
  INV_X1    g670(.A(G120gat), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n872_), .B1(new_n614_), .B2(KEYINPUT60), .ZN(new_n873_));
  OAI211_X1 g672(.A(new_n857_), .B(new_n873_), .C1(KEYINPUT60), .C2(new_n872_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n871_), .A2(new_n874_), .ZN(G1341gat));
  OAI21_X1  g674(.A(G127gat), .B1(new_n866_), .B2(new_n485_), .ZN(new_n876_));
  OR3_X1    g675(.A1(new_n868_), .A2(G127gat), .A3(new_n485_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1342gat));
  INV_X1    g677(.A(new_n567_), .ZN(new_n879_));
  OAI21_X1  g678(.A(G134gat), .B1(new_n866_), .B2(new_n879_), .ZN(new_n880_));
  OR3_X1    g679(.A1(new_n868_), .A2(G134gat), .A3(new_n650_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n880_), .A2(new_n881_), .ZN(G1343gat));
  NAND2_X1  g681(.A1(new_n847_), .A2(new_n856_), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n400_), .A2(new_n275_), .A3(new_n333_), .A4(new_n430_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n886_), .A2(new_n286_), .A3(new_n635_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G141gat), .B1(new_n885_), .B2(new_n636_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1344gat));
  NAND3_X1  g688(.A1(new_n886_), .A2(new_n287_), .A3(new_n615_), .ZN(new_n890_));
  OAI21_X1  g689(.A(G148gat), .B1(new_n885_), .B2(new_n614_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(G1345gat));
  XNOR2_X1  g691(.A(KEYINPUT61), .B(G155gat), .ZN(new_n893_));
  OR3_X1    g692(.A1(new_n885_), .A2(new_n485_), .A3(new_n893_), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n893_), .B1(new_n885_), .B2(new_n485_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(G1346gat));
  INV_X1    g695(.A(G162gat), .ZN(new_n897_));
  NOR3_X1   g696(.A1(new_n885_), .A2(new_n897_), .A3(new_n709_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n886_), .A2(new_n649_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n897_), .B2(new_n899_), .ZN(G1347gat));
  NAND2_X1  g699(.A1(new_n643_), .A2(new_n400_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(KEYINPUT123), .ZN(new_n902_));
  OR3_X1    g701(.A1(new_n902_), .A2(KEYINPUT124), .A3(new_n636_), .ZN(new_n903_));
  OAI21_X1  g702(.A(KEYINPUT124), .B1(new_n902_), .B2(new_n636_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n903_), .A2(new_n430_), .A3(new_n904_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n860_), .A2(new_n856_), .ZN(new_n906_));
  OAI21_X1  g705(.A(G169gat), .B1(new_n905_), .B2(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT62), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n902_), .A2(new_n426_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n906_), .A2(new_n910_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n911_), .A2(new_n347_), .A3(new_n635_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n908_), .A2(new_n912_), .ZN(G1348gat));
  AOI21_X1  g712(.A(new_n910_), .B1(new_n847_), .B2(new_n856_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n614_), .A2(new_n348_), .ZN(new_n916_));
  AND3_X1   g715(.A1(new_n914_), .A2(new_n915_), .A3(new_n916_), .ZN(new_n917_));
  AOI21_X1  g716(.A(G176gat), .B1(new_n911_), .B2(new_n615_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n915_), .B1(new_n914_), .B2(new_n916_), .ZN(new_n919_));
  NOR3_X1   g718(.A1(new_n917_), .A2(new_n918_), .A3(new_n919_), .ZN(G1349gat));
  AOI21_X1  g719(.A(G183gat), .B1(new_n914_), .B2(new_n484_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n485_), .A2(new_n221_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n921_), .B1(new_n911_), .B2(new_n922_), .ZN(G1350gat));
  NAND3_X1  g722(.A1(new_n911_), .A2(new_n352_), .A3(new_n649_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n911_), .ZN(new_n925_));
  OAI21_X1  g724(.A(G190gat), .B1(new_n925_), .B2(new_n879_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n924_), .A2(new_n926_), .ZN(G1351gat));
  NAND2_X1  g726(.A1(new_n448_), .A2(new_n451_), .ZN(new_n928_));
  OR2_X1    g727(.A1(new_n928_), .A2(KEYINPUT126), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(KEYINPUT126), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n929_), .A2(new_n400_), .A3(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n931_), .B1(new_n847_), .B2(new_n856_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n932_), .A2(new_n635_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g733(.A1(new_n932_), .A2(new_n615_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G204gat), .ZN(G1353gat));
  AOI211_X1 g735(.A(KEYINPUT63), .B(G211gat), .C1(new_n932_), .C2(new_n484_), .ZN(new_n937_));
  AND2_X1   g736(.A1(new_n932_), .A2(new_n484_), .ZN(new_n938_));
  XOR2_X1   g737(.A(KEYINPUT63), .B(G211gat), .Z(new_n939_));
  AOI21_X1  g738(.A(new_n937_), .B1(new_n938_), .B2(new_n939_), .ZN(G1354gat));
  INV_X1    g739(.A(KEYINPUT127), .ZN(new_n941_));
  INV_X1    g740(.A(G218gat), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n942_), .B1(new_n932_), .B2(new_n567_), .ZN(new_n943_));
  INV_X1    g742(.A(new_n931_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n650_), .A2(G218gat), .ZN(new_n945_));
  AND3_X1   g744(.A1(new_n883_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  OAI21_X1  g745(.A(new_n941_), .B1(new_n943_), .B2(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n932_), .A2(new_n945_), .ZN(new_n948_));
  AOI211_X1 g747(.A(new_n879_), .B(new_n931_), .C1(new_n847_), .C2(new_n856_), .ZN(new_n949_));
  OAI211_X1 g748(.A(new_n948_), .B(KEYINPUT127), .C1(new_n949_), .C2(new_n942_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n947_), .A2(new_n950_), .ZN(G1355gat));
endmodule


