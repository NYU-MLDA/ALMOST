//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0 1 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 0 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n941_, new_n942_,
    new_n943_, new_n945_, new_n946_, new_n947_, new_n949_, new_n950_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n957_, new_n958_,
    new_n959_;
  INV_X1    g000(.A(KEYINPUT79), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  AOI21_X1  g002(.A(new_n202_), .B1(new_n203_), .B2(KEYINPUT23), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(KEYINPUT23), .ZN(new_n205_));
  AOI21_X1  g004(.A(new_n204_), .B1(new_n205_), .B2(new_n202_), .ZN(new_n206_));
  INV_X1    g005(.A(G183gat), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT77), .B(G190gat), .Z(new_n208_));
  AOI21_X1  g007(.A(new_n206_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  OR2_X1    g008(.A1(new_n209_), .A2(KEYINPUT80), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(KEYINPUT80), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT22), .B(G169gat), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n214_), .A2(KEYINPUT78), .ZN(new_n215_));
  INV_X1    g014(.A(G169gat), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n216_), .A2(KEYINPUT22), .ZN(new_n217_));
  AOI21_X1  g016(.A(G176gat), .B1(new_n217_), .B2(KEYINPUT78), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n213_), .B1(new_n215_), .B2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n210_), .A2(new_n211_), .A3(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n212_), .A2(KEYINPUT24), .ZN(new_n221_));
  INV_X1    g020(.A(G176gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n216_), .A2(new_n222_), .ZN(new_n223_));
  MUX2_X1   g022(.A(KEYINPUT24), .B(new_n221_), .S(new_n223_), .Z(new_n224_));
  MUX2_X1   g023(.A(G190gat), .B(new_n208_), .S(KEYINPUT26), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n207_), .A2(KEYINPUT25), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT76), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n207_), .A2(KEYINPUT76), .A3(KEYINPUT25), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n207_), .A2(KEYINPUT25), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n224_), .B(new_n205_), .C1(new_n225_), .C2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n220_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G71gat), .B(G99gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n234_), .B(G43gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n233_), .B(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT81), .B(KEYINPUT31), .Z(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  XOR2_X1   g037(.A(G127gat), .B(G134gat), .Z(new_n239_));
  XOR2_X1   g038(.A(G113gat), .B(G120gat), .Z(new_n240_));
  XOR2_X1   g039(.A(new_n239_), .B(new_n240_), .Z(new_n241_));
  NAND2_X1  g040(.A1(G227gat), .A2(G233gat), .ZN(new_n242_));
  INV_X1    g041(.A(G15gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT30), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n241_), .B(new_n245_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n238_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n238_), .A2(new_n246_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G8gat), .B(G36gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT18), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G64gat), .B(G92gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n252_), .B(new_n253_), .Z(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT32), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G197gat), .B(G204gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT85), .ZN(new_n257_));
  INV_X1    g056(.A(G204gat), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(G197gat), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n257_), .B(KEYINPUT21), .C1(KEYINPUT85), .C2(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT86), .ZN(new_n261_));
  XOR2_X1   g060(.A(G211gat), .B(G218gat), .Z(new_n262_));
  INV_X1    g061(.A(KEYINPUT21), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n262_), .B1(new_n263_), .B2(new_n256_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n256_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n266_), .A2(KEYINPUT21), .A3(new_n262_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n265_), .A2(new_n267_), .ZN(new_n268_));
  OR2_X1    g067(.A1(G183gat), .A2(G190gat), .ZN(new_n269_));
  AND2_X1   g068(.A1(new_n205_), .A2(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n213_), .B1(new_n214_), .B2(new_n222_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT26), .B(G190gat), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n274_), .A2(new_n226_), .A3(new_n230_), .ZN(new_n275_));
  AND2_X1   g074(.A1(new_n224_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n206_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n273_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n268_), .A2(new_n279_), .ZN(new_n280_));
  OAI211_X1 g079(.A(new_n280_), .B(KEYINPUT20), .C1(new_n233_), .C2(new_n268_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G226gat), .A2(G233gat), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n282_), .B(KEYINPUT19), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n283_), .B(KEYINPUT89), .Z(new_n284_));
  NOR2_X1   g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT20), .ZN(new_n286_));
  AND2_X1   g085(.A1(new_n265_), .A2(new_n267_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n286_), .B1(new_n287_), .B2(new_n278_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n233_), .A2(new_n268_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(new_n283_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT92), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n285_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n283_), .ZN(new_n294_));
  AOI211_X1 g093(.A(new_n292_), .B(new_n294_), .C1(new_n288_), .C2(new_n289_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n255_), .B1(new_n293_), .B2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G225gat), .A2(G233gat), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G141gat), .A2(G148gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G141gat), .A2(G148gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NOR2_X1   g100(.A1(G155gat), .A2(G162gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n302_), .B1(KEYINPUT1), .B2(new_n303_), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n303_), .A2(KEYINPUT1), .ZN(new_n305_));
  AOI211_X1 g104(.A(new_n299_), .B(new_n301_), .C1(new_n304_), .C2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G155gat), .B(G162gat), .Z(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT83), .ZN(new_n308_));
  AOI21_X1  g107(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT82), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT3), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n299_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n301_), .A2(KEYINPUT2), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .A4(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n306_), .B1(new_n308_), .B2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n241_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n318_), .A2(KEYINPUT90), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n317_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(KEYINPUT4), .A3(new_n320_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(KEYINPUT4), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n322_), .A2(KEYINPUT90), .A3(new_n318_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n298_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G1gat), .B(G29gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(G85gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(KEYINPUT0), .B(G57gat), .ZN(new_n327_));
  XOR2_X1   g126(.A(new_n326_), .B(new_n327_), .Z(new_n328_));
  XNOR2_X1  g127(.A(new_n316_), .B(new_n241_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n298_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  OR3_X1    g130(.A1(new_n324_), .A2(new_n328_), .A3(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n328_), .B1(new_n324_), .B2(new_n331_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n284_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n287_), .A2(new_n220_), .A3(new_n232_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n286_), .B1(new_n268_), .B2(new_n279_), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n335_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n288_), .A2(new_n289_), .A3(new_n294_), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n340_), .A3(new_n255_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n334_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT33), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n333_), .A2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(KEYINPUT33), .B(new_n328_), .C1(new_n324_), .C2(new_n331_), .ZN(new_n345_));
  OR2_X1    g144(.A1(new_n329_), .A2(KEYINPUT91), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n329_), .A2(KEYINPUT91), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n346_), .A2(new_n347_), .A3(new_n330_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n328_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n321_), .A2(new_n298_), .A3(new_n323_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n348_), .A2(new_n349_), .A3(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n344_), .A2(new_n345_), .A3(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n254_), .ZN(new_n353_));
  AND3_X1   g152(.A1(new_n288_), .A2(new_n289_), .A3(new_n294_), .ZN(new_n354_));
  OAI21_X1  g153(.A(new_n353_), .B1(new_n354_), .B2(new_n338_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n339_), .A2(new_n340_), .A3(new_n254_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OAI22_X1  g156(.A1(new_n297_), .A2(new_n342_), .B1(new_n352_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(G228gat), .A2(G233gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n359_), .B(KEYINPUT84), .Z(new_n360_));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n316_), .A2(new_n361_), .ZN(new_n362_));
  OAI211_X1 g161(.A(KEYINPUT87), .B(new_n360_), .C1(new_n287_), .C2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n362_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n360_), .A2(KEYINPUT87), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n360_), .A2(KEYINPUT87), .ZN(new_n366_));
  NAND4_X1  g165(.A1(new_n268_), .A2(new_n364_), .A3(new_n365_), .A4(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n363_), .A2(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G78gat), .B(G106gat), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n363_), .A2(new_n369_), .A3(new_n367_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n316_), .A2(new_n361_), .ZN(new_n373_));
  XOR2_X1   g172(.A(G22gat), .B(G50gat), .Z(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT28), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n373_), .B(new_n375_), .ZN(new_n376_));
  AND4_X1   g175(.A1(KEYINPUT88), .A2(new_n371_), .A3(new_n372_), .A4(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT88), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n372_), .A2(new_n378_), .ZN(new_n379_));
  AOI22_X1  g178(.A1(new_n379_), .A2(new_n376_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n377_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n358_), .A2(new_n382_), .A3(KEYINPUT93), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT27), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n354_), .A2(new_n338_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n384_), .B1(new_n385_), .B2(new_n254_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n294_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n387_));
  OAI22_X1  g186(.A1(new_n387_), .A2(KEYINPUT92), .B1(new_n284_), .B2(new_n281_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n353_), .B1(new_n388_), .B2(new_n295_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n386_), .A2(new_n389_), .B1(new_n357_), .B2(new_n384_), .ZN(new_n390_));
  NOR3_X1   g189(.A1(new_n377_), .A2(new_n380_), .A3(new_n334_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n383_), .A2(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT93), .B1(new_n358_), .B2(new_n382_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n250_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n334_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n249_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n382_), .A2(new_n390_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n395_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT94), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G15gat), .B(G22gat), .ZN(new_n403_));
  INV_X1    g202(.A(G1gat), .ZN(new_n404_));
  INV_X1    g203(.A(G8gat), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT14), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G1gat), .B(G8gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G29gat), .B(G36gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G43gat), .B(G50gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(new_n410_), .B(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n409_), .B(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT74), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G229gat), .A2(G233gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  XOR2_X1   g216(.A(new_n410_), .B(new_n411_), .Z(new_n418_));
  OR2_X1    g217(.A1(new_n409_), .A2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n412_), .B(KEYINPUT15), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n409_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n415_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n417_), .A2(KEYINPUT75), .A3(new_n423_), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n423_), .A2(KEYINPUT75), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G113gat), .B(G141gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(G169gat), .B(G197gat), .ZN(new_n428_));
  XOR2_X1   g227(.A(new_n427_), .B(new_n428_), .Z(new_n429_));
  OR2_X1    g228(.A1(new_n426_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n429_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n401_), .A2(new_n402_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT93), .ZN(new_n434_));
  INV_X1    g233(.A(new_n357_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n352_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n385_), .A2(new_n255_), .B1(new_n332_), .B2(new_n333_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n255_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n438_), .B1(new_n388_), .B2(new_n295_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n435_), .A2(new_n436_), .B1(new_n437_), .B2(new_n439_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n434_), .B1(new_n440_), .B2(new_n381_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n441_), .A2(new_n392_), .A3(new_n383_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n399_), .B1(new_n442_), .B2(new_n250_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n432_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT94), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n433_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447_));
  OR2_X1    g246(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n448_));
  INV_X1    g247(.A(G106gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT64), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT64), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n451_), .A2(G106gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n448_), .A2(new_n450_), .A3(new_n452_), .A4(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G99gat), .A2(G106gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT6), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n457_), .A2(G99gat), .A3(G106gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n456_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  OR2_X1    g259(.A1(new_n460_), .A2(KEYINPUT9), .ZN(new_n461_));
  INV_X1    g260(.A(G85gat), .ZN(new_n462_));
  INV_X1    g261(.A(G92gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n464_), .A2(KEYINPUT9), .A3(new_n460_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n454_), .A2(new_n459_), .A3(new_n461_), .A4(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(new_n460_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n456_), .A2(new_n458_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT7), .ZN(new_n471_));
  INV_X1    g270(.A(G99gat), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(new_n472_), .A3(new_n449_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n469_), .B1(new_n470_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(KEYINPUT8), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n457_), .B1(G99gat), .B2(G106gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n455_), .A2(KEYINPUT6), .ZN(new_n479_));
  OAI211_X1 g278(.A(new_n474_), .B(new_n473_), .C1(new_n478_), .C2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT8), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n469_), .ZN(new_n482_));
  AOI21_X1  g281(.A(new_n467_), .B1(new_n477_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n412_), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT69), .ZN(new_n485_));
  INV_X1    g284(.A(new_n474_), .ZN(new_n486_));
  NOR3_X1   g285(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  AOI211_X1 g287(.A(KEYINPUT8), .B(new_n468_), .C1(new_n488_), .C2(new_n459_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n481_), .B1(new_n480_), .B2(new_n469_), .ZN(new_n490_));
  NOR3_X1   g289(.A1(new_n489_), .A2(new_n490_), .A3(KEYINPUT66), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT66), .ZN(new_n492_));
  AOI21_X1  g291(.A(new_n492_), .B1(new_n477_), .B2(new_n482_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n466_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  AND2_X1   g293(.A1(new_n494_), .A2(new_n421_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G232gat), .A2(G233gat), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT34), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n497_), .A2(KEYINPUT35), .ZN(new_n498_));
  NOR3_X1   g297(.A1(new_n485_), .A2(new_n495_), .A3(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(KEYINPUT35), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  OAI211_X1 g300(.A(KEYINPUT35), .B(new_n497_), .C1(new_n485_), .C2(new_n495_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(KEYINPUT72), .ZN(new_n503_));
  XOR2_X1   g302(.A(G190gat), .B(G218gat), .Z(new_n504_));
  XNOR2_X1  g303(.A(G134gat), .B(G162gat), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n504_), .B(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n503_), .B1(KEYINPUT36), .B2(new_n508_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n508_), .A2(KEYINPUT36), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n501_), .A2(new_n502_), .A3(KEYINPUT72), .A4(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n509_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n508_), .A2(KEYINPUT36), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n513_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n447_), .B1(new_n512_), .B2(new_n515_), .ZN(new_n516_));
  AOI211_X1 g315(.A(KEYINPUT37), .B(new_n514_), .C1(new_n509_), .C2(new_n511_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT12), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G57gat), .B(G64gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G71gat), .B(G78gat), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n520_), .A2(new_n521_), .A3(KEYINPUT11), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(KEYINPUT11), .ZN(new_n523_));
  INV_X1    g322(.A(new_n521_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n520_), .A2(KEYINPUT11), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n522_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n519_), .B1(new_n483_), .B2(new_n527_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n527_), .B(new_n466_), .C1(new_n489_), .C2(new_n490_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n527_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT12), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n494_), .A2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT67), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n530_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(G230gat), .A2(G233gat), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n494_), .A2(KEYINPUT67), .A3(new_n533_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n536_), .A2(KEYINPUT68), .A3(new_n537_), .A4(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT66), .B1(new_n489_), .B2(new_n490_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n477_), .A2(new_n492_), .A3(new_n482_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n467_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n535_), .B1(new_n542_), .B2(new_n532_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n466_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT12), .B1(new_n544_), .B2(new_n531_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n529_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NAND4_X1  g346(.A1(new_n538_), .A2(new_n543_), .A3(new_n537_), .A4(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT68), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n546_), .A2(KEYINPUT65), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n483_), .A2(new_n527_), .ZN(new_n552_));
  OR2_X1    g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n537_), .B1(new_n552_), .B2(KEYINPUT65), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n539_), .A2(new_n550_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G120gat), .B(G148gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT5), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G176gat), .B(G204gat), .ZN(new_n558_));
  XOR2_X1   g357(.A(new_n557_), .B(new_n558_), .Z(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n555_), .A2(new_n560_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n561_), .A2(KEYINPUT13), .A3(new_n562_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n409_), .B(new_n527_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G231gat), .A2(G233gat), .ZN(new_n569_));
  XOR2_X1   g368(.A(new_n568_), .B(new_n569_), .Z(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT17), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G127gat), .B(G155gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G183gat), .B(G211gat), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  OR3_X1    g376(.A1(new_n571_), .A2(new_n572_), .A3(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(KEYINPUT17), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n571_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n578_), .A2(new_n580_), .ZN(new_n581_));
  NOR3_X1   g380(.A1(new_n518_), .A2(new_n567_), .A3(new_n581_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n396_), .A2(G1gat), .ZN(new_n583_));
  AND4_X1   g382(.A1(KEYINPUT95), .A2(new_n446_), .A3(new_n582_), .A4(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n582_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n585_), .B1(new_n433_), .B2(new_n445_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT95), .B1(new_n586_), .B2(new_n583_), .ZN(new_n587_));
  OAI21_X1  g386(.A(KEYINPUT96), .B1(new_n584_), .B2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n446_), .A2(new_n582_), .A3(new_n583_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT95), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n586_), .A2(KEYINPUT95), .A3(new_n583_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT96), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n591_), .A2(new_n592_), .A3(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n588_), .A2(KEYINPUT38), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n567_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n581_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(new_n432_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n512_), .A2(new_n515_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n401_), .A2(KEYINPUT97), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT97), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n602_), .B1(new_n443_), .B2(new_n599_), .ZN(new_n603_));
  AOI21_X1  g402(.A(new_n598_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n604_), .A2(new_n334_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(G1gat), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n595_), .A2(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT38), .B1(new_n588_), .B2(new_n594_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT98), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n588_), .A2(new_n594_), .ZN(new_n610_));
  INV_X1    g409(.A(KEYINPUT38), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT98), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n612_), .A2(new_n613_), .A3(new_n606_), .A4(new_n595_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n609_), .A2(new_n614_), .ZN(G1324gat));
  INV_X1    g414(.A(new_n390_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n586_), .A2(new_n405_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n604_), .A2(KEYINPUT99), .A3(new_n616_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n619_), .A2(G8gat), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n604_), .A2(new_n616_), .ZN(new_n621_));
  INV_X1    g420(.A(KEYINPUT99), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n618_), .B1(new_n620_), .B2(new_n623_), .ZN(new_n624_));
  AND4_X1   g423(.A1(new_n618_), .A2(new_n623_), .A3(G8gat), .A4(new_n619_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n617_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT40), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  OAI211_X1 g427(.A(KEYINPUT40), .B(new_n617_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(G1325gat));
  NAND3_X1  g429(.A1(new_n586_), .A2(new_n243_), .A3(new_n249_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n604_), .A2(new_n249_), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n632_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT41), .B1(new_n632_), .B2(G15gat), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n631_), .B1(new_n633_), .B2(new_n634_), .ZN(G1326gat));
  INV_X1    g434(.A(G22gat), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n586_), .A2(new_n636_), .A3(new_n381_), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT42), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n604_), .A2(new_n381_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n638_), .B1(new_n639_), .B2(G22gat), .ZN(new_n640_));
  AOI211_X1 g439(.A(KEYINPUT42), .B(new_n636_), .C1(new_n604_), .C2(new_n381_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n637_), .B1(new_n640_), .B2(new_n641_), .ZN(G1327gat));
  NOR2_X1   g441(.A1(new_n600_), .A2(new_n597_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(new_n596_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n644_), .B1(new_n433_), .B2(new_n445_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  OR3_X1    g445(.A1(new_n646_), .A2(G29gat), .A3(new_n396_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n567_), .A2(new_n444_), .A3(new_n597_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n649_), .B1(new_n401_), .B2(new_n518_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n516_), .A2(new_n517_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n443_), .A2(KEYINPUT43), .A3(new_n651_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n648_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n401_), .A2(new_n649_), .A3(new_n518_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT43), .B1(new_n443_), .B2(new_n651_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(KEYINPUT44), .A3(new_n648_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n655_), .A2(new_n334_), .A3(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(KEYINPUT100), .A3(G29gat), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT100), .B1(new_n660_), .B2(G29gat), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n647_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT101), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n665_), .B(new_n647_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(G1328gat));
  INV_X1    g466(.A(KEYINPUT45), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n390_), .A2(G36gat), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n645_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n669_), .B1(new_n645_), .B2(new_n670_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n668_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n673_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n675_), .A2(KEYINPUT45), .A3(new_n671_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n674_), .A2(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT44), .B1(new_n658_), .B2(new_n648_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n648_), .ZN(new_n681_));
  AOI211_X1 g480(.A(new_n654_), .B(new_n681_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  AOI21_X1  g482(.A(KEYINPUT102), .B1(new_n683_), .B2(new_n616_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n655_), .A2(new_n616_), .A3(new_n659_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n686_));
  OAI21_X1  g485(.A(G36gat), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  OAI211_X1 g486(.A(new_n677_), .B(new_n679_), .C1(new_n684_), .C2(new_n687_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n684_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n674_), .A2(new_n676_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n678_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n688_), .A2(new_n691_), .ZN(G1329gat));
  NOR3_X1   g491(.A1(new_n646_), .A2(G43gat), .A3(new_n250_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n683_), .A2(new_n249_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n693_), .B1(new_n694_), .B2(G43gat), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g495(.A1(new_n646_), .A2(G50gat), .A3(new_n382_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n655_), .A2(new_n381_), .A3(new_n659_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT105), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n698_), .A2(new_n699_), .A3(G50gat), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n699_), .B1(new_n698_), .B2(G50gat), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(KEYINPUT106), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n704_));
  OAI211_X1 g503(.A(new_n704_), .B(new_n697_), .C1(new_n700_), .C2(new_n701_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n703_), .A2(new_n705_), .ZN(G1331gat));
  NOR2_X1   g505(.A1(new_n443_), .A2(new_n432_), .ZN(new_n707_));
  AND4_X1   g506(.A1(new_n567_), .A2(new_n707_), .A3(new_n597_), .A4(new_n651_), .ZN(new_n708_));
  AOI21_X1  g507(.A(G57gat), .B1(new_n708_), .B2(new_n334_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n567_), .A2(new_n444_), .A3(new_n597_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n710_), .B1(new_n601_), .B2(new_n603_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n396_), .A2(KEYINPUT107), .ZN(new_n712_));
  MUX2_X1   g511(.A(KEYINPUT107), .B(new_n712_), .S(G57gat), .Z(new_n713_));
  AOI21_X1  g512(.A(new_n709_), .B1(new_n711_), .B2(new_n713_), .ZN(G1332gat));
  INV_X1    g513(.A(G64gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n708_), .A2(new_n715_), .A3(new_n616_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n715_), .B1(new_n711_), .B2(new_n616_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n717_), .A2(new_n718_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n719_), .B2(new_n720_), .ZN(G1333gat));
  INV_X1    g520(.A(G71gat), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n249_), .A2(new_n722_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT108), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n708_), .A2(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n722_), .B1(new_n711_), .B2(new_n249_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT49), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n726_), .A2(new_n727_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1334gat));
  INV_X1    g529(.A(G78gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n708_), .A2(new_n731_), .A3(new_n381_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n711_), .B2(new_n381_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT50), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n733_), .A2(new_n734_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(G1335gat));
  NAND3_X1  g536(.A1(new_n567_), .A2(new_n444_), .A3(new_n581_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G85gat), .B1(new_n740_), .B2(new_n396_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n707_), .A2(new_n567_), .A3(new_n643_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n742_), .A2(new_n462_), .A3(new_n334_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1336gat));
  OAI21_X1  g543(.A(G92gat), .B1(new_n740_), .B2(new_n390_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n742_), .A2(new_n463_), .A3(new_n616_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(G1337gat));
  NAND4_X1  g546(.A1(new_n742_), .A2(new_n249_), .A3(new_n448_), .A4(new_n453_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n739_), .A2(new_n249_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(G99gat), .ZN(new_n751_));
  AOI211_X1 g550(.A(KEYINPUT109), .B(new_n472_), .C1(new_n739_), .C2(new_n249_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g553(.A(KEYINPUT110), .B(KEYINPUT53), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT52), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(G106gat), .C1(new_n740_), .C2(new_n382_), .ZN(new_n758_));
  AOI211_X1 g557(.A(new_n382_), .B(new_n738_), .C1(new_n656_), .C2(new_n657_), .ZN(new_n759_));
  OAI21_X1  g558(.A(KEYINPUT52), .B1(new_n759_), .B2(new_n449_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT111), .ZN(new_n762_));
  NAND4_X1  g561(.A1(new_n742_), .A2(new_n381_), .A3(new_n450_), .A4(new_n452_), .ZN(new_n763_));
  AND3_X1   g562(.A1(new_n761_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n762_), .B1(new_n761_), .B2(new_n763_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n756_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT111), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n761_), .A2(new_n762_), .A3(new_n763_), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n769_), .A3(new_n755_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n766_), .A2(new_n770_), .ZN(G1339gat));
  NOR3_X1   g570(.A1(new_n398_), .A2(new_n250_), .A3(new_n396_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n773_), .A2(KEYINPUT59), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT54), .B1(new_n585_), .B2(new_n432_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT54), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n582_), .A2(new_n776_), .A3(new_n444_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n414_), .A2(new_n415_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n429_), .B1(new_n422_), .B2(new_n416_), .ZN(new_n780_));
  AOI22_X1  g579(.A1(new_n426_), .A2(new_n429_), .B1(new_n779_), .B2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n562_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784_));
  AND2_X1   g583(.A1(new_n548_), .A2(new_n549_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n548_), .A2(new_n549_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n784_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n537_), .A2(new_n789_), .ZN(new_n790_));
  AND4_X1   g589(.A1(new_n538_), .A2(new_n543_), .A3(new_n547_), .A4(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n791_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n537_), .A2(new_n784_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n538_), .A2(new_n543_), .A3(new_n547_), .A4(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n790_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n792_), .A2(new_n796_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n787_), .A2(new_n788_), .A3(new_n797_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT55), .B1(new_n539_), .B2(new_n550_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n791_), .B1(new_n795_), .B2(new_n794_), .ZN(new_n800_));
  OAI21_X1  g599(.A(KEYINPUT113), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n798_), .A2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT56), .B1(new_n802_), .B2(new_n559_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT56), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n804_), .B(new_n560_), .C1(new_n798_), .C2(new_n801_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n783_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT58), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n518_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT117), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n806_), .A2(new_n807_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n651_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT117), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n811_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n788_), .B1(new_n787_), .B2(new_n797_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n799_), .A2(new_n800_), .A3(KEYINPUT113), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT56), .B(new_n559_), .C1(new_n815_), .C2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT115), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n559_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n818_), .A2(new_n804_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n820_), .A2(KEYINPUT114), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n560_), .B1(new_n798_), .B2(new_n801_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n821_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n819_), .A2(new_n823_), .A3(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n432_), .A2(new_n562_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n827_), .A2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n563_), .A2(new_n781_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n599_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n810_), .A2(new_n814_), .B1(new_n832_), .B2(KEYINPUT57), .ZN(new_n833_));
  INV_X1    g632(.A(new_n831_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n827_), .B2(new_n829_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT116), .B1(new_n835_), .B2(new_n599_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT116), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n825_), .B1(new_n802_), .B2(new_n559_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n838_), .A2(new_n822_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n828_), .B1(new_n839_), .B2(new_n826_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n837_), .B(new_n600_), .C1(new_n840_), .C2(new_n834_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n836_), .A2(new_n841_), .A3(new_n842_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n597_), .B1(new_n833_), .B2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n778_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  AOI211_X1 g645(.A(KEYINPUT119), .B(new_n597_), .C1(new_n833_), .C2(new_n843_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n774_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n778_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n810_), .A2(new_n814_), .A3(KEYINPUT118), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n820_), .A2(new_n804_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n782_), .B1(new_n852_), .B2(new_n817_), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n813_), .B(new_n518_), .C1(new_n853_), .C2(KEYINPUT58), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(KEYINPUT58), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n813_), .B1(new_n808_), .B2(new_n518_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n851_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n832_), .A2(KEYINPUT57), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n843_), .A2(new_n850_), .A3(new_n858_), .A4(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n849_), .B1(new_n860_), .B2(new_n581_), .ZN(new_n861_));
  OAI21_X1  g660(.A(KEYINPUT59), .B1(new_n861_), .B2(new_n773_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n432_), .A2(G113gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT120), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n848_), .A2(new_n862_), .A3(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n860_), .A2(new_n581_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n778_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n867_), .A2(new_n432_), .A3(new_n772_), .ZN(new_n868_));
  INV_X1    g667(.A(G113gat), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n865_), .A2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT121), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n865_), .A2(KEYINPUT121), .A3(new_n870_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1340gat));
  NAND3_X1  g674(.A1(new_n848_), .A2(new_n567_), .A3(new_n862_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(G120gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n867_), .A2(new_n772_), .ZN(new_n878_));
  INV_X1    g677(.A(G120gat), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n596_), .B2(KEYINPUT60), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(KEYINPUT60), .B2(new_n879_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n877_), .B1(new_n878_), .B2(new_n881_), .ZN(G1341gat));
  INV_X1    g681(.A(G127gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n878_), .B2(new_n581_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT122), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886_));
  OAI211_X1 g685(.A(new_n886_), .B(new_n883_), .C1(new_n878_), .C2(new_n581_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n848_), .A2(new_n862_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n581_), .A2(new_n883_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n885_), .A2(new_n887_), .B1(new_n888_), .B2(new_n889_), .ZN(G1342gat));
  NAND2_X1  g689(.A1(new_n518_), .A2(G134gat), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(KEYINPUT123), .ZN(new_n892_));
  INV_X1    g691(.A(G134gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n867_), .A2(new_n599_), .A3(new_n772_), .ZN(new_n894_));
  AOI22_X1  g693(.A1(new_n888_), .A2(new_n892_), .B1(new_n893_), .B2(new_n894_), .ZN(G1343gat));
  NOR4_X1   g694(.A1(new_n616_), .A2(new_n249_), .A3(new_n382_), .A4(new_n396_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n861_), .A2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n432_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n567_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g701(.A(KEYINPUT61), .B(G155gat), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n867_), .A2(new_n896_), .ZN(new_n904_));
  OAI21_X1  g703(.A(KEYINPUT124), .B1(new_n904_), .B2(new_n581_), .ZN(new_n905_));
  NOR4_X1   g704(.A1(new_n861_), .A2(KEYINPUT124), .A3(new_n581_), .A4(new_n897_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n903_), .B1(new_n905_), .B2(new_n907_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT124), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n909_), .B1(new_n898_), .B2(new_n597_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n903_), .ZN(new_n911_));
  NOR3_X1   g710(.A1(new_n910_), .A2(new_n906_), .A3(new_n911_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n908_), .A2(new_n912_), .ZN(G1346gat));
  OR3_X1    g712(.A1(new_n904_), .A2(G162gat), .A3(new_n600_), .ZN(new_n914_));
  OAI21_X1  g713(.A(G162gat), .B1(new_n904_), .B2(new_n651_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1347gat));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n616_), .A2(new_n249_), .A3(new_n396_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n381_), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n432_), .B(new_n919_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n920_));
  INV_X1    g719(.A(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n917_), .B1(new_n921_), .B2(new_n216_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n214_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n920_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n922_), .A2(new_n923_), .A3(new_n924_), .ZN(G1348gat));
  NAND2_X1  g724(.A1(new_n867_), .A2(new_n382_), .ZN(new_n926_));
  NOR4_X1   g725(.A1(new_n926_), .A2(new_n222_), .A3(new_n596_), .A4(new_n918_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n567_), .B(new_n919_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n929_));
  INV_X1    g728(.A(new_n929_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n928_), .B1(new_n930_), .B2(G176gat), .ZN(new_n931_));
  NAND3_X1  g730(.A1(new_n929_), .A2(KEYINPUT125), .A3(new_n222_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n927_), .B1(new_n931_), .B2(new_n932_), .ZN(G1349gat));
  OR3_X1    g732(.A1(new_n926_), .A2(new_n581_), .A3(new_n918_), .ZN(new_n934_));
  OR2_X1    g733(.A1(new_n846_), .A2(new_n847_), .ZN(new_n935_));
  AND2_X1   g734(.A1(new_n935_), .A2(new_n919_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n581_), .B1(new_n226_), .B2(new_n230_), .ZN(new_n937_));
  AOI22_X1  g736(.A1(new_n207_), .A2(new_n934_), .B1(new_n936_), .B2(new_n937_), .ZN(G1350gat));
  NAND4_X1  g737(.A1(new_n935_), .A2(new_n274_), .A3(new_n599_), .A4(new_n919_), .ZN(new_n939_));
  OAI211_X1 g738(.A(new_n518_), .B(new_n919_), .C1(new_n846_), .C2(new_n847_), .ZN(new_n940_));
  INV_X1    g739(.A(KEYINPUT126), .ZN(new_n941_));
  AND3_X1   g740(.A1(new_n940_), .A2(new_n941_), .A3(G190gat), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n940_), .B2(G190gat), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n939_), .B1(new_n942_), .B2(new_n943_), .ZN(G1351gat));
  NAND3_X1  g743(.A1(new_n250_), .A2(new_n616_), .A3(new_n391_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n861_), .A2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(new_n432_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(G197gat), .ZN(G1352gat));
  NOR3_X1   g747(.A1(new_n861_), .A2(new_n596_), .A3(new_n945_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n949_), .B1(KEYINPUT127), .B2(new_n258_), .ZN(new_n950_));
  XNOR2_X1  g749(.A(KEYINPUT127), .B(G204gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n949_), .B2(new_n951_), .ZN(G1353gat));
  NOR3_X1   g751(.A1(new_n861_), .A2(new_n581_), .A3(new_n945_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n953_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954_));
  XOR2_X1   g753(.A(KEYINPUT63), .B(G211gat), .Z(new_n955_));
  AOI21_X1  g754(.A(new_n954_), .B1(new_n953_), .B2(new_n955_), .ZN(G1354gat));
  INV_X1    g755(.A(G218gat), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n946_), .A2(new_n957_), .A3(new_n599_), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n861_), .A2(new_n651_), .A3(new_n945_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n959_), .B2(new_n957_), .ZN(G1355gat));
endmodule


