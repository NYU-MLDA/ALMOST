//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 1 1 0 1 1 0 1 0 0 1 1 1 1 0 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n918_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n931_;
  NOR2_X1   g000(.A1(KEYINPUT71), .A2(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XOR2_X1   g002(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n204_));
  INV_X1    g003(.A(KEYINPUT7), .ZN(new_n205_));
  INV_X1    g004(.A(G99gat), .ZN(new_n206_));
  INV_X1    g005(.A(G106gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT6), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n213_));
  NAND4_X1  g012(.A1(new_n208_), .A2(new_n211_), .A3(new_n212_), .A4(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G85gat), .A2(G92gat), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n214_), .A2(KEYINPUT66), .A3(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT8), .ZN(new_n219_));
  NAND3_X1  g018(.A1(new_n218_), .A2(KEYINPUT67), .A3(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n216_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT9), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT9), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n216_), .A2(new_n221_), .A3(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n215_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT65), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n206_), .A2(KEYINPUT10), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT10), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n229_), .A2(G99gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(G106gat), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n211_), .A2(new_n212_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n223_), .A2(new_n234_), .A3(new_n215_), .A4(new_n225_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n227_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n218_), .A2(KEYINPUT67), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n214_), .A2(new_n238_), .A3(new_n217_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n239_), .A2(KEYINPUT8), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n220_), .B(new_n236_), .C1(new_n237_), .C2(new_n240_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G57gat), .B(G64gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT11), .ZN(new_n243_));
  XNOR2_X1  g042(.A(G71gat), .B(G78gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  XOR2_X1   g044(.A(new_n242_), .B(KEYINPUT11), .Z(new_n246_));
  OAI21_X1  g045(.A(new_n245_), .B1(new_n246_), .B2(new_n244_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n204_), .B1(new_n241_), .B2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n241_), .A2(new_n247_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n236_), .A2(KEYINPUT68), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n252_));
  NAND4_X1  g051(.A1(new_n227_), .A2(new_n252_), .A3(new_n233_), .A4(new_n235_), .ZN(new_n253_));
  AND2_X1   g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n218_), .A2(KEYINPUT67), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT8), .A3(new_n239_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n220_), .ZN(new_n257_));
  OAI211_X1 g056(.A(KEYINPUT12), .B(new_n247_), .C1(new_n254_), .C2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G230gat), .A2(G233gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n250_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n241_), .A2(new_n247_), .ZN(new_n261_));
  OAI211_X1 g060(.A(G230gat), .B(G233gat), .C1(new_n261_), .C2(new_n249_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT5), .B(G176gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n263_), .B(G204gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G120gat), .B(G148gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n264_), .B(new_n265_), .Z(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n260_), .A2(new_n262_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n267_), .B1(new_n260_), .B2(new_n262_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n270_));
  NOR3_X1   g069(.A1(new_n268_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n260_), .A2(new_n262_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n272_), .A2(new_n266_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n260_), .A2(new_n262_), .A3(new_n267_), .ZN(new_n274_));
  AOI21_X1  g073(.A(KEYINPUT70), .B1(new_n273_), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n203_), .B1(new_n271_), .B2(new_n275_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n270_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n273_), .A2(KEYINPUT70), .A3(new_n274_), .ZN(new_n278_));
  XOR2_X1   g077(.A(KEYINPUT71), .B(KEYINPUT13), .Z(new_n279_));
  INV_X1    g078(.A(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n277_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n276_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G29gat), .B(G36gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G43gat), .B(G50gat), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n286_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n284_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n287_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT15), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G15gat), .B(G22gat), .ZN(new_n293_));
  INV_X1    g092(.A(G1gat), .ZN(new_n294_));
  INV_X1    g093(.A(G8gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(KEYINPUT14), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G8gat), .ZN(new_n298_));
  OR2_X1    g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n298_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n292_), .A2(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G229gat), .A2(G233gat), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n299_), .A2(new_n300_), .A3(new_n287_), .A4(new_n289_), .ZN(new_n304_));
  AND3_X1   g103(.A1(new_n302_), .A2(new_n303_), .A3(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n303_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n290_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(new_n304_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n307_), .A2(KEYINPUT77), .A3(new_n304_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n305_), .B1(new_n306_), .B2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT78), .B(G169gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(G197gat), .ZN(new_n315_));
  XOR2_X1   g114(.A(G113gat), .B(G141gat), .Z(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  XOR2_X1   g116(.A(new_n313_), .B(new_n317_), .Z(new_n318_));
  NOR2_X1   g117(.A1(new_n283_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT27), .ZN(new_n321_));
  NAND2_X1  g120(.A1(G183gat), .A2(G190gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT82), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT82), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n324_), .A2(G183gat), .A3(G190gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(KEYINPUT23), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT84), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n328_), .B1(new_n322_), .B2(KEYINPUT23), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n330_), .A2(KEYINPUT84), .A3(G183gat), .A4(G190gat), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(new_n329_), .A3(new_n331_), .ZN(new_n332_));
  NOR2_X1   g131(.A1(G183gat), .A2(G190gat), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n332_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT22), .B(G169gat), .ZN(new_n336_));
  INV_X1    g135(.A(G176gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n335_), .A2(new_n341_), .ZN(new_n342_));
  XOR2_X1   g141(.A(G197gat), .B(G204gat), .Z(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(KEYINPUT21), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G197gat), .B(G204gat), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT21), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G211gat), .B(G218gat), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n344_), .A2(new_n347_), .A3(new_n348_), .ZN(new_n349_));
  OR3_X1    g148(.A1(new_n345_), .A2(new_n348_), .A3(new_n346_), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n323_), .A2(new_n325_), .A3(new_n330_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n352_), .A2(KEYINPUT83), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n322_), .A2(KEYINPUT23), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT83), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n323_), .A2(new_n325_), .A3(new_n355_), .A4(new_n330_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n353_), .A2(new_n354_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT80), .ZN(new_n358_));
  INV_X1    g157(.A(G190gat), .ZN(new_n359_));
  OAI21_X1  g158(.A(KEYINPUT79), .B1(new_n359_), .B2(KEYINPUT26), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT79), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT26), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n361_), .A2(new_n362_), .A3(G190gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n360_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n359_), .A2(KEYINPUT26), .ZN(new_n365_));
  AND2_X1   g164(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n366_));
  NOR2_X1   g165(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n365_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n358_), .B1(new_n364_), .B2(new_n368_), .ZN(new_n369_));
  OR2_X1    g168(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n370_), .A2(new_n371_), .B1(KEYINPUT26), .B2(new_n359_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n372_), .A2(KEYINPUT80), .A3(new_n363_), .A4(new_n360_), .ZN(new_n373_));
  NOR2_X1   g172(.A1(G169gat), .A2(G176gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT81), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT81), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n376_), .B1(G169gat), .B2(G176gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT24), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n379_), .B1(G169gat), .B2(G176gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  NAND4_X1  g180(.A1(new_n357_), .A2(new_n369_), .A3(new_n373_), .A4(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n375_), .A2(new_n379_), .A3(new_n377_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  OAI211_X1 g183(.A(new_n342_), .B(new_n351_), .C1(new_n382_), .C2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n349_), .A2(new_n350_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n380_), .A2(KEYINPUT98), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT98), .ZN(new_n388_));
  INV_X1    g187(.A(new_n339_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n388_), .B1(new_n389_), .B2(new_n379_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n387_), .A2(new_n378_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n362_), .A2(G190gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n372_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n374_), .A2(new_n379_), .ZN(new_n394_));
  AND4_X1   g193(.A1(new_n332_), .A2(new_n391_), .A3(new_n393_), .A4(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n340_), .B1(new_n357_), .B2(new_n334_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n386_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n385_), .A2(new_n397_), .A3(KEYINPUT20), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G226gat), .A2(G233gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n398_), .A2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT99), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n398_), .A2(KEYINPUT99), .A3(new_n402_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(G8gat), .B(G36gat), .ZN(new_n408_));
  INV_X1    g207(.A(G92gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n408_), .B(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT18), .B(G64gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n410_), .B(new_n411_), .Z(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT100), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n373_), .A2(new_n369_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n415_), .A2(new_n383_), .A3(new_n357_), .A4(new_n381_), .ZN(new_n416_));
  AOI211_X1 g215(.A(new_n414_), .B(new_n351_), .C1(new_n416_), .C2(new_n342_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n342_), .B1(new_n382_), .B2(new_n384_), .ZN(new_n418_));
  AOI21_X1  g217(.A(KEYINPUT100), .B1(new_n418_), .B2(new_n386_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n417_), .A2(new_n419_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n395_), .A2(new_n396_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n421_), .A2(new_n351_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n420_), .A2(KEYINPUT20), .A3(new_n401_), .A4(new_n422_), .ZN(new_n423_));
  AND3_X1   g222(.A1(new_n407_), .A2(new_n413_), .A3(new_n423_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n413_), .B1(new_n407_), .B2(new_n423_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n321_), .B1(new_n424_), .B2(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(G113gat), .B(G120gat), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n427_), .B(G134gat), .ZN(new_n428_));
  XNOR2_X1  g227(.A(KEYINPUT88), .B(G127gat), .ZN(new_n429_));
  OR2_X1    g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n428_), .A2(new_n429_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OR2_X1    g231(.A1(G155gat), .A2(G162gat), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G155gat), .A2(G162gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT92), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G141gat), .A2(G148gat), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT91), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT3), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT91), .B1(new_n439_), .B2(KEYINPUT92), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n438_), .A2(new_n439_), .B1(new_n436_), .B2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G141gat), .A2(G148gat), .ZN(new_n442_));
  XOR2_X1   g241(.A(new_n442_), .B(KEYINPUT2), .Z(new_n443_));
  OAI211_X1 g242(.A(new_n433_), .B(new_n434_), .C1(new_n441_), .C2(new_n443_), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n434_), .A2(KEYINPUT1), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n434_), .A2(KEYINPUT1), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n433_), .A3(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n436_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n447_), .A2(new_n448_), .A3(new_n442_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n432_), .A2(new_n450_), .ZN(new_n451_));
  NAND4_X1  g250(.A1(new_n430_), .A2(new_n444_), .A3(new_n449_), .A4(new_n431_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(KEYINPUT4), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT4), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n432_), .A2(new_n454_), .A3(new_n450_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G225gat), .A2(G233gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(KEYINPUT101), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n453_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n451_), .A2(new_n452_), .A3(new_n456_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  XOR2_X1   g259(.A(G57gat), .B(G85gat), .Z(new_n461_));
  XNOR2_X1  g260(.A(G1gat), .B(G29gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(KEYINPUT102), .B(KEYINPUT0), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n460_), .A2(new_n466_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n458_), .A2(new_n459_), .A3(new_n465_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n407_), .A2(new_n423_), .A3(new_n413_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n398_), .A2(new_n402_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT104), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n421_), .A2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(KEYINPUT104), .B1(new_n395_), .B2(new_n396_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n351_), .A3(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n420_), .A2(KEYINPUT20), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n472_), .B1(new_n477_), .B2(new_n402_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n471_), .B(KEYINPUT27), .C1(new_n478_), .C2(new_n413_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n426_), .A2(new_n470_), .A3(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n351_), .B1(new_n450_), .B2(KEYINPUT29), .ZN(new_n481_));
  INV_X1    g280(.A(G233gat), .ZN(new_n482_));
  AND2_X1   g281(.A1(new_n482_), .A2(KEYINPUT93), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n482_), .A2(KEYINPUT93), .ZN(new_n484_));
  OAI21_X1  g283(.A(G228gat), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NOR2_X1   g284(.A1(new_n481_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT95), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n481_), .A2(new_n485_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT94), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G78gat), .B(G106gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  OR3_X1    g292(.A1(new_n450_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n494_));
  OAI21_X1  g293(.A(KEYINPUT28), .B1(new_n450_), .B2(KEYINPUT29), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G22gat), .B(G50gat), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n496_), .A2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT96), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n496_), .A2(new_n498_), .ZN(new_n502_));
  OR3_X1    g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  OAI21_X1  g302(.A(new_n501_), .B1(new_n500_), .B2(new_n502_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n492_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n488_), .A2(new_n490_), .A3(new_n505_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n493_), .A2(new_n503_), .A3(new_n504_), .A4(new_n506_), .ZN(new_n507_));
  NOR3_X1   g306(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n508_));
  AND3_X1   g307(.A1(new_n488_), .A2(new_n490_), .A3(new_n505_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n505_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n507_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n480_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n507_), .A2(new_n511_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n453_), .A2(new_n456_), .A3(new_n455_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n451_), .A2(new_n452_), .A3(new_n457_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n466_), .A3(new_n516_), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT103), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n468_), .B(KEYINPUT33), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n407_), .A2(new_n423_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(new_n412_), .ZN(new_n521_));
  NAND4_X1  g320(.A1(new_n518_), .A2(new_n519_), .A3(new_n521_), .A4(new_n471_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n413_), .A2(KEYINPUT32), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n407_), .A2(new_n423_), .A3(new_n523_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n469_), .B(new_n524_), .C1(new_n478_), .C2(new_n523_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n514_), .A2(new_n522_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT85), .B(KEYINPUT30), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n342_), .B(new_n528_), .C1(new_n382_), .C2(new_n384_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n528_), .B1(new_n416_), .B2(new_n342_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n527_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n528_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n418_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(KEYINPUT87), .A3(new_n529_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G15gat), .B(G43gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G71gat), .B(G99gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G227gat), .A2(G233gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT86), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n538_), .B(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n532_), .A2(new_n535_), .A3(new_n542_), .ZN(new_n543_));
  NAND4_X1  g342(.A1(new_n534_), .A2(KEYINPUT87), .A3(new_n529_), .A4(new_n541_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT90), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n547_));
  XOR2_X1   g346(.A(new_n432_), .B(new_n547_), .Z(new_n548_));
  INV_X1    g347(.A(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n546_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT90), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n543_), .A2(new_n544_), .A3(new_n551_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n551_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n550_), .B1(new_n549_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n513_), .A2(new_n526_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT105), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n555_), .B1(new_n480_), .B2(new_n512_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT105), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n560_), .A3(new_n526_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n426_), .A2(new_n479_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n563_), .A2(new_n470_), .A3(new_n555_), .A4(new_n514_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n320_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT76), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n290_), .B(KEYINPUT15), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n256_), .A2(new_n220_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n251_), .A2(new_n253_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n567_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  XOR2_X1   g369(.A(KEYINPUT72), .B(KEYINPUT34), .Z(new_n571_));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n571_), .B(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT35), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n575_), .B(KEYINPUT73), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n570_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n573_), .A2(new_n574_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n578_), .B1(new_n241_), .B2(new_n290_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n566_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n581_));
  NOR4_X1   g380(.A1(new_n570_), .A2(new_n579_), .A3(new_n576_), .A4(KEYINPUT76), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT74), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n579_), .B1(new_n570_), .B2(new_n584_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n585_), .B1(new_n584_), .B2(new_n570_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n576_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G190gat), .B(G218gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(G162gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT75), .B(G134gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  OR2_X1    g393(.A1(new_n592_), .A2(new_n593_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n588_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  NAND4_X1  g395(.A1(new_n583_), .A2(new_n587_), .A3(new_n593_), .A4(new_n592_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT37), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n596_), .A2(KEYINPUT37), .A3(new_n597_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G231gat), .A2(G233gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n301_), .B(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n604_), .B(new_n247_), .Z(new_n605_));
  XNOR2_X1  g404(.A(G127gat), .B(G155gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(G211gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT16), .B(G183gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n609_), .A2(KEYINPUT17), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n605_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n609_), .B(KEYINPUT17), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n605_), .A2(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n602_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n565_), .A2(new_n616_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n617_), .A2(G1gat), .A3(new_n470_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(KEYINPUT106), .B(KEYINPUT38), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n565_), .A2(KEYINPUT107), .A3(new_n614_), .A4(new_n598_), .ZN(new_n621_));
  AND4_X1   g420(.A1(new_n560_), .A2(new_n513_), .A3(new_n556_), .A4(new_n526_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n560_), .B1(new_n559_), .B2(new_n526_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n564_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n624_), .A2(new_n319_), .A3(new_n614_), .A4(new_n598_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT107), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n470_), .B1(new_n621_), .B2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n620_), .B1(new_n628_), .B2(new_n294_), .ZN(G1324gat));
  OAI21_X1  g428(.A(G8gat), .B1(new_n625_), .B2(new_n563_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n630_), .A2(KEYINPUT108), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT108), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n632_), .B(G8gat), .C1(new_n625_), .C2(new_n563_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n563_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n565_), .A2(new_n295_), .A3(new_n637_), .A4(new_n616_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n631_), .A2(KEYINPUT39), .A3(new_n633_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n636_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT40), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n636_), .A2(KEYINPUT40), .A3(new_n638_), .A4(new_n639_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1325gat));
  INV_X1    g443(.A(G15gat), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n565_), .A2(new_n645_), .A3(new_n555_), .A4(new_n616_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n625_), .A2(new_n626_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n625_), .A2(new_n626_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n555_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(KEYINPUT41), .B1(new_n649_), .B2(G15gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n556_), .B1(new_n621_), .B2(new_n627_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n652_));
  NOR3_X1   g451(.A1(new_n651_), .A2(new_n652_), .A3(new_n645_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n646_), .B1(new_n650_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT109), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(KEYINPUT109), .B(new_n646_), .C1(new_n650_), .C2(new_n653_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(G1326gat));
  OR3_X1    g457(.A1(new_n617_), .A2(G22gat), .A3(new_n514_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n512_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT42), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n660_), .A2(new_n661_), .A3(G22gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n661_), .B1(new_n660_), .B2(G22gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n662_), .B2(new_n663_), .ZN(G1327gat));
  INV_X1    g463(.A(KEYINPUT112), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n624_), .A2(new_n319_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n598_), .A2(new_n614_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n665_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n565_), .A2(KEYINPUT112), .A3(new_n667_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n671_), .A2(G29gat), .A3(new_n470_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT111), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n624_), .A2(new_n602_), .ZN(new_n674_));
  XOR2_X1   g473(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n624_), .A2(KEYINPUT110), .A3(KEYINPUT43), .A4(new_n602_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n676_), .A2(new_n319_), .A3(new_n615_), .A4(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n679_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n680_), .A2(new_n469_), .A3(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n673_), .B1(new_n682_), .B2(G29gat), .ZN(new_n683_));
  INV_X1    g482(.A(new_n681_), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n469_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n673_), .B(G29gat), .C1(new_n684_), .C2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n672_), .B1(new_n683_), .B2(new_n687_), .ZN(G1328gat));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n689_));
  INV_X1    g488(.A(G36gat), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n563_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n680_), .B2(new_n691_), .ZN(new_n692_));
  NAND4_X1  g491(.A1(new_n669_), .A2(new_n670_), .A3(new_n690_), .A4(new_n637_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT45), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n689_), .B1(new_n692_), .B2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n681_), .A2(new_n637_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n678_), .A2(new_n679_), .ZN(new_n698_));
  OAI21_X1  g497(.A(G36gat), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n693_), .B(KEYINPUT45), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n699_), .A2(KEYINPUT46), .A3(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n696_), .A2(new_n701_), .ZN(G1329gat));
  NAND3_X1  g501(.A1(new_n669_), .A2(new_n670_), .A3(new_n555_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT113), .ZN(new_n704_));
  INV_X1    g503(.A(G43gat), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n704_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n681_), .A2(new_n555_), .ZN(new_n708_));
  OAI21_X1  g507(.A(G43gat), .B1(new_n678_), .B2(new_n679_), .ZN(new_n709_));
  OAI22_X1  g508(.A1(new_n706_), .A2(new_n707_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT47), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712_));
  OAI221_X1 g511(.A(new_n712_), .B1(new_n708_), .B2(new_n709_), .C1(new_n707_), .C2(new_n706_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1330gat));
  NOR3_X1   g513(.A1(new_n684_), .A2(new_n698_), .A3(new_n514_), .ZN(new_n715_));
  INV_X1    g514(.A(G50gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n514_), .A2(G50gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT114), .ZN(new_n718_));
  OAI22_X1  g517(.A1(new_n715_), .A2(new_n716_), .B1(new_n671_), .B2(new_n718_), .ZN(G1331gat));
  INV_X1    g518(.A(new_n318_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n282_), .A2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n722_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(new_n616_), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(G57gat), .B1(new_n725_), .B2(new_n469_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT115), .ZN(new_n727_));
  INV_X1    g526(.A(G57gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n596_), .A2(new_n597_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n730_), .A2(new_n615_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n723_), .A2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n728_), .B1(new_n469_), .B2(new_n727_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n726_), .B1(new_n729_), .B2(new_n734_), .ZN(G1332gat));
  OAI21_X1  g534(.A(G64gat), .B1(new_n732_), .B2(new_n563_), .ZN(new_n736_));
  XNOR2_X1  g535(.A(new_n736_), .B(KEYINPUT48), .ZN(new_n737_));
  OR2_X1    g536(.A1(new_n563_), .A2(G64gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n737_), .B1(new_n724_), .B2(new_n738_), .ZN(G1333gat));
  OR3_X1    g538(.A1(new_n724_), .A2(G71gat), .A3(new_n556_), .ZN(new_n740_));
  OAI21_X1  g539(.A(G71gat), .B1(new_n732_), .B2(new_n556_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(KEYINPUT49), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(KEYINPUT49), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n740_), .B1(new_n742_), .B2(new_n743_), .ZN(G1334gat));
  OR3_X1    g543(.A1(new_n724_), .A2(G78gat), .A3(new_n514_), .ZN(new_n745_));
  OAI21_X1  g544(.A(G78gat), .B1(new_n732_), .B2(new_n514_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(KEYINPUT50), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n746_), .A2(KEYINPUT50), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n745_), .B1(new_n747_), .B2(new_n748_), .ZN(G1335gat));
  NAND2_X1  g548(.A1(new_n723_), .A2(new_n667_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(G85gat), .B1(new_n751_), .B2(new_n469_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n722_), .A2(new_n614_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n676_), .A2(new_n677_), .A3(new_n753_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n754_), .A2(new_n470_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n752_), .B1(new_n755_), .B2(G85gat), .ZN(G1336gat));
  NOR3_X1   g555(.A1(new_n754_), .A2(new_n409_), .A3(new_n563_), .ZN(new_n757_));
  AOI21_X1  g556(.A(G92gat), .B1(new_n751_), .B2(new_n637_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n754_), .B2(new_n556_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n556_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n751_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  XNOR2_X1  g562(.A(KEYINPUT116), .B(KEYINPUT51), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n763_), .B(new_n764_), .ZN(G1338gat));
  NAND4_X1  g564(.A1(new_n676_), .A2(new_n512_), .A3(new_n677_), .A4(new_n753_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT117), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT52), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n766_), .A2(G106gat), .A3(new_n768_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n767_), .A2(KEYINPUT52), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n751_), .A2(new_n207_), .A3(new_n512_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n770_), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n766_), .A2(G106gat), .A3(new_n773_), .A4(new_n768_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n771_), .A2(new_n772_), .A3(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT53), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777_));
  NAND4_X1  g576(.A1(new_n771_), .A2(new_n777_), .A3(new_n772_), .A4(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(G1339gat));
  AND3_X1   g578(.A1(new_n277_), .A2(new_n278_), .A3(new_n280_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n202_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n781_));
  OAI211_X1 g580(.A(new_n318_), .B(new_n614_), .C1(new_n780_), .C2(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT118), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n282_), .A2(KEYINPUT118), .A3(new_n318_), .A4(new_n614_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n602_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787_));
  XNOR2_X1  g586(.A(new_n786_), .B(new_n787_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n259_), .B1(new_n250_), .B2(new_n258_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n260_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n250_), .A2(new_n258_), .A3(KEYINPUT55), .A4(new_n259_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n793_), .A2(new_n266_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT56), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n267_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT119), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n795_), .A2(new_n799_), .A3(new_n720_), .A4(new_n274_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT120), .B1(new_n302_), .B2(new_n304_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n801_), .A2(new_n303_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n302_), .A2(KEYINPUT120), .A3(new_n304_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n317_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n312_), .A2(new_n303_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n804_), .A2(new_n805_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n806_), .B1(new_n271_), .B2(new_n275_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n800_), .A2(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n598_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n808_), .A2(KEYINPUT57), .A3(new_n598_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n797_), .B(KEYINPUT56), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n806_), .A2(new_n274_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT121), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n806_), .A2(new_n816_), .A3(new_n274_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n813_), .A2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n813_), .A2(new_n818_), .A3(KEYINPUT58), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n821_), .A2(new_n602_), .A3(new_n822_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n811_), .A2(KEYINPUT122), .A3(new_n812_), .A4(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n615_), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT57), .B1(new_n808_), .B2(new_n598_), .ZN(new_n826_));
  AOI211_X1 g625(.A(new_n810_), .B(new_n730_), .C1(new_n800_), .C2(new_n807_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT122), .B1(new_n828_), .B2(new_n823_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n788_), .B1(new_n825_), .B2(new_n829_), .ZN(new_n830_));
  NOR4_X1   g629(.A1(new_n637_), .A2(new_n556_), .A3(new_n470_), .A4(new_n512_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(G113gat), .B1(new_n832_), .B2(new_n720_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(KEYINPUT59), .A3(new_n831_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT123), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n831_), .A2(new_n835_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n831_), .A2(new_n835_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n614_), .B1(new_n828_), .B2(new_n823_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n784_), .A2(new_n785_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n602_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n787_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n841_));
  AOI211_X1 g640(.A(KEYINPUT54), .B(new_n602_), .C1(new_n784_), .C2(new_n785_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n836_), .B(new_n837_), .C1(new_n838_), .C2(new_n843_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT59), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n834_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n318_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n833_), .B1(new_n849_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g649(.A(KEYINPUT124), .ZN(new_n851_));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n852_), .B1(new_n847_), .B2(new_n283_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n282_), .B2(KEYINPUT60), .ZN(new_n854_));
  OR2_X1    g653(.A1(new_n852_), .A2(KEYINPUT60), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n832_), .A2(new_n854_), .A3(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n851_), .B1(new_n853_), .B2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n282_), .B1(new_n834_), .B2(new_n846_), .ZN(new_n859_));
  OAI211_X1 g658(.A(KEYINPUT124), .B(new_n856_), .C1(new_n859_), .C2(new_n852_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(G1341gat));
  AOI21_X1  g660(.A(G127gat), .B1(new_n832_), .B2(new_n614_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n848_), .A2(new_n615_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n863_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g663(.A(G134gat), .B1(new_n832_), .B2(new_n730_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n848_), .A2(new_n840_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(G134gat), .ZN(G1343gat));
  AND2_X1   g666(.A1(new_n830_), .A2(new_n512_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n637_), .A2(new_n555_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n868_), .A2(new_n469_), .A3(new_n869_), .ZN(new_n870_));
  OR3_X1    g669(.A1(new_n870_), .A2(G141gat), .A3(new_n318_), .ZN(new_n871_));
  OAI21_X1  g670(.A(G141gat), .B1(new_n870_), .B2(new_n318_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n871_), .A2(new_n872_), .ZN(G1344gat));
  OR3_X1    g672(.A1(new_n870_), .A2(G148gat), .A3(new_n282_), .ZN(new_n874_));
  OAI21_X1  g673(.A(G148gat), .B1(new_n870_), .B2(new_n282_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(G1345gat));
  AND2_X1   g675(.A1(new_n868_), .A2(new_n469_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT61), .B(G155gat), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n877_), .A2(new_n614_), .A3(new_n869_), .A4(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n878_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n880_), .B1(new_n870_), .B2(new_n615_), .ZN(new_n881_));
  AND2_X1   g680(.A1(new_n879_), .A2(new_n881_), .ZN(G1346gat));
  INV_X1    g681(.A(G162gat), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n870_), .A2(new_n883_), .A3(new_n840_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n877_), .A2(new_n730_), .A3(new_n869_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n883_), .B2(new_n885_), .ZN(G1347gat));
  OR2_X1    g685(.A1(new_n838_), .A2(new_n843_), .ZN(new_n887_));
  NOR4_X1   g686(.A1(new_n556_), .A2(new_n563_), .A3(new_n469_), .A4(new_n512_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(G169gat), .B1(new_n889_), .B2(new_n318_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT62), .ZN(new_n891_));
  OR2_X1    g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n889_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n893_), .A2(new_n720_), .A3(new_n336_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n890_), .A2(new_n891_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n892_), .A2(new_n894_), .A3(new_n895_), .ZN(G1348gat));
  AND2_X1   g695(.A1(new_n830_), .A2(new_n888_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n897_), .A2(G176gat), .A3(new_n283_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT125), .ZN(new_n899_));
  AND2_X1   g698(.A1(new_n898_), .A2(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n898_), .A2(new_n899_), .ZN(new_n901_));
  AOI21_X1  g700(.A(G176gat), .B1(new_n893_), .B2(new_n283_), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(G1349gat));
  NAND3_X1  g702(.A1(new_n897_), .A2(KEYINPUT126), .A3(new_n614_), .ZN(new_n904_));
  INV_X1    g703(.A(G183gat), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n830_), .A2(new_n614_), .A3(new_n888_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT126), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n906_), .A2(new_n907_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n904_), .A2(new_n905_), .A3(new_n908_), .ZN(new_n909_));
  NAND4_X1  g708(.A1(new_n893_), .A2(new_n370_), .A3(new_n371_), .A4(new_n614_), .ZN(new_n910_));
  AND2_X1   g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1350gat));
  OAI21_X1  g710(.A(G190gat), .B1(new_n889_), .B2(new_n840_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n730_), .A2(new_n365_), .A3(new_n392_), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n912_), .B1(new_n889_), .B2(new_n913_), .ZN(G1351gat));
  NOR3_X1   g713(.A1(new_n563_), .A2(new_n469_), .A3(new_n555_), .ZN(new_n915_));
  NAND3_X1  g714(.A1(new_n868_), .A2(new_n720_), .A3(new_n915_), .ZN(new_n916_));
  XNOR2_X1  g715(.A(new_n916_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g716(.A1(new_n868_), .A2(new_n283_), .A3(new_n915_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g718(.A1(new_n868_), .A2(new_n614_), .A3(new_n915_), .ZN(new_n920_));
  NOR2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  AND2_X1   g720(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n922_));
  NOR3_X1   g721(.A1(new_n920_), .A2(new_n921_), .A3(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n920_), .A2(new_n921_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(KEYINPUT127), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n920_), .A2(new_n926_), .A3(new_n921_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n923_), .B1(new_n925_), .B2(new_n927_), .ZN(G1354gat));
  AND4_X1   g727(.A1(G218gat), .A2(new_n868_), .A3(new_n602_), .A4(new_n915_), .ZN(new_n929_));
  INV_X1    g728(.A(G218gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n868_), .A2(new_n730_), .A3(new_n915_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n929_), .B1(new_n930_), .B2(new_n931_), .ZN(G1355gat));
endmodule


