//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:20 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n631_, new_n632_, new_n633_, new_n634_, new_n636_,
    new_n637_, new_n638_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n872_, new_n873_, new_n874_, new_n876_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_;
  INV_X1    g000(.A(KEYINPUT27), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT87), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n204_), .A2(G183gat), .A3(G190gat), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT80), .ZN(new_n206_));
  OR2_X1    g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G183gat), .ZN(new_n208_));
  INV_X1    g007(.A(G190gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT23), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n210_), .A2(new_n206_), .A3(new_n205_), .ZN(new_n211_));
  AND2_X1   g010(.A1(new_n207_), .A2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  XNOR2_X1  g012(.A(KEYINPUT25), .B(G183gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT24), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n216_), .B1(G169gat), .B2(G176gat), .ZN(new_n217_));
  INV_X1    g016(.A(G169gat), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n217_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n215_), .A2(KEYINPUT86), .A3(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n216_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n212_), .A2(new_n222_), .A3(new_n223_), .ZN(new_n224_));
  AOI22_X1  g023(.A1(new_n213_), .A2(new_n214_), .B1(new_n217_), .B2(new_n220_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n225_), .A2(KEYINPUT86), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n203_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n207_), .A2(new_n211_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(KEYINPUT86), .B2(new_n225_), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n225_), .A2(KEYINPUT86), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n229_), .A2(KEYINPUT87), .A3(new_n230_), .A4(new_n223_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n210_), .A2(new_n205_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n208_), .A2(new_n209_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT88), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT22), .B(G169gat), .Z(new_n238_));
  MUX2_X1   g037(.A(new_n218_), .B(new_n238_), .S(new_n219_), .Z(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n232_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT89), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G211gat), .B(G218gat), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n243_), .A2(KEYINPUT21), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(KEYINPUT21), .ZN(new_n245_));
  XOR2_X1   g044(.A(G197gat), .B(G204gat), .Z(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  OR2_X1    g046(.A1(new_n245_), .A2(new_n246_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  NAND3_X1  g048(.A1(new_n241_), .A2(new_n242_), .A3(new_n249_), .ZN(new_n250_));
  AOI22_X1  g049(.A1(new_n227_), .A2(new_n231_), .B1(new_n239_), .B2(new_n237_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n249_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT89), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT81), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n212_), .A2(new_n254_), .A3(new_n234_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n207_), .A2(new_n211_), .A3(new_n234_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT81), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n239_), .A3(new_n257_), .ZN(new_n258_));
  OR2_X1    g057(.A1(new_n213_), .A2(KEYINPUT79), .ZN(new_n259_));
  OR2_X1    g058(.A1(new_n214_), .A2(KEYINPUT78), .ZN(new_n260_));
  OAI21_X1  g059(.A(KEYINPUT78), .B1(new_n208_), .B2(KEYINPUT25), .ZN(new_n261_));
  OAI21_X1  g060(.A(KEYINPUT79), .B1(new_n209_), .B2(KEYINPUT26), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n259_), .A2(new_n260_), .A3(new_n261_), .A4(new_n262_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n263_), .A2(new_n233_), .A3(new_n221_), .A4(new_n223_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n258_), .A2(new_n264_), .A3(new_n252_), .ZN(new_n265_));
  AND2_X1   g064(.A1(new_n265_), .A2(KEYINPUT20), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n250_), .A2(new_n253_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n268_), .B(KEYINPUT85), .Z(new_n269_));
  XOR2_X1   g068(.A(new_n269_), .B(KEYINPUT19), .Z(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n267_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT18), .B(G64gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n273_), .B(G92gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G8gat), .B(G36gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n274_), .B(new_n275_), .Z(new_n276_));
  AOI21_X1  g075(.A(new_n249_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n232_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n258_), .A2(new_n264_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n279_), .A2(new_n249_), .ZN(new_n280_));
  NAND4_X1  g079(.A1(new_n278_), .A2(KEYINPUT20), .A3(new_n280_), .A4(new_n270_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n272_), .A2(new_n276_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n276_), .B1(new_n272_), .B2(new_n281_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n202_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n277_), .B1(new_n226_), .B2(new_n224_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n280_), .A2(new_n286_), .A3(KEYINPUT20), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(new_n271_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n288_), .B1(new_n267_), .B2(new_n271_), .ZN(new_n289_));
  INV_X1    g088(.A(new_n276_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(KEYINPUT27), .A3(new_n282_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n285_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT93), .ZN(new_n295_));
  INV_X1    g094(.A(G120gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(G127gat), .B(G134gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(G113gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(new_n297_), .A2(G113gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n296_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n300_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(G120gat), .A3(new_n298_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  AND2_X1   g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305_));
  NOR2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n308_));
  NOR2_X1   g107(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n308_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n312_));
  NOR2_X1   g111(.A1(G141gat), .A2(G148gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n311_), .A2(new_n312_), .A3(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n310_), .A2(new_n308_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n307_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n313_), .B1(new_n307_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n305_), .A2(KEYINPUT1), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n320_), .A2(new_n310_), .A3(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n304_), .A2(new_n323_), .ZN(new_n324_));
  OR2_X1    g123(.A1(new_n324_), .A2(KEYINPUT4), .ZN(new_n325_));
  NAND2_X1  g124(.A1(G225gat), .A2(G233gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT90), .ZN(new_n327_));
  NAND4_X1  g126(.A1(new_n301_), .A2(new_n303_), .A3(new_n318_), .A4(new_n322_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n324_), .A2(KEYINPUT4), .A3(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n325_), .A2(new_n327_), .A3(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n324_), .A2(new_n326_), .A3(new_n328_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(KEYINPUT0), .B(G57gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n332_), .B(G85gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(G1gat), .B(G29gat), .Z(new_n334_));
  XOR2_X1   g133(.A(new_n333_), .B(new_n334_), .Z(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n330_), .A2(new_n331_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n336_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n295_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n339_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n341_), .A2(KEYINPUT93), .A3(new_n337_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n340_), .A2(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n318_), .B2(new_n322_), .ZN(new_n345_));
  OR3_X1    g144(.A1(new_n252_), .A2(new_n345_), .A3(G22gat), .ZN(new_n346_));
  OAI21_X1  g145(.A(G22gat), .B1(new_n252_), .B2(new_n345_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n318_), .A2(new_n322_), .A3(new_n344_), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n349_), .B(KEYINPUT28), .Z(new_n350_));
  NOR2_X1   g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n348_), .A2(new_n350_), .ZN(new_n353_));
  INV_X1    g152(.A(G228gat), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT84), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n355_), .A2(G233gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(G233gat), .ZN(new_n357_));
  AOI21_X1  g156(.A(new_n354_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(G50gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  XOR2_X1   g159(.A(G78gat), .B(G106gat), .Z(new_n361_));
  XNOR2_X1  g160(.A(new_n360_), .B(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n352_), .A2(new_n353_), .A3(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n362_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n279_), .A2(new_n304_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n279_), .A2(new_n304_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n366_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n369_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n366_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n371_), .A2(new_n367_), .A3(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G71gat), .B(G99gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT31), .ZN(new_n375_));
  XOR2_X1   g174(.A(G15gat), .B(G43gat), .Z(new_n376_));
  XNOR2_X1  g175(.A(new_n375_), .B(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G227gat), .A2(G233gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n370_), .A2(new_n373_), .A3(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n379_), .B1(new_n370_), .B2(new_n373_), .ZN(new_n382_));
  OAI22_X1  g181(.A1(new_n364_), .A2(new_n365_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n382_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n362_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n353_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n385_), .B1(new_n386_), .B2(new_n351_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n384_), .A2(new_n363_), .A3(new_n387_), .A4(new_n380_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n343_), .B1(new_n383_), .B2(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n384_), .A2(new_n380_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n272_), .A2(new_n281_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(new_n290_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n324_), .A2(new_n328_), .A3(new_n327_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n335_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT91), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT91), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n393_), .A2(new_n396_), .A3(new_n335_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n325_), .A2(new_n326_), .A3(new_n329_), .ZN(new_n399_));
  AOI21_X1  g198(.A(KEYINPUT92), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  AND4_X1   g199(.A1(KEYINPUT92), .A2(new_n395_), .A3(new_n399_), .A4(new_n397_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n337_), .B(KEYINPUT33), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n392_), .A2(new_n402_), .A3(new_n282_), .A4(new_n403_), .ZN(new_n404_));
  AND2_X1   g203(.A1(new_n276_), .A2(KEYINPUT32), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n289_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n341_), .A2(new_n337_), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n406_), .B(new_n407_), .C1(new_n405_), .C2(new_n391_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n390_), .B1(new_n404_), .B2(new_n408_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n364_), .A2(new_n365_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI22_X1  g210(.A1(new_n294_), .A2(new_n389_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT67), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n413_), .A2(G71gat), .ZN(new_n414_));
  INV_X1    g213(.A(G71gat), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n415_), .A2(KEYINPUT67), .ZN(new_n416_));
  OAI21_X1  g215(.A(G78gat), .B1(new_n414_), .B2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(G57gat), .A2(G64gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT11), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G57gat), .A2(G64gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n419_), .A2(new_n420_), .A3(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n421_), .ZN(new_n423_));
  OAI21_X1  g222(.A(KEYINPUT11), .B1(new_n423_), .B2(new_n418_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n415_), .A2(KEYINPUT67), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n413_), .A2(G71gat), .ZN(new_n426_));
  INV_X1    g225(.A(G78gat), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n417_), .A2(new_n422_), .A3(new_n424_), .A4(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n420_), .B1(new_n419_), .B2(new_n421_), .ZN(new_n430_));
  AND3_X1   g229(.A1(new_n425_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n427_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n432_));
  OAI21_X1  g231(.A(new_n430_), .B1(new_n431_), .B2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n429_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G85gat), .ZN(new_n435_));
  INV_X1    g234(.A(G92gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT65), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT9), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G85gat), .A2(G92gat), .ZN(new_n440_));
  NAND4_X1  g239(.A1(new_n437_), .A2(new_n438_), .A3(new_n439_), .A4(new_n440_), .ZN(new_n441_));
  AND2_X1   g240(.A1(G85gat), .A2(G92gat), .ZN(new_n442_));
  NOR2_X1   g241(.A1(G85gat), .A2(G92gat), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n442_), .A2(new_n443_), .A3(KEYINPUT65), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n443_), .A2(KEYINPUT9), .ZN(new_n445_));
  OAI211_X1 g244(.A(KEYINPUT66), .B(new_n441_), .C1(new_n444_), .C2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(G99gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT10), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT10), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(G99gat), .ZN(new_n450_));
  AOI21_X1  g249(.A(G106gat), .B1(new_n448_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G99gat), .A2(G106gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT6), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n440_), .A2(new_n439_), .A3(KEYINPUT66), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n451_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n446_), .A2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT8), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT7), .ZN(new_n461_));
  INV_X1    g260(.A(G106gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n461_), .A2(new_n447_), .A3(new_n462_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n463_), .A2(new_n454_), .A3(new_n455_), .A4(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n442_), .A2(new_n443_), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n460_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  AND3_X1   g266(.A1(new_n465_), .A2(new_n460_), .A3(new_n466_), .ZN(new_n468_));
  OAI211_X1 g267(.A(new_n434_), .B(new_n459_), .C1(new_n467_), .C2(new_n468_), .ZN(new_n469_));
  XOR2_X1   g268(.A(KEYINPUT69), .B(KEYINPUT12), .Z(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n465_), .A2(new_n466_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT8), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n465_), .A2(new_n460_), .A3(new_n466_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(new_n459_), .ZN(new_n476_));
  INV_X1    g275(.A(new_n434_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT68), .B1(new_n468_), .B2(new_n467_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT68), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n473_), .A2(new_n480_), .A3(new_n474_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n479_), .A2(new_n481_), .A3(new_n459_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n429_), .A2(new_n433_), .A3(KEYINPUT12), .ZN(new_n483_));
  AOI22_X1  g282(.A1(new_n471_), .A2(new_n478_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G230gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT64), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n484_), .A2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n478_), .A2(new_n469_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n486_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G120gat), .B(G148gat), .ZN(new_n492_));
  INV_X1    g291(.A(G204gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT5), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(new_n219_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n491_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT70), .ZN(new_n499_));
  INV_X1    g298(.A(new_n491_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n499_), .B1(new_n500_), .B2(new_n496_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(new_n491_), .A2(KEYINPUT70), .A3(new_n497_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n498_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(KEYINPUT13), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT13), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n505_), .B(new_n498_), .C1(new_n501_), .C2(new_n502_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT15), .ZN(new_n508_));
  INV_X1    g307(.A(G29gat), .ZN(new_n509_));
  INV_X1    g308(.A(G36gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G29gat), .A2(G36gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(G43gat), .ZN(new_n514_));
  INV_X1    g313(.A(G43gat), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n511_), .A2(new_n515_), .A3(new_n512_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(G50gat), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(G50gat), .B1(new_n514_), .B2(new_n516_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n508_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n514_), .A2(new_n516_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n359_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n522_), .A2(KEYINPUT15), .A3(new_n517_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n520_), .A2(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G15gat), .B(G22gat), .ZN(new_n525_));
  INV_X1    g324(.A(G1gat), .ZN(new_n526_));
  INV_X1    g325(.A(G8gat), .ZN(new_n527_));
  OAI21_X1  g326(.A(KEYINPUT14), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G1gat), .B(G8gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n524_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n531_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n518_), .A2(new_n519_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G229gat), .A2(G233gat), .ZN(new_n536_));
  XOR2_X1   g335(.A(new_n536_), .B(KEYINPUT76), .Z(new_n537_));
  NAND3_X1  g336(.A1(new_n532_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n538_), .A2(KEYINPUT77), .ZN(new_n539_));
  OR3_X1    g338(.A1(new_n533_), .A2(new_n534_), .A3(KEYINPUT75), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n531_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n535_), .A2(KEYINPUT75), .A3(new_n541_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n540_), .A2(new_n542_), .A3(G229gat), .A4(G233gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n538_), .A2(KEYINPUT77), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n539_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G113gat), .B(G141gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(new_n218_), .ZN(new_n547_));
  INV_X1    g346(.A(G197gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n545_), .A2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n549_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n539_), .A2(new_n543_), .A3(new_n544_), .A4(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n507_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n412_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT34), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(KEYINPUT71), .B(KEYINPUT35), .Z(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n482_), .A2(new_n524_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT72), .ZN(new_n566_));
  AOI22_X1  g365(.A1(new_n473_), .A2(new_n474_), .B1(new_n446_), .B2(new_n458_), .ZN(new_n567_));
  AOI22_X1  g366(.A1(new_n567_), .A2(new_n534_), .B1(new_n560_), .B2(new_n562_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n565_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n566_), .B1(new_n565_), .B2(new_n568_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n564_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n565_), .A2(new_n568_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT72), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n565_), .A2(new_n566_), .A3(new_n568_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n563_), .A3(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n571_), .A2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G190gat), .B(G218gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(G134gat), .ZN(new_n578_));
  INV_X1    g377(.A(G162gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT36), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n580_), .A2(new_n581_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n576_), .A2(new_n583_), .A3(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT74), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT37), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n576_), .A2(KEYINPUT74), .A3(new_n583_), .A4(new_n584_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n584_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n571_), .A2(new_n575_), .A3(new_n590_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n587_), .A2(new_n588_), .A3(new_n589_), .A4(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT73), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n571_), .A2(new_n575_), .A3(KEYINPUT73), .A4(new_n590_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n594_), .A2(new_n585_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT37), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n592_), .A2(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n434_), .B(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(new_n533_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT16), .B(G183gat), .ZN(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(G211gat), .ZN(new_n603_));
  XOR2_X1   g402(.A(G127gat), .B(G155gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT17), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n601_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n605_), .B(KEYINPUT17), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n608_), .B1(new_n601_), .B2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n598_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n557_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n616_), .A2(new_n526_), .A3(new_n343_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT38), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n587_), .A2(new_n589_), .A3(new_n591_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(new_n611_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n557_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n343_), .ZN(new_n623_));
  OAI21_X1  g422(.A(G1gat), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n618_), .A2(new_n624_), .ZN(G1324gat));
  OAI21_X1  g424(.A(G8gat), .B1(new_n622_), .B2(new_n294_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT39), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n616_), .A2(new_n527_), .A3(new_n293_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n629_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g429(.A(new_n390_), .ZN(new_n631_));
  OAI21_X1  g430(.A(G15gat), .B1(new_n622_), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT41), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n615_), .A2(G15gat), .A3(new_n631_), .ZN(new_n634_));
  OR2_X1    g433(.A1(new_n633_), .A2(new_n634_), .ZN(G1326gat));
  OAI21_X1  g434(.A(G22gat), .B1(new_n622_), .B2(new_n411_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT94), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT42), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n411_), .A2(G22gat), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT95), .Z(new_n641_));
  NAND2_X1  g440(.A1(new_n616_), .A2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n639_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT96), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT96), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n639_), .A2(new_n645_), .A3(new_n642_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(G1327gat));
  NOR2_X1   g446(.A1(new_n619_), .A2(new_n612_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n557_), .A2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT97), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n649_), .B(new_n650_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(new_n509_), .A3(new_n343_), .ZN(new_n652_));
  OAI21_X1  g451(.A(KEYINPUT43), .B1(new_n412_), .B2(new_n598_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n404_), .A2(new_n408_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n654_), .A2(new_n411_), .A3(new_n631_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n389_), .A2(new_n285_), .A3(new_n292_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n592_), .A2(new_n597_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n653_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n611_), .A3(new_n555_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT44), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n661_), .A2(KEYINPUT44), .A3(new_n611_), .A4(new_n555_), .ZN(new_n665_));
  AND2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n666_), .A2(new_n343_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n652_), .B1(new_n667_), .B2(new_n509_), .ZN(G1328gat));
  NAND3_X1  g467(.A1(new_n651_), .A2(new_n510_), .A3(new_n293_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT45), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n664_), .A2(new_n293_), .A3(new_n665_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT98), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND4_X1  g472(.A1(new_n664_), .A2(KEYINPUT98), .A3(new_n293_), .A4(new_n665_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(G36gat), .A3(new_n674_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n670_), .A2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT46), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(KEYINPUT99), .A3(new_n677_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n677_), .A2(KEYINPUT99), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n670_), .A2(new_n675_), .A3(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n678_), .A2(new_n680_), .ZN(G1329gat));
  NAND3_X1  g480(.A1(new_n666_), .A2(G43gat), .A3(new_n390_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n651_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n515_), .B1(new_n683_), .B2(new_n631_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g485(.A1(new_n651_), .A2(new_n359_), .A3(new_n410_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT100), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n666_), .A2(new_n410_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n688_), .B1(new_n689_), .B2(G50gat), .ZN(new_n690_));
  AOI211_X1 g489(.A(KEYINPUT100), .B(new_n359_), .C1(new_n666_), .C2(new_n410_), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n687_), .B1(new_n690_), .B2(new_n691_), .ZN(G1331gat));
  NAND2_X1  g491(.A1(new_n657_), .A2(new_n554_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(new_n507_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n614_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G57gat), .B1(new_n698_), .B2(new_n343_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n657_), .A2(new_n621_), .A3(new_n554_), .A4(new_n507_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n700_), .A2(new_n623_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n699_), .B1(G57gat), .B2(new_n701_), .ZN(G1332gat));
  OAI21_X1  g501(.A(G64gat), .B1(new_n700_), .B2(new_n294_), .ZN(new_n703_));
  XOR2_X1   g502(.A(new_n703_), .B(KEYINPUT102), .Z(new_n704_));
  XOR2_X1   g503(.A(new_n704_), .B(KEYINPUT48), .Z(new_n705_));
  NOR3_X1   g504(.A1(new_n697_), .A2(G64gat), .A3(new_n294_), .ZN(new_n706_));
  OR2_X1    g505(.A1(new_n705_), .A2(new_n706_), .ZN(G1333gat));
  OAI21_X1  g506(.A(G71gat), .B1(new_n700_), .B2(new_n631_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT49), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n390_), .A2(new_n415_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n697_), .B2(new_n710_), .ZN(G1334gat));
  OAI21_X1  g510(.A(G78gat), .B1(new_n700_), .B2(new_n411_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT50), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n410_), .A2(new_n427_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n713_), .B1(new_n697_), .B2(new_n714_), .ZN(G1335gat));
  NAND3_X1  g514(.A1(new_n695_), .A2(new_n507_), .A3(new_n648_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(G85gat), .B1(new_n717_), .B2(new_n343_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n507_), .A2(new_n611_), .A3(new_n554_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NAND4_X1  g520(.A1(new_n507_), .A2(KEYINPUT103), .A3(new_n611_), .A4(new_n554_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n661_), .A2(new_n723_), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n724_), .A2(KEYINPUT104), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(KEYINPUT104), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n623_), .A2(new_n435_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n718_), .B1(new_n727_), .B2(new_n728_), .ZN(G1336gat));
  AOI21_X1  g528(.A(G92gat), .B1(new_n717_), .B2(new_n293_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n294_), .A2(new_n436_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n727_), .B2(new_n731_), .ZN(G1337gat));
  NAND3_X1  g531(.A1(new_n725_), .A2(new_n390_), .A3(new_n726_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(G99gat), .ZN(new_n734_));
  NAND2_X1  g533(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n448_), .A2(new_n450_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n717_), .A2(new_n736_), .A3(new_n390_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n734_), .A2(new_n735_), .A3(new_n737_), .ZN(new_n738_));
  OR2_X1    g537(.A1(KEYINPUT105), .A2(KEYINPUT51), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n738_), .B(new_n739_), .ZN(G1338gat));
  AOI21_X1  g539(.A(new_n658_), .B1(new_n657_), .B2(new_n659_), .ZN(new_n741_));
  AOI211_X1 g540(.A(KEYINPUT43), .B(new_n598_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n410_), .B(new_n723_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n661_), .A2(KEYINPUT106), .A3(new_n410_), .A4(new_n723_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n745_), .A2(new_n746_), .A3(G106gat), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(KEYINPUT52), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT52), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n745_), .A2(new_n746_), .A3(new_n749_), .A4(G106gat), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n410_), .A2(new_n462_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n716_), .A2(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n751_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT107), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT107), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n751_), .A2(new_n757_), .A3(new_n754_), .ZN(new_n758_));
  AOI21_X1  g557(.A(KEYINPUT53), .B1(new_n756_), .B2(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n757_), .B1(new_n751_), .B2(new_n754_), .ZN(new_n760_));
  AOI211_X1 g559(.A(KEYINPUT107), .B(new_n753_), .C1(new_n748_), .C2(new_n750_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT53), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n760_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n759_), .A2(new_n763_), .ZN(G1339gat));
  INV_X1    g563(.A(KEYINPUT109), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n434_), .B1(new_n475_), .B2(new_n459_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n767_));
  AND2_X1   g566(.A1(new_n482_), .A2(new_n483_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n489_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n765_), .B1(new_n769_), .B2(KEYINPUT55), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n765_), .B(KEYINPUT55), .C1(new_n484_), .C2(new_n486_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n487_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n484_), .A2(new_n486_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  OAI21_X1  g574(.A(KEYINPUT109), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n487_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n776_), .A2(new_n777_), .A3(new_n771_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n773_), .A2(new_n497_), .A3(new_n778_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT56), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n773_), .A2(new_n778_), .A3(KEYINPUT56), .A4(new_n497_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n540_), .A2(new_n542_), .A3(new_n537_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n532_), .A2(new_n535_), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n784_), .B(new_n549_), .C1(new_n785_), .C2(new_n537_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n552_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n788_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n789_));
  INV_X1    g588(.A(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT58), .B1(new_n783_), .B2(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(KEYINPUT112), .B1(new_n791_), .B2(new_n598_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT112), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n789_), .B1(new_n781_), .B2(new_n782_), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n659_), .B(new_n793_), .C1(KEYINPUT58), .C2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(KEYINPUT58), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(KEYINPUT113), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT113), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n794_), .A2(new_n798_), .A3(KEYINPUT58), .ZN(new_n799_));
  NAND4_X1  g598(.A1(new_n792_), .A2(new_n795_), .A3(new_n797_), .A4(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n503_), .A2(new_n788_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(KEYINPUT110), .B(KEYINPUT56), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n779_), .A2(KEYINPUT111), .A3(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(KEYINPUT111), .B1(new_n779_), .B2(new_n802_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n782_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n803_), .A2(new_n804_), .A3(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n501_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n502_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n553_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n801_), .B1(new_n806_), .B2(new_n810_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT57), .A3(new_n619_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT57), .ZN(new_n813_));
  INV_X1    g612(.A(new_n801_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n779_), .A2(new_n802_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n779_), .A2(KEYINPUT111), .A3(new_n802_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n782_), .A3(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n810_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n814_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n813_), .B1(new_n821_), .B2(new_n620_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n800_), .A2(new_n812_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n611_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT108), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n504_), .A2(new_n506_), .ZN(new_n828_));
  NAND4_X1  g627(.A1(new_n598_), .A2(new_n612_), .A3(new_n828_), .A4(new_n554_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n827_), .B1(new_n829_), .B2(KEYINPUT54), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n611_), .B(new_n553_), .C1(new_n592_), .C2(new_n597_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n831_), .A2(KEYINPUT108), .A3(new_n832_), .A4(new_n828_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n829_), .A2(KEYINPUT54), .ZN(new_n834_));
  AND3_X1   g633(.A1(new_n830_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n823_), .A2(KEYINPUT115), .A3(new_n611_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n826_), .A2(new_n836_), .A3(new_n837_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n293_), .A2(new_n623_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n840_), .A2(new_n383_), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT59), .B1(new_n841_), .B2(KEYINPUT114), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n842_), .B1(KEYINPUT114), .B2(new_n841_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n838_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n824_), .A2(new_n836_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n841_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT59), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n845_), .A2(new_n848_), .ZN(new_n849_));
  AND3_X1   g648(.A1(new_n849_), .A2(G113gat), .A3(new_n553_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n847_), .ZN(new_n851_));
  AOI21_X1  g650(.A(G113gat), .B1(new_n851_), .B2(new_n553_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n850_), .A2(new_n852_), .ZN(G1340gat));
  NAND3_X1  g652(.A1(new_n845_), .A2(new_n507_), .A3(new_n848_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT116), .B(G120gat), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n845_), .A2(new_n848_), .A3(KEYINPUT117), .A4(new_n507_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n857_), .A3(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT60), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n828_), .B2(new_n857_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n851_), .B(new_n861_), .C1(new_n860_), .C2(new_n857_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n859_), .A2(new_n862_), .ZN(G1341gat));
  AOI21_X1  g662(.A(G127gat), .B1(new_n851_), .B2(new_n612_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n612_), .A2(G127gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n864_), .B1(new_n849_), .B2(new_n865_), .ZN(G1342gat));
  NAND3_X1  g665(.A1(new_n849_), .A2(G134gat), .A3(new_n659_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  AOI21_X1  g667(.A(G134gat), .B1(new_n851_), .B2(new_n620_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(KEYINPUT118), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n868_), .A2(new_n870_), .ZN(G1343gat));
  AOI21_X1  g670(.A(new_n835_), .B1(new_n823_), .B2(new_n611_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n872_), .A2(new_n388_), .A3(new_n840_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n553_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n873_), .A2(new_n507_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n612_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT61), .B(G155gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1346gat));
  AOI21_X1  g679(.A(G162gat), .B1(new_n873_), .B2(new_n620_), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n882_));
  OR2_X1    g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n882_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n598_), .A2(new_n579_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n883_), .A2(new_n884_), .B1(new_n873_), .B2(new_n885_), .ZN(G1347gat));
  NOR2_X1   g685(.A1(new_n294_), .A2(new_n343_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(new_n390_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT120), .ZN(new_n889_));
  NAND4_X1  g688(.A1(new_n838_), .A2(new_n553_), .A3(new_n411_), .A4(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(G169gat), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n890_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n893_), .B(new_n894_), .C1(new_n238_), .C2(new_n890_), .ZN(G1348gat));
  NOR2_X1   g694(.A1(new_n872_), .A2(new_n410_), .ZN(new_n896_));
  AND4_X1   g695(.A1(G176gat), .A2(new_n896_), .A3(new_n507_), .A4(new_n889_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n838_), .A2(new_n411_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n898_), .A2(new_n507_), .A3(new_n889_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n897_), .B1(new_n899_), .B2(new_n219_), .ZN(G1349gat));
  NOR2_X1   g699(.A1(new_n611_), .A2(new_n214_), .ZN(new_n901_));
  NAND4_X1  g700(.A1(new_n838_), .A2(new_n411_), .A3(new_n889_), .A4(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n902_), .A2(new_n903_), .ZN(new_n905_));
  NAND3_X1  g704(.A1(new_n896_), .A2(new_n612_), .A3(new_n889_), .ZN(new_n906_));
  AOI211_X1 g705(.A(new_n904_), .B(new_n905_), .C1(new_n208_), .C2(new_n906_), .ZN(G1350gat));
  NAND4_X1  g706(.A1(new_n838_), .A2(new_n411_), .A3(new_n659_), .A4(new_n889_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT122), .ZN(new_n909_));
  AND3_X1   g708(.A1(new_n908_), .A2(new_n909_), .A3(G190gat), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n909_), .B1(new_n908_), .B2(G190gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n898_), .A2(new_n889_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n620_), .A2(new_n213_), .ZN(new_n913_));
  OAI22_X1  g712(.A1(new_n910_), .A2(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(G1351gat));
  AOI21_X1  g713(.A(new_n388_), .B1(new_n824_), .B2(new_n836_), .ZN(new_n915_));
  AOI21_X1  g714(.A(KEYINPUT123), .B1(new_n915_), .B2(new_n887_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT123), .ZN(new_n917_));
  INV_X1    g716(.A(new_n887_), .ZN(new_n918_));
  NOR4_X1   g717(.A1(new_n872_), .A2(new_n917_), .A3(new_n388_), .A4(new_n918_), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n916_), .A2(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n553_), .ZN(new_n921_));
  XNOR2_X1  g720(.A(new_n921_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g721(.A1(new_n920_), .A2(new_n507_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n493_), .A2(KEYINPUT124), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  AOI22_X1  g724(.A1(new_n920_), .A2(new_n507_), .B1(KEYINPUT124), .B2(new_n493_), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(new_n924_), .ZN(G1353gat));
  INV_X1    g726(.A(KEYINPUT63), .ZN(new_n928_));
  INV_X1    g727(.A(G211gat), .ZN(new_n929_));
  OAI21_X1  g728(.A(new_n612_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT125), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n920_), .A2(new_n931_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n928_), .A2(new_n929_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1354gat));
  OAI21_X1  g733(.A(new_n620_), .B1(new_n916_), .B2(new_n919_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n935_), .A2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(G218gat), .ZN(new_n938_));
  OAI211_X1 g737(.A(KEYINPUT126), .B(new_n620_), .C1(new_n916_), .C2(new_n919_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n937_), .A2(new_n938_), .A3(new_n939_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n659_), .A2(G218gat), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(KEYINPUT127), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n920_), .A2(new_n942_), .ZN(new_n943_));
  AND2_X1   g742(.A1(new_n940_), .A2(new_n943_), .ZN(G1355gat));
endmodule


