//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n591_, new_n592_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n599_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_;
  INV_X1    g000(.A(KEYINPUT20), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G183gat), .A2(G190gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT23), .ZN(new_n204_));
  OAI21_X1  g003(.A(new_n204_), .B1(G183gat), .B2(G190gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G169gat), .A2(G176gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(G176gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT22), .B(G169gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT91), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n207_), .B1(new_n208_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT92), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n206_), .A2(KEYINPUT24), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215_));
  MUX2_X1   g014(.A(new_n214_), .B(KEYINPUT24), .S(new_n215_), .Z(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT26), .B(G190gat), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  XOR2_X1   g017(.A(KEYINPUT25), .B(G183gat), .Z(new_n219_));
  OAI211_X1 g018(.A(new_n216_), .B(new_n204_), .C1(new_n218_), .C2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n213_), .A2(new_n220_), .ZN(new_n221_));
  XOR2_X1   g020(.A(G211gat), .B(G218gat), .Z(new_n222_));
  INV_X1    g021(.A(KEYINPUT21), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G197gat), .B(G204gat), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n222_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n224_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT21), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n226_), .A2(new_n222_), .A3(KEYINPUT21), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n202_), .B1(new_n221_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT22), .ZN(new_n232_));
  INV_X1    g031(.A(G169gat), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n233_), .A2(KEYINPUT80), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT80), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(G169gat), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n232_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n237_), .B(KEYINPUT81), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n208_), .B1(new_n233_), .B2(KEYINPUT22), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n206_), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT79), .B(G183gat), .Z(new_n241_));
  INV_X1    g040(.A(G190gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  AOI22_X1  g042(.A1(new_n240_), .A2(KEYINPUT82), .B1(new_n204_), .B2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n244_), .B1(KEYINPUT82), .B2(new_n240_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n230_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT25), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n241_), .A2(new_n247_), .ZN(new_n248_));
  NOR2_X1   g047(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n217_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(new_n204_), .A3(new_n216_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n245_), .A2(new_n246_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n231_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(G226gat), .A2(G233gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(KEYINPUT89), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n257_), .B(KEYINPUT90), .Z(new_n258_));
  NAND2_X1  g057(.A1(new_n253_), .A2(new_n258_), .ZN(new_n259_));
  XOR2_X1   g058(.A(G8gat), .B(G36gat), .Z(new_n260_));
  XNOR2_X1  g059(.A(G64gat), .B(G92gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n257_), .A2(new_n202_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n265_), .B1(new_n221_), .B2(new_n230_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n246_), .B1(new_n245_), .B2(new_n251_), .ZN(new_n267_));
  OR2_X1    g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n259_), .A2(new_n264_), .A3(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n264_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n258_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n271_), .B1(new_n231_), .B2(new_n252_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n266_), .A2(new_n267_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n270_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT27), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n246_), .A2(new_n220_), .ZN(new_n278_));
  OAI21_X1  g077(.A(KEYINPUT20), .B1(new_n278_), .B2(new_n211_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n257_), .B1(new_n267_), .B2(new_n279_), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n280_), .B1(new_n253_), .B2(new_n258_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n270_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(KEYINPUT27), .A3(new_n269_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n277_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G155gat), .A2(G162gat), .ZN(new_n286_));
  NOR2_X1   g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NOR2_X1   g087(.A1(G141gat), .A2(G148gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n289_), .B(KEYINPUT3), .Z(new_n290_));
  NAND2_X1  g089(.A1(G141gat), .A2(G148gat), .ZN(new_n291_));
  XOR2_X1   g090(.A(new_n291_), .B(KEYINPUT2), .Z(new_n292_));
  OAI211_X1 g091(.A(new_n286_), .B(new_n288_), .C1(new_n290_), .C2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n287_), .B1(KEYINPUT1), .B2(new_n286_), .ZN(new_n294_));
  OAI21_X1  g093(.A(new_n294_), .B1(KEYINPUT1), .B2(new_n286_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n289_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(new_n296_), .A3(new_n291_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n293_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT29), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G22gat), .B(G50gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n230_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n305_));
  INV_X1    g104(.A(G233gat), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n306_), .A2(KEYINPUT86), .ZN(new_n307_));
  NOR2_X1   g106(.A1(new_n306_), .A2(KEYINPUT86), .ZN(new_n308_));
  OAI21_X1  g107(.A(G228gat), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n305_), .A2(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(new_n230_), .B(new_n309_), .C1(new_n299_), .C2(new_n300_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G78gat), .B(G106gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(KEYINPUT85), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT87), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n312_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n314_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n315_), .A2(new_n316_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n319_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT85), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n322_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT87), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(KEYINPUT84), .B(KEYINPUT28), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  AND3_X1   g125(.A1(new_n320_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n326_), .B1(new_n320_), .B2(new_n324_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n304_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n320_), .A2(new_n324_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n330_), .A2(new_n325_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n320_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n331_), .A2(new_n303_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  XOR2_X1   g133(.A(G1gat), .B(G29gat), .Z(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G57gat), .B(G85gat), .ZN(new_n338_));
  XOR2_X1   g137(.A(new_n337_), .B(new_n338_), .Z(new_n339_));
  XNOR2_X1  g138(.A(G127gat), .B(G134gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G113gat), .B(G120gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n298_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  OR3_X1    g146(.A1(new_n299_), .A2(KEYINPUT95), .A3(new_n342_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n299_), .A2(new_n342_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(new_n348_), .A2(KEYINPUT4), .A3(new_n349_), .ZN(new_n350_));
  OR4_X1    g149(.A1(KEYINPUT95), .A2(new_n299_), .A3(KEYINPUT4), .A4(new_n342_), .ZN(new_n351_));
  AND2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  OAI211_X1 g151(.A(new_n339_), .B(new_n347_), .C1(new_n352_), .C2(new_n344_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n339_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n344_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n354_), .B1(new_n355_), .B2(new_n346_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n353_), .A2(new_n356_), .A3(KEYINPUT97), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT97), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n358_), .B(new_n354_), .C1(new_n355_), .C2(new_n346_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n245_), .A2(new_n251_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G71gat), .B(G99gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n362_), .B(G43gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n361_), .B(new_n363_), .ZN(new_n364_));
  XOR2_X1   g163(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n365_));
  XNOR2_X1  g164(.A(new_n364_), .B(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G227gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(G15gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT30), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(new_n342_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n366_), .B(new_n370_), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n285_), .A2(new_n334_), .A3(new_n360_), .A4(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT94), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n275_), .A2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n269_), .A2(KEYINPUT94), .A3(new_n274_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT33), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n356_), .A2(new_n376_), .ZN(new_n377_));
  OAI211_X1 g176(.A(KEYINPUT33), .B(new_n354_), .C1(new_n355_), .C2(new_n346_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n352_), .A2(new_n344_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n354_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n377_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n374_), .A2(new_n375_), .A3(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n357_), .A2(new_n359_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT98), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n264_), .A2(KEYINPUT32), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n259_), .A2(new_n268_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n281_), .A2(KEYINPUT32), .A3(new_n264_), .ZN(new_n388_));
  NAND4_X1  g187(.A1(new_n384_), .A2(new_n385_), .A3(new_n387_), .A4(new_n388_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n388_), .A2(new_n387_), .A3(new_n359_), .A4(new_n357_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(KEYINPUT98), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n383_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n329_), .A2(new_n333_), .A3(new_n360_), .ZN(new_n393_));
  AOI22_X1  g192(.A1(new_n392_), .A2(new_n334_), .B1(new_n393_), .B2(new_n285_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n372_), .B1(new_n394_), .B2(new_n371_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(G229gat), .A2(G233gat), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G1gat), .B(G8gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT75), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G15gat), .B(G22gat), .ZN(new_n401_));
  INV_X1    g200(.A(G1gat), .ZN(new_n402_));
  INV_X1    g201(.A(G8gat), .ZN(new_n403_));
  OAI21_X1  g202(.A(KEYINPUT14), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n400_), .A2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n398_), .B(KEYINPUT75), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n405_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G29gat), .B(G36gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G43gat), .B(G50gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n410_), .A2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT77), .ZN(new_n415_));
  AND3_X1   g214(.A1(new_n410_), .A2(new_n415_), .A3(new_n413_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n415_), .B1(new_n410_), .B2(new_n413_), .ZN(new_n417_));
  OAI211_X1 g216(.A(new_n397_), .B(new_n414_), .C1(new_n416_), .C2(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT78), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n408_), .A2(new_n405_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n400_), .A2(new_n406_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n413_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT77), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n410_), .A2(new_n415_), .A3(new_n413_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n410_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n413_), .B(KEYINPUT15), .ZN(new_n426_));
  AOI22_X1  g225(.A1(new_n423_), .A2(new_n424_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n418_), .B(new_n419_), .C1(new_n427_), .C2(new_n397_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G113gat), .B(G141gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G169gat), .B(G197gat), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n429_), .B(new_n430_), .Z(new_n431_));
  XNOR2_X1  g230(.A(new_n428_), .B(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n395_), .A2(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT68), .ZN(new_n434_));
  AND2_X1   g233(.A1(G85gat), .A2(G92gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(G85gat), .A2(G92gat), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G99gat), .A2(G106gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT6), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT6), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(G99gat), .A3(G106gat), .ZN(new_n441_));
  AND2_X1   g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT7), .ZN(new_n443_));
  INV_X1    g242(.A(G99gat), .ZN(new_n444_));
  INV_X1    g243(.A(G106gat), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n437_), .B1(new_n442_), .B2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(KEYINPUT8), .B1(new_n437_), .B2(KEYINPUT65), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OAI221_X1 g250(.A(new_n437_), .B1(KEYINPUT65), .B2(KEYINPUT8), .C1(new_n442_), .C2(new_n448_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(KEYINPUT9), .A2(G92gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT9), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n455_), .A2(KEYINPUT64), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n455_), .A2(KEYINPUT64), .ZN(new_n457_));
  OAI221_X1 g256(.A(new_n454_), .B1(new_n435_), .B2(new_n436_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n459_));
  NOR2_X1   g258(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n461_), .A2(new_n445_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n463_), .B1(new_n437_), .B2(new_n453_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n458_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n451_), .A2(new_n452_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT66), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n451_), .A2(new_n452_), .A3(new_n465_), .A4(KEYINPUT66), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G57gat), .B(G64gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT11), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT67), .B(G71gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(G78gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(G78gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n473_), .B(new_n476_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n471_), .A2(KEYINPUT11), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n475_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n470_), .A2(new_n480_), .ZN(new_n481_));
  AND2_X1   g280(.A1(new_n475_), .A2(new_n479_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n468_), .A2(new_n482_), .A3(new_n469_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G230gat), .A2(G233gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n434_), .B1(new_n484_), .B2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT12), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n481_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n480_), .A2(new_n466_), .A3(KEYINPUT12), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n483_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n491_), .A3(new_n485_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n487_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n483_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n482_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n434_), .B(new_n486_), .C1(new_n494_), .C2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  XOR2_X1   g296(.A(G120gat), .B(G148gat), .Z(new_n498_));
  XNOR2_X1  g297(.A(G176gat), .B(G204gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n498_), .B(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n501_));
  XOR2_X1   g300(.A(new_n500_), .B(new_n501_), .Z(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n497_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n496_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n505_), .B1(new_n487_), .B2(new_n492_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n506_), .A2(new_n502_), .ZN(new_n507_));
  AND2_X1   g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT70), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT13), .ZN(new_n510_));
  OAI21_X1  g309(.A(new_n508_), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n512_));
  OAI21_X1  g311(.A(new_n511_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n513_), .B(KEYINPUT71), .Z(new_n514_));
  INV_X1    g313(.A(KEYINPUT35), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G232gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT34), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI22_X1  g317(.A1(new_n426_), .A2(new_n466_), .B1(new_n515_), .B2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n468_), .A2(new_n413_), .A3(new_n469_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n518_), .A2(new_n515_), .ZN(new_n522_));
  AND2_X1   g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n521_), .A2(new_n522_), .ZN(new_n524_));
  NOR2_X1   g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G190gat), .B(G218gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT72), .ZN(new_n527_));
  XNOR2_X1  g326(.A(G134gat), .B(G162gat), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n527_), .B(new_n528_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n529_), .A2(KEYINPUT36), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n525_), .A2(new_n530_), .ZN(new_n531_));
  XOR2_X1   g330(.A(new_n529_), .B(KEYINPUT36), .Z(new_n532_));
  OAI21_X1  g331(.A(new_n532_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(KEYINPUT37), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n533_), .A2(KEYINPUT74), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT73), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n531_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n525_), .A2(KEYINPUT73), .A3(new_n530_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n533_), .A2(KEYINPUT74), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n536_), .A2(new_n538_), .A3(new_n539_), .A4(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n535_), .B1(new_n541_), .B2(KEYINPUT37), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G231gat), .A2(G233gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n410_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(new_n482_), .ZN(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G127gat), .B(G155gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G183gat), .B(G211gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n550_), .B(new_n551_), .ZN(new_n552_));
  OR3_X1    g351(.A1(new_n546_), .A2(new_n547_), .A3(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(KEYINPUT17), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n546_), .A2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n542_), .A2(new_n556_), .ZN(new_n557_));
  AND2_X1   g356(.A1(new_n514_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n433_), .A2(new_n558_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(KEYINPUT99), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT99), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n433_), .A2(new_n561_), .A3(new_n558_), .ZN(new_n562_));
  AND2_X1   g361(.A1(new_n560_), .A2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(new_n402_), .A3(new_n384_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT38), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n563_), .A2(KEYINPUT38), .A3(new_n402_), .A4(new_n384_), .ZN(new_n567_));
  AND2_X1   g366(.A1(new_n395_), .A2(new_n534_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n513_), .A2(new_n432_), .ZN(new_n569_));
  NOR2_X1   g368(.A1(new_n569_), .A2(new_n556_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(G1gat), .B1(new_n571_), .B2(new_n360_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n566_), .A2(new_n567_), .A3(new_n572_), .ZN(G1324gat));
  XOR2_X1   g372(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT100), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n568_), .A2(new_n284_), .A3(new_n570_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT39), .ZN(new_n577_));
  AND3_X1   g376(.A1(new_n576_), .A2(new_n577_), .A3(G8gat), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n577_), .B1(new_n576_), .B2(G8gat), .ZN(new_n579_));
  OR2_X1    g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n560_), .A2(new_n403_), .A3(new_n284_), .A4(new_n562_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n575_), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n581_), .B(new_n575_), .C1(new_n578_), .C2(new_n579_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n582_), .A2(new_n584_), .ZN(G1325gat));
  INV_X1    g384(.A(new_n371_), .ZN(new_n586_));
  OAI21_X1  g385(.A(G15gat), .B1(new_n571_), .B2(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT41), .ZN(new_n588_));
  NOR3_X1   g387(.A1(new_n559_), .A2(G15gat), .A3(new_n586_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n588_), .A2(new_n589_), .ZN(G1326gat));
  AND2_X1   g389(.A1(new_n329_), .A2(new_n333_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n568_), .A2(new_n591_), .A3(new_n570_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT42), .ZN(new_n593_));
  AND3_X1   g392(.A1(new_n592_), .A2(new_n593_), .A3(G22gat), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n593_), .B1(new_n592_), .B2(G22gat), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n334_), .A2(G22gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n596_), .B(KEYINPUT102), .Z(new_n597_));
  OAI22_X1  g396(.A1(new_n594_), .A2(new_n595_), .B1(new_n559_), .B2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT103), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n598_), .B(new_n599_), .ZN(G1327gat));
  INV_X1    g399(.A(new_n556_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n569_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n542_), .A2(KEYINPUT104), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT43), .ZN(new_n604_));
  AND3_X1   g403(.A1(new_n395_), .A2(new_n542_), .A3(new_n604_), .ZN(new_n605_));
  AOI21_X1  g404(.A(new_n604_), .B1(new_n395_), .B2(new_n542_), .ZN(new_n606_));
  OAI211_X1 g405(.A(KEYINPUT44), .B(new_n602_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n602_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n395_), .A2(new_n542_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n604_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n395_), .A2(new_n542_), .A3(new_n604_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n608_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n614_));
  OAI21_X1  g413(.A(new_n607_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n384_), .A2(G29gat), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n513_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n534_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n556_), .A2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  AND2_X1   g421(.A1(new_n433_), .A2(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(G29gat), .B1(new_n623_), .B2(new_n384_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n618_), .A2(new_n624_), .ZN(G1328gat));
  INV_X1    g424(.A(KEYINPUT46), .ZN(new_n626_));
  AOI21_X1  g425(.A(KEYINPUT107), .B1(new_n626_), .B2(KEYINPUT106), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT108), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n607_), .B(new_n284_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(G36gat), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n626_), .A2(KEYINPUT107), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n285_), .A2(G36gat), .ZN(new_n632_));
  NAND4_X1  g431(.A1(new_n395_), .A2(new_n432_), .A3(new_n622_), .A4(new_n632_), .ZN(new_n633_));
  AND2_X1   g432(.A1(new_n633_), .A2(KEYINPUT45), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(KEYINPUT45), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n631_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n628_), .B1(new_n630_), .B2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n628_), .ZN(new_n639_));
  AOI211_X1 g438(.A(new_n639_), .B(new_n636_), .C1(new_n629_), .C2(G36gat), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n638_), .A2(new_n640_), .ZN(G1329gat));
  NAND2_X1  g440(.A1(new_n623_), .A2(new_n371_), .ZN(new_n642_));
  INV_X1    g441(.A(G43gat), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n371_), .A2(G43gat), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n644_), .B1(new_n615_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g446(.A1(new_n334_), .A2(G50gat), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT110), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n623_), .A2(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n607_), .B(new_n591_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n651_), .A2(KEYINPUT109), .ZN(new_n652_));
  OAI21_X1  g451(.A(G50gat), .B1(new_n651_), .B2(KEYINPUT109), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n650_), .B1(new_n652_), .B2(new_n653_), .ZN(G1331gat));
  INV_X1    g453(.A(new_n432_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n395_), .A2(new_n655_), .ZN(new_n656_));
  NOR4_X1   g455(.A1(new_n656_), .A2(new_n513_), .A3(new_n556_), .A4(new_n542_), .ZN(new_n657_));
  INV_X1    g456(.A(G57gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(new_n658_), .A3(new_n384_), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n514_), .A2(new_n432_), .A3(new_n556_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n568_), .A2(new_n660_), .ZN(new_n661_));
  OAI21_X1  g460(.A(G57gat), .B1(new_n661_), .B2(new_n360_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n659_), .A2(new_n662_), .ZN(G1332gat));
  OAI21_X1  g462(.A(G64gat), .B1(new_n661_), .B2(new_n285_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT48), .ZN(new_n665_));
  INV_X1    g464(.A(G64gat), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n657_), .A2(new_n666_), .A3(new_n284_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1333gat));
  INV_X1    g467(.A(G71gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n657_), .A2(new_n669_), .A3(new_n371_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G71gat), .B1(new_n661_), .B2(new_n586_), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n671_), .A2(KEYINPUT49), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n671_), .A2(KEYINPUT49), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n670_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT111), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT111), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n676_), .B(new_n670_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1334gat));
  OAI21_X1  g477(.A(G78gat), .B1(new_n661_), .B2(new_n334_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT50), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n657_), .A2(new_n476_), .A3(new_n591_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1335gat));
  NOR3_X1   g481(.A1(new_n513_), .A2(new_n432_), .A3(new_n601_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n683_), .B(KEYINPUT112), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n684_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n685_));
  OAI21_X1  g484(.A(G85gat), .B1(new_n685_), .B2(new_n360_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n656_), .A2(new_n514_), .A3(new_n621_), .ZN(new_n687_));
  INV_X1    g486(.A(G85gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n384_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n686_), .A2(new_n689_), .ZN(G1336gat));
  OAI21_X1  g489(.A(G92gat), .B1(new_n685_), .B2(new_n285_), .ZN(new_n691_));
  INV_X1    g490(.A(G92gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n687_), .A2(new_n692_), .A3(new_n284_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n691_), .A2(new_n693_), .ZN(G1337gat));
  OAI211_X1 g493(.A(new_n371_), .B(new_n684_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n371_), .A2(new_n461_), .ZN(new_n696_));
  AOI22_X1  g495(.A1(new_n695_), .A2(G99gat), .B1(new_n687_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT114), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT113), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n699_), .A2(KEYINPUT51), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n697_), .A2(new_n698_), .A3(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n697_), .A2(new_n698_), .ZN(new_n702_));
  OAI21_X1  g501(.A(KEYINPUT51), .B1(new_n697_), .B2(new_n699_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n701_), .B1(new_n702_), .B2(new_n703_), .ZN(G1338gat));
  NAND3_X1  g503(.A1(new_n687_), .A2(new_n445_), .A3(new_n591_), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n591_), .B(new_n684_), .C1(new_n605_), .C2(new_n606_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT52), .ZN(new_n707_));
  AND3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(G106gat), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n707_), .B1(new_n706_), .B2(G106gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT53), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT53), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n712_), .B(new_n705_), .C1(new_n708_), .C2(new_n709_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1339gat));
  NAND4_X1  g513(.A1(new_n285_), .A2(new_n334_), .A3(new_n384_), .A4(new_n371_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n432_), .B1(new_n506_), .B2(new_n502_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT55), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n483_), .B(new_n490_), .C1(new_n495_), .C2(KEYINPUT12), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n718_), .B2(new_n486_), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n718_), .A2(new_n486_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(new_n720_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n718_), .A2(new_n717_), .A3(new_n486_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n502_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT56), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n485_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n492_), .B1(new_n726_), .B2(new_n717_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n722_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n729_), .A2(KEYINPUT56), .A3(new_n502_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n716_), .B1(new_n725_), .B2(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n418_), .B1(new_n427_), .B2(new_n397_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n732_), .A2(new_n431_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n423_), .A2(new_n424_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(new_n414_), .ZN(new_n735_));
  MUX2_X1   g534(.A(new_n427_), .B(new_n735_), .S(new_n396_), .Z(new_n736_));
  OAI21_X1  g535(.A(new_n733_), .B1(new_n736_), .B2(new_n431_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n504_), .B2(new_n507_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n534_), .B1(new_n731_), .B2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT57), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n737_), .B1(new_n497_), .B2(new_n503_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT56), .B1(new_n729_), .B2(new_n502_), .ZN(new_n743_));
  AOI211_X1 g542(.A(new_n724_), .B(new_n503_), .C1(new_n727_), .C2(new_n728_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n742_), .B1(new_n743_), .B2(new_n744_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(KEYINPUT115), .A2(KEYINPUT58), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n746_), .ZN(new_n748_));
  OAI211_X1 g547(.A(new_n742_), .B(new_n748_), .C1(new_n743_), .C2(new_n744_), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n747_), .A2(new_n542_), .A3(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(KEYINPUT57), .B(new_n534_), .C1(new_n731_), .C2(new_n738_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n741_), .A2(new_n750_), .A3(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT116), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n741_), .A2(new_n750_), .A3(KEYINPUT116), .A4(new_n751_), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n754_), .A2(new_n556_), .A3(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n513_), .A2(new_n557_), .A3(new_n655_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(KEYINPUT54), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n759_));
  NAND4_X1  g558(.A1(new_n513_), .A2(new_n557_), .A3(new_n759_), .A4(new_n655_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n758_), .A2(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n715_), .B1(new_n756_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(G113gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n762_), .A2(new_n763_), .A3(new_n432_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n601_), .B1(new_n752_), .B2(new_n753_), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n765_), .A2(new_n755_), .B1(new_n758_), .B2(new_n760_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT59), .B1(new_n766_), .B2(new_n715_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n752_), .A2(new_n556_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n761_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT59), .ZN(new_n770_));
  OR2_X1    g569(.A1(new_n715_), .A2(KEYINPUT117), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n715_), .A2(KEYINPUT117), .ZN(new_n772_));
  NAND4_X1  g571(.A1(new_n769_), .A2(new_n770_), .A3(new_n771_), .A4(new_n772_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n767_), .A2(new_n773_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(new_n432_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n764_), .B1(new_n776_), .B2(new_n763_), .ZN(G1340gat));
  INV_X1    g576(.A(new_n514_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n778_), .B(new_n773_), .C1(new_n762_), .C2(new_n770_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n779_), .A2(KEYINPUT118), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT118), .ZN(new_n781_));
  NAND4_X1  g580(.A1(new_n767_), .A2(new_n781_), .A3(new_n778_), .A4(new_n773_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(G120gat), .A3(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(G120gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n513_), .B2(KEYINPUT60), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n762_), .B(new_n785_), .C1(KEYINPUT60), .C2(new_n784_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n783_), .A2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT119), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n783_), .A2(KEYINPUT119), .A3(new_n786_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1341gat));
  INV_X1    g590(.A(G127gat), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n762_), .A2(new_n792_), .A3(new_n601_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n774_), .A2(new_n601_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n793_), .B1(new_n795_), .B2(new_n792_), .ZN(G1342gat));
  INV_X1    g595(.A(G134gat), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n762_), .A2(new_n797_), .A3(new_n620_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n774_), .A2(new_n542_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n798_), .B1(new_n800_), .B2(new_n797_), .ZN(G1343gat));
  NAND2_X1  g600(.A1(new_n756_), .A2(new_n761_), .ZN(new_n802_));
  NOR2_X1   g601(.A1(new_n334_), .A2(new_n371_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n284_), .A2(new_n360_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n802_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT120), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT120), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n802_), .A2(new_n807_), .A3(new_n803_), .A4(new_n804_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n432_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g610(.A1(new_n809_), .A2(new_n778_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g612(.A(KEYINPUT61), .B(G155gat), .ZN(new_n814_));
  INV_X1    g613(.A(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT121), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n816_), .B1(new_n809_), .B2(new_n601_), .ZN(new_n817_));
  AOI211_X1 g616(.A(KEYINPUT121), .B(new_n556_), .C1(new_n806_), .C2(new_n808_), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n815_), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n803_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n766_), .A2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n807_), .B1(new_n821_), .B2(new_n804_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n808_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n601_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT121), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n809_), .A2(new_n816_), .A3(new_n601_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n825_), .A2(new_n826_), .A3(new_n814_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n819_), .A2(new_n827_), .ZN(G1346gat));
  INV_X1    g627(.A(new_n809_), .ZN(new_n829_));
  OR3_X1    g628(.A1(new_n829_), .A2(G162gat), .A3(new_n534_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n542_), .ZN(new_n831_));
  OAI21_X1  g630(.A(G162gat), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1347gat));
  NOR2_X1   g632(.A1(new_n285_), .A2(new_n384_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(new_n371_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n769_), .A2(new_n334_), .A3(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n432_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(G169gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n837_), .A2(new_n655_), .ZN(new_n842_));
  AOI22_X1  g641(.A1(new_n840_), .A2(new_n841_), .B1(new_n842_), .B2(new_n210_), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n840_), .B2(new_n841_), .ZN(G1348gat));
  OAI21_X1  g643(.A(new_n208_), .B1(new_n837_), .B2(new_n513_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n845_), .B(KEYINPUT123), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n766_), .A2(new_n591_), .ZN(new_n847_));
  NOR3_X1   g646(.A1(new_n514_), .A2(new_n208_), .A3(new_n835_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n846_), .B1(new_n847_), .B2(new_n848_), .ZN(G1349gat));
  NAND3_X1  g648(.A1(new_n847_), .A2(new_n601_), .A3(new_n836_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n601_), .A2(new_n219_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n850_), .A2(new_n241_), .B1(new_n838_), .B2(new_n851_), .ZN(G1350gat));
  OAI21_X1  g651(.A(G190gat), .B1(new_n837_), .B2(new_n831_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n620_), .A2(new_n217_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n837_), .B2(new_n854_), .ZN(new_n855_));
  XOR2_X1   g654(.A(new_n855_), .B(KEYINPUT124), .Z(G1351gat));
  AND3_X1   g655(.A1(new_n802_), .A2(new_n803_), .A3(new_n834_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n432_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g658(.A(G204gat), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n857_), .B(new_n778_), .C1(KEYINPUT125), .C2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(KEYINPUT125), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1353gat));
  AOI21_X1  g662(.A(new_n556_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n857_), .A2(new_n864_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT126), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT126), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n857_), .A2(new_n867_), .A3(new_n864_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n866_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n869_), .B(new_n870_), .ZN(G1354gat));
  AND3_X1   g670(.A1(new_n857_), .A2(G218gat), .A3(new_n542_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n857_), .A2(new_n620_), .ZN(new_n873_));
  OR2_X1    g672(.A1(new_n873_), .A2(KEYINPUT127), .ZN(new_n874_));
  AOI21_X1  g673(.A(G218gat), .B1(new_n873_), .B2(KEYINPUT127), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n872_), .B1(new_n874_), .B2(new_n875_), .ZN(G1355gat));
endmodule


