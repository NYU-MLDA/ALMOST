//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n829_, new_n830_, new_n831_, new_n832_, new_n833_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n909_, new_n911_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n938_, new_n940_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT8), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G99gat), .A2(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT6), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n208_));
  NAND3_X1  g007(.A1(new_n206_), .A2(new_n207_), .A3(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT7), .ZN(new_n210_));
  INV_X1    g009(.A(G99gat), .ZN(new_n211_));
  INV_X1    g010(.A(G106gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n210_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT68), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT68), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(new_n210_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n209_), .B1(new_n214_), .B2(new_n217_), .ZN(new_n218_));
  AND2_X1   g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G85gat), .A2(G92gat), .ZN(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT69), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(G85gat), .ZN(new_n222_));
  INV_X1    g021(.A(G92gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT69), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G85gat), .A2(G92gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n224_), .A2(new_n225_), .A3(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n221_), .A2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n203_), .B1(new_n218_), .B2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n203_), .B1(new_n221_), .B2(new_n227_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n204_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT70), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n232_), .A2(KEYINPUT6), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n205_), .A2(KEYINPUT70), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n231_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n205_), .A2(KEYINPUT70), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(KEYINPUT6), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n204_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n235_), .A2(new_n208_), .A3(new_n238_), .ZN(new_n239_));
  NOR4_X1   g038(.A1(KEYINPUT68), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n216_), .B1(new_n215_), .B2(new_n210_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n230_), .B1(new_n239_), .B2(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n223_), .A2(KEYINPUT65), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G92gat), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n222_), .B1(new_n245_), .B2(new_n247_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n244_), .B1(new_n248_), .B2(KEYINPUT9), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT9), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT65), .B(G92gat), .ZN(new_n251_));
  OAI211_X1 g050(.A(KEYINPUT66), .B(new_n250_), .C1(new_n251_), .C2(new_n222_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n219_), .A2(KEYINPUT67), .A3(KEYINPUT9), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n219_), .A2(KEYINPUT9), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n224_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  AOI22_X1  g055(.A1(new_n249_), .A2(new_n252_), .B1(new_n253_), .B2(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n206_), .A2(new_n207_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT64), .ZN(new_n260_));
  XOR2_X1   g059(.A(KEYINPUT10), .B(G99gat), .Z(new_n261_));
  AOI21_X1  g060(.A(new_n260_), .B1(new_n261_), .B2(new_n212_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT10), .B(G99gat), .ZN(new_n263_));
  NOR3_X1   g062(.A1(new_n263_), .A2(KEYINPUT64), .A3(G106gat), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n259_), .B1(new_n262_), .B2(new_n264_), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n229_), .B(new_n243_), .C1(new_n257_), .C2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT71), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n256_), .A2(new_n253_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n245_), .A2(new_n247_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(G85gat), .ZN(new_n271_));
  AOI21_X1  g070(.A(KEYINPUT66), .B1(new_n271_), .B2(new_n250_), .ZN(new_n272_));
  NOR3_X1   g071(.A1(new_n248_), .A2(new_n244_), .A3(KEYINPUT9), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n269_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n264_), .ZN(new_n275_));
  OAI21_X1  g074(.A(KEYINPUT64), .B1(new_n263_), .B2(G106gat), .ZN(new_n276_));
  AOI21_X1  g075(.A(new_n258_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n274_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n221_), .A2(new_n227_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(new_n242_), .B2(new_n209_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n208_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT70), .B(KEYINPUT6), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n281_), .B1(new_n282_), .B2(new_n204_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n214_), .A2(new_n217_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(new_n235_), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n203_), .A2(new_n280_), .B1(new_n285_), .B2(new_n230_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n278_), .A2(new_n286_), .A3(KEYINPUT71), .ZN(new_n287_));
  INV_X1    g086(.A(G36gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(G29gat), .ZN(new_n289_));
  INV_X1    g088(.A(G29gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(G36gat), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n292_));
  AND3_X1   g091(.A1(new_n289_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n292_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n294_));
  OAI21_X1  g093(.A(G43gat), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n290_), .A2(G36gat), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n288_), .A2(G29gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(KEYINPUT73), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(G43gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n289_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n298_), .A2(new_n299_), .A3(new_n300_), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n295_), .A2(new_n301_), .A3(G50gat), .ZN(new_n302_));
  AOI21_X1  g101(.A(G50gat), .B1(new_n295_), .B2(new_n301_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n268_), .A2(new_n287_), .A3(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(KEYINPUT74), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n307_));
  NAND4_X1  g106(.A1(new_n268_), .A2(new_n287_), .A3(new_n307_), .A4(new_n304_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(G50gat), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n293_), .A2(new_n294_), .A3(G43gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n299_), .B1(new_n298_), .B2(new_n300_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n310_), .B1(new_n311_), .B2(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n295_), .A2(new_n301_), .A3(G50gat), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n313_), .A2(KEYINPUT15), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(KEYINPUT15), .B1(new_n313_), .B2(new_n314_), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n266_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G232gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT34), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(KEYINPUT35), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n319_), .A2(KEYINPUT35), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n317_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n309_), .A2(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(G134gat), .B(G162gat), .Z(new_n327_));
  XNOR2_X1  g126(.A(G190gat), .B(G218gat), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n327_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(KEYINPUT77), .B(KEYINPUT36), .Z(new_n333_));
  NOR2_X1   g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n326_), .A2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n320_), .B1(new_n309_), .B2(new_n317_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n202_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n309_), .A2(new_n317_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n321_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n324_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n334_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(KEYINPUT78), .A3(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n337_), .A2(new_n343_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n339_), .A2(new_n326_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT80), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n331_), .B(KEYINPUT36), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n347_), .B1(new_n336_), .B2(new_n340_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT80), .ZN(new_n350_));
  XOR2_X1   g149(.A(KEYINPUT81), .B(KEYINPUT37), .Z(new_n351_));
  AND4_X1   g150(.A1(new_n344_), .A2(new_n348_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT79), .ZN(new_n353_));
  AOI22_X1  g152(.A1(new_n337_), .A2(new_n343_), .B1(new_n345_), .B2(new_n347_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT37), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n335_), .A2(new_n202_), .A3(new_n336_), .ZN(new_n357_));
  AOI21_X1  g156(.A(KEYINPUT78), .B1(new_n339_), .B2(new_n342_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n349_), .B1(new_n357_), .B2(new_n358_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(KEYINPUT79), .A3(KEYINPUT37), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n352_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G127gat), .B(G134gat), .Z(new_n362_));
  XOR2_X1   g161(.A(G113gat), .B(G120gat), .Z(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT31), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT30), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G183gat), .A2(G190gat), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n368_), .A2(KEYINPUT23), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT23), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n370_), .A2(G183gat), .A3(G190gat), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT84), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n369_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  OR2_X1    g172(.A1(G183gat), .A2(G190gat), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n368_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n373_), .A2(new_n374_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G169gat), .A2(G176gat), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT22), .B(G169gat), .ZN(new_n379_));
  INV_X1    g178(.A(G176gat), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n378_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n376_), .A2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(KEYINPUT25), .B(G183gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT26), .B(G190gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n369_), .A2(new_n371_), .ZN(new_n386_));
  OR3_X1    g185(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n387_));
  INV_X1    g186(.A(G169gat), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n380_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(KEYINPUT24), .A3(new_n377_), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n385_), .A2(new_n386_), .A3(new_n387_), .A4(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n382_), .A2(KEYINPUT85), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(KEYINPUT85), .B1(new_n382_), .B2(new_n391_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n367_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n394_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(KEYINPUT30), .A3(new_n392_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G15gat), .B(G43gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399_));
  XNOR2_X1  g198(.A(new_n398_), .B(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G71gat), .B(G99gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n395_), .A2(new_n397_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT86), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n402_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n366_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n406_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n408_), .A2(new_n404_), .A3(new_n403_), .A4(new_n365_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G78gat), .B(G106gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT29), .ZN(new_n413_));
  XOR2_X1   g212(.A(G155gat), .B(G162gat), .Z(new_n414_));
  OR3_X1    g213(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT2), .ZN(new_n417_));
  AOI21_X1  g216(.A(KEYINPUT87), .B1(G141gat), .B2(G148gat), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n415_), .B(new_n416_), .C1(new_n417_), .C2(new_n418_), .ZN(new_n419_));
  AND2_X1   g218(.A1(new_n418_), .A2(new_n417_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n414_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT1), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n414_), .A2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(G141gat), .B(G148gat), .Z(new_n425_));
  NAND3_X1  g224(.A1(new_n423_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n413_), .B1(new_n421_), .B2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT90), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT89), .ZN(new_n429_));
  INV_X1    g228(.A(G197gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n429_), .B1(new_n430_), .B2(G204gat), .ZN(new_n431_));
  INV_X1    g230(.A(G204gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT21), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(G204gat), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n431_), .A2(new_n433_), .A3(new_n434_), .A4(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(G211gat), .B(G218gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G197gat), .B(G204gat), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n438_), .B1(new_n439_), .B2(new_n434_), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n428_), .B1(new_n437_), .B2(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n435_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n430_), .A2(G204gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT21), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  NAND4_X1  g243(.A1(new_n444_), .A2(new_n436_), .A3(KEYINPUT90), .A4(new_n438_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n431_), .A2(new_n435_), .A3(new_n433_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n438_), .A2(new_n434_), .ZN(new_n447_));
  AOI22_X1  g246(.A1(new_n441_), .A2(new_n445_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n448_));
  AND2_X1   g247(.A1(G228gat), .A2(G233gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  AOI211_X1 g249(.A(new_n427_), .B(new_n448_), .C1(KEYINPUT88), .C2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n450_), .B1(new_n448_), .B2(KEYINPUT88), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n448_), .A2(new_n427_), .ZN(new_n453_));
  NOR2_X1   g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n412_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT91), .ZN(new_n456_));
  INV_X1    g255(.A(new_n427_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n441_), .A2(new_n445_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n447_), .A2(new_n446_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n461_), .A2(new_n463_), .A3(new_n450_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n452_), .A2(new_n453_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n464_), .A2(new_n411_), .A3(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n421_), .A2(new_n426_), .ZN(new_n467_));
  NOR2_X1   g266(.A1(new_n467_), .A2(KEYINPUT29), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G22gat), .B(G50gat), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n469_), .B(KEYINPUT28), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n468_), .B(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n455_), .A2(new_n456_), .A3(new_n466_), .A4(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n466_), .A2(KEYINPUT91), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n474_), .A2(new_n471_), .B1(new_n455_), .B2(new_n466_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n410_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G225gat), .A2(G233gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT4), .ZN(new_n479_));
  INV_X1    g278(.A(new_n467_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT96), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n364_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n364_), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n483_), .B1(new_n467_), .B2(KEYINPUT96), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n479_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n480_), .A2(new_n483_), .A3(KEYINPUT4), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n478_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n482_), .A2(new_n484_), .A3(new_n477_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G57gat), .B(G85gat), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G1gat), .B(G29gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  XNOR2_X1  g291(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n489_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT33), .ZN(new_n497_));
  OR3_X1    g296(.A1(new_n485_), .A2(new_n478_), .A3(new_n486_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n482_), .A2(new_n484_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n495_), .B1(new_n499_), .B2(new_n478_), .ZN(new_n500_));
  AOI22_X1  g299(.A1(new_n496_), .A2(new_n497_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G8gat), .B(G36gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT18), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(G64gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(new_n223_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n373_), .A2(new_n375_), .A3(new_n387_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT93), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  XOR2_X1   g308(.A(KEYINPUT26), .B(G190gat), .Z(new_n510_));
  INV_X1    g309(.A(KEYINPUT92), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n384_), .A2(KEYINPUT92), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n383_), .A3(new_n513_), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n373_), .A2(KEYINPUT93), .A3(new_n375_), .A4(new_n387_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n509_), .A2(new_n514_), .A3(new_n390_), .A4(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n386_), .A2(new_n374_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n381_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n448_), .A2(new_n516_), .A3(new_n518_), .ZN(new_n519_));
  AND2_X1   g318(.A1(new_n519_), .A2(KEYINPUT20), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G226gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT19), .ZN(new_n522_));
  INV_X1    g321(.A(new_n522_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n460_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n520_), .A2(KEYINPUT95), .A3(new_n523_), .A4(new_n524_), .ZN(new_n525_));
  NAND4_X1  g324(.A1(new_n524_), .A2(KEYINPUT20), .A3(new_n523_), .A4(new_n519_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n525_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT20), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n516_), .A2(new_n518_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n531_), .B1(new_n532_), .B2(new_n460_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n396_), .A2(new_n448_), .A3(new_n392_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n523_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n535_), .A2(KEYINPUT94), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT94), .ZN(new_n537_));
  AOI211_X1 g336(.A(new_n537_), .B(new_n523_), .C1(new_n533_), .C2(new_n534_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n506_), .B1(new_n530_), .B2(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n529_), .B(new_n505_), .C1(new_n536_), .C2(new_n538_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n489_), .A2(KEYINPUT33), .A3(new_n495_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n501_), .A2(new_n540_), .A3(new_n541_), .A4(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT98), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n544_), .B1(new_n489_), .B2(new_n495_), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n487_), .A2(new_n488_), .A3(KEYINPUT98), .A4(new_n494_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n545_), .A2(new_n546_), .A3(new_n496_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n535_), .B(KEYINPUT94), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n505_), .A2(KEYINPUT32), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n529_), .A3(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n533_), .A2(new_n523_), .A3(new_n534_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n524_), .A2(KEYINPUT20), .A3(new_n519_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(new_n523_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n553_), .A2(KEYINPUT32), .A3(new_n505_), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n547_), .A2(new_n550_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n476_), .B1(new_n543_), .B2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT27), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n557_), .B1(new_n553_), .B2(new_n506_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n541_), .A2(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT99), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n541_), .A2(KEYINPUT99), .A3(new_n558_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  AND2_X1   g362(.A1(new_n407_), .A2(new_n409_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n474_), .A2(new_n471_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n455_), .A2(new_n466_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n568_), .A2(new_n472_), .A3(new_n410_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n547_), .B1(new_n565_), .B2(new_n569_), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n563_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n541_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n505_), .B1(new_n548_), .B2(new_n529_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n557_), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT100), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n540_), .A2(new_n541_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n577_), .A2(KEYINPUT100), .A3(new_n557_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n576_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n556_), .B1(new_n571_), .B2(new_n579_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n361_), .A2(new_n580_), .ZN(new_n581_));
  AND2_X1   g380(.A1(G230gat), .A2(G233gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(G71gat), .B(G78gat), .Z(new_n583_));
  XNOR2_X1  g382(.A(G57gat), .B(G64gat), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n583_), .B1(KEYINPUT11), .B2(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(KEYINPUT11), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n585_), .B(new_n586_), .Z(new_n587_));
  NAND3_X1  g386(.A1(new_n268_), .A2(new_n287_), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n587_), .B1(new_n268_), .B2(new_n287_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n582_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n266_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT12), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n587_), .A2(new_n593_), .ZN(new_n594_));
  OAI221_X1 g393(.A(new_n588_), .B1(new_n592_), .B2(new_n594_), .C1(new_n590_), .C2(KEYINPUT12), .ZN(new_n595_));
  OAI21_X1  g394(.A(new_n591_), .B1(new_n595_), .B2(new_n582_), .ZN(new_n596_));
  XOR2_X1   g395(.A(KEYINPUT72), .B(KEYINPUT5), .Z(new_n597_));
  XNOR2_X1  g396(.A(G120gat), .B(G148gat), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n599_), .B(new_n600_), .Z(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n596_), .A2(new_n602_), .ZN(new_n603_));
  OAI211_X1 g402(.A(new_n591_), .B(new_n601_), .C1(new_n595_), .C2(new_n582_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT13), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n603_), .A2(KEYINPUT13), .A3(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G15gat), .B(G22gat), .ZN(new_n611_));
  INV_X1    g410(.A(G1gat), .ZN(new_n612_));
  INV_X1    g411(.A(G8gat), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT14), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G1gat), .B(G8gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n615_), .B(new_n616_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n617_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n618_), .A2(KEYINPUT82), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(KEYINPUT82), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n304_), .ZN(new_n622_));
  OR2_X1    g421(.A1(new_n622_), .A2(new_n617_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(G229gat), .A2(G233gat), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n621_), .A2(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n622_), .A2(new_n617_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n623_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n624_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(G113gat), .B(G141gat), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(G169gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(new_n430_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n627_), .A2(new_n631_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n634_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n625_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n631_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n636_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT83), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n635_), .A2(new_n639_), .A3(new_n640_), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n640_), .B1(new_n635_), .B2(new_n639_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n610_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n617_), .B(new_n646_), .ZN(new_n647_));
  XOR2_X1   g446(.A(new_n647_), .B(new_n587_), .Z(new_n648_));
  XNOR2_X1  g447(.A(G127gat), .B(G155gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT16), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(G183gat), .ZN(new_n651_));
  INV_X1    g450(.A(G211gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n651_), .B(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT17), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n653_), .A2(new_n654_), .ZN(new_n656_));
  OR3_X1    g455(.A1(new_n648_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n648_), .A2(new_n656_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n645_), .A2(new_n659_), .ZN(new_n660_));
  AND2_X1   g459(.A1(new_n581_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n612_), .A3(new_n547_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n663_), .A2(KEYINPUT38), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT101), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n344_), .A2(new_n348_), .A3(new_n350_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n580_), .A2(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n668_), .A2(new_n660_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n612_), .B1(new_n669_), .B2(new_n547_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n663_), .B2(KEYINPUT38), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n665_), .A2(new_n671_), .ZN(G1324gat));
  NAND2_X1  g471(.A1(new_n579_), .A2(new_n563_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n613_), .B1(new_n669_), .B2(new_n673_), .ZN(new_n674_));
  XOR2_X1   g473(.A(new_n674_), .B(KEYINPUT39), .Z(new_n675_));
  NAND3_X1  g474(.A1(new_n661_), .A2(new_n613_), .A3(new_n673_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n678_));
  XNOR2_X1  g477(.A(new_n677_), .B(new_n678_), .ZN(G1325gat));
  NAND2_X1  g478(.A1(new_n669_), .A2(new_n564_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n680_), .A2(G15gat), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT102), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n680_), .A2(new_n683_), .A3(G15gat), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(G15gat), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n661_), .A2(new_n688_), .A3(new_n564_), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n682_), .A2(KEYINPUT41), .A3(new_n684_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n687_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(KEYINPUT103), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n687_), .A2(new_n693_), .A3(new_n689_), .A4(new_n690_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n692_), .A2(new_n694_), .ZN(G1326gat));
  INV_X1    g494(.A(G22gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n473_), .A2(new_n475_), .ZN(new_n697_));
  NAND3_X1  g496(.A1(new_n661_), .A2(new_n696_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n696_), .B1(new_n669_), .B2(new_n697_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT104), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n700_), .A2(KEYINPUT42), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(KEYINPUT42), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n701_), .B2(new_n702_), .ZN(G1327gat));
  NAND3_X1  g502(.A1(new_n610_), .A2(new_n644_), .A3(new_n659_), .ZN(new_n704_));
  NOR3_X1   g503(.A1(new_n580_), .A2(new_n704_), .A3(new_n666_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G29gat), .B1(new_n705_), .B2(new_n547_), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n344_), .A2(new_n348_), .A3(new_n350_), .A4(new_n351_), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n354_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n708_));
  AOI21_X1  g507(.A(KEYINPUT79), .B1(new_n359_), .B2(KEYINPUT37), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n707_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(KEYINPUT43), .B1(new_n710_), .B2(new_n580_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n556_), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT100), .B1(new_n577_), .B2(new_n557_), .ZN(new_n713_));
  AOI211_X1 g512(.A(new_n575_), .B(KEYINPUT27), .C1(new_n540_), .C2(new_n541_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n713_), .A2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n563_), .A2(new_n570_), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT43), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n361_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n711_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n704_), .ZN(new_n721_));
  AND4_X1   g520(.A1(KEYINPUT105), .A2(new_n720_), .A3(KEYINPUT44), .A4(new_n721_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n704_), .B1(new_n711_), .B2(new_n719_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT105), .B1(new_n723_), .B2(KEYINPUT44), .ZN(new_n724_));
  OR2_X1    g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n723_), .A2(KEYINPUT44), .ZN(new_n726_));
  INV_X1    g525(.A(new_n547_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n726_), .A2(new_n290_), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n706_), .B1(new_n725_), .B2(new_n728_), .ZN(G1328gat));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n705_), .A2(new_n288_), .A3(new_n673_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT45), .Z(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n673_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n726_), .A2(new_n736_), .ZN(new_n737_));
  AND2_X1   g536(.A1(new_n725_), .A2(new_n737_), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n732_), .B(new_n735_), .C1(new_n738_), .C2(new_n288_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n288_), .B1(new_n725_), .B2(new_n737_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n730_), .B(new_n731_), .C1(new_n740_), .C2(new_n734_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(G1329gat));
  XNOR2_X1  g541(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n564_), .A2(G43gat), .ZN(new_n744_));
  AND3_X1   g543(.A1(new_n361_), .A2(new_n718_), .A3(new_n717_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n718_), .B1(new_n361_), .B2(new_n717_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n721_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT44), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT107), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT107), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n752_), .B(new_n749_), .C1(new_n722_), .C2(new_n724_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(G43gat), .B1(new_n705_), .B2(new_n564_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n743_), .B1(new_n754_), .B2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n743_), .ZN(new_n758_));
  AOI211_X1 g557(.A(new_n758_), .B(new_n755_), .C1(new_n751_), .C2(new_n753_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n757_), .A2(new_n759_), .ZN(G1330gat));
  AOI21_X1  g559(.A(G50gat), .B1(new_n705_), .B2(new_n697_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n697_), .ZN(new_n762_));
  NOR3_X1   g561(.A1(new_n726_), .A2(new_n310_), .A3(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n761_), .B1(new_n725_), .B2(new_n763_), .ZN(G1331gat));
  NOR3_X1   g563(.A1(new_n610_), .A2(new_n644_), .A3(new_n659_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n668_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n766_), .B(new_n767_), .ZN(new_n768_));
  XOR2_X1   g567(.A(KEYINPUT110), .B(G57gat), .Z(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(new_n547_), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n771_));
  OR2_X1    g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(G57gat), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n581_), .A2(new_n765_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(new_n727_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n770_), .A2(new_n771_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n772_), .A2(new_n775_), .A3(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n772_), .A2(KEYINPUT112), .A3(new_n775_), .A4(new_n776_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(G1332gat));
  INV_X1    g580(.A(G64gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n768_), .B2(new_n673_), .ZN(new_n783_));
  XOR2_X1   g582(.A(new_n783_), .B(KEYINPUT48), .Z(new_n784_));
  INV_X1    g583(.A(new_n774_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n785_), .A2(new_n782_), .A3(new_n673_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1333gat));
  INV_X1    g586(.A(G71gat), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(new_n788_), .A3(new_n564_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n768_), .A2(new_n564_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n790_), .B1(new_n791_), .B2(G71gat), .ZN(new_n792_));
  AOI211_X1 g591(.A(KEYINPUT49), .B(new_n788_), .C1(new_n768_), .C2(new_n564_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n789_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT113), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  OAI211_X1 g595(.A(KEYINPUT113), .B(new_n789_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(G1334gat));
  NAND2_X1  g597(.A1(new_n768_), .A2(new_n697_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(G78gat), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n800_), .B(new_n801_), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n762_), .A2(G78gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n802_), .B1(new_n774_), .B2(new_n803_), .ZN(G1335gat));
  INV_X1    g603(.A(new_n659_), .ZN(new_n805_));
  NOR3_X1   g604(.A1(new_n610_), .A2(new_n644_), .A3(new_n805_), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n806_), .A2(new_n717_), .A3(new_n667_), .ZN(new_n807_));
  AOI21_X1  g606(.A(G85gat), .B1(new_n807_), .B2(new_n547_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n806_), .B(KEYINPUT115), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n720_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(KEYINPUT116), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n809_), .A2(new_n812_), .A3(new_n720_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n811_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n547_), .A2(G85gat), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n815_), .B(KEYINPUT117), .Z(new_n816_));
  AOI21_X1  g615(.A(new_n808_), .B1(new_n814_), .B2(new_n816_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT118), .ZN(G1336gat));
  AOI21_X1  g617(.A(G92gat), .B1(new_n807_), .B2(new_n673_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n736_), .A2(new_n251_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n819_), .B1(new_n814_), .B2(new_n820_), .ZN(G1337gat));
  NAND3_X1  g620(.A1(new_n807_), .A2(new_n261_), .A3(new_n564_), .ZN(new_n822_));
  XOR2_X1   g621(.A(new_n822_), .B(KEYINPUT119), .Z(new_n823_));
  AOI21_X1  g622(.A(new_n410_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n824_));
  OAI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(new_n211_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT51), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(KEYINPUT120), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n825_), .B(new_n827_), .ZN(G1338gat));
  NAND3_X1  g627(.A1(new_n807_), .A2(new_n212_), .A3(new_n697_), .ZN(new_n829_));
  OAI21_X1  g628(.A(G106gat), .B1(new_n810_), .B2(new_n762_), .ZN(new_n830_));
  AND2_X1   g629(.A1(new_n830_), .A2(KEYINPUT52), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(KEYINPUT52), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n829_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g633(.A(new_n565_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n736_), .A2(new_n547_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n604_), .B1(new_n641_), .B2(new_n642_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n839_), .B1(new_n595_), .B2(new_n582_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n595_), .A2(new_n582_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NOR3_X1   g641(.A1(new_n595_), .A2(new_n839_), .A3(new_n582_), .ZN(new_n843_));
  OAI211_X1 g642(.A(KEYINPUT56), .B(new_n602_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n602_), .B1(new_n842_), .B2(new_n843_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT56), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n838_), .B1(new_n844_), .B2(new_n847_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n621_), .A2(new_n623_), .A3(new_n630_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n634_), .B1(new_n629_), .B2(new_n624_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n635_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n605_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT121), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(KEYINPUT121), .A3(new_n605_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n666_), .B1(new_n848_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(KEYINPUT57), .B(new_n666_), .C1(new_n848_), .C2(new_n857_), .ZN(new_n861_));
  AND2_X1   g660(.A1(new_n860_), .A2(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n847_), .A2(KEYINPUT122), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n845_), .A2(new_n864_), .A3(new_n846_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n863_), .A2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n844_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n867_), .A2(KEYINPUT58), .A3(new_n604_), .A4(new_n852_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT58), .ZN(new_n869_));
  INV_X1    g668(.A(new_n844_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(new_n863_), .B2(new_n865_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n852_), .A2(new_n604_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n869_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n868_), .A2(new_n361_), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n805_), .B1(new_n862_), .B2(new_n874_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n710_), .A2(new_n643_), .A3(new_n610_), .A4(new_n805_), .ZN(new_n876_));
  XOR2_X1   g675(.A(new_n876_), .B(KEYINPUT54), .Z(new_n877_));
  OAI211_X1 g676(.A(new_n835_), .B(new_n837_), .C1(new_n875_), .C2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(KEYINPUT59), .ZN(new_n879_));
  AND3_X1   g678(.A1(new_n868_), .A2(new_n361_), .A3(new_n873_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n860_), .A2(new_n861_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n659_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n876_), .B(KEYINPUT54), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  XOR2_X1   g683(.A(KEYINPUT123), .B(KEYINPUT59), .Z(new_n885_));
  NAND4_X1  g684(.A1(new_n884_), .A2(new_n835_), .A3(new_n837_), .A4(new_n885_), .ZN(new_n886_));
  NAND3_X1  g685(.A1(new_n879_), .A2(new_n886_), .A3(new_n644_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(G113gat), .ZN(new_n888_));
  OR3_X1    g687(.A1(new_n878_), .A2(G113gat), .A3(new_n643_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1340gat));
  NAND3_X1  g689(.A1(new_n879_), .A2(new_n886_), .A3(new_n609_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(G120gat), .ZN(new_n892_));
  INV_X1    g691(.A(G120gat), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n893_), .A2(KEYINPUT60), .ZN(new_n894_));
  AOI21_X1  g693(.A(KEYINPUT60), .B1(new_n609_), .B2(new_n893_), .ZN(new_n895_));
  OR3_X1    g694(.A1(new_n878_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n892_), .A2(new_n896_), .ZN(G1341gat));
  NAND3_X1  g696(.A1(new_n879_), .A2(new_n886_), .A3(new_n805_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G127gat), .ZN(new_n899_));
  OR3_X1    g698(.A1(new_n878_), .A2(G127gat), .A3(new_n659_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1342gat));
  NAND3_X1  g700(.A1(new_n879_), .A2(new_n886_), .A3(new_n361_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(G134gat), .ZN(new_n903_));
  OR3_X1    g702(.A1(new_n878_), .A2(G134gat), .A3(new_n666_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(G1343gat));
  AOI21_X1  g704(.A(new_n569_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n906_), .A2(new_n644_), .A3(new_n837_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g707(.A1(new_n906_), .A2(new_n609_), .A3(new_n837_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g709(.A1(new_n906_), .A2(new_n805_), .A3(new_n837_), .ZN(new_n911_));
  XOR2_X1   g710(.A(KEYINPUT61), .B(G155gat), .Z(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT124), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n911_), .B(new_n913_), .ZN(G1346gat));
  NAND2_X1  g713(.A1(new_n906_), .A2(new_n837_), .ZN(new_n915_));
  OAI21_X1  g714(.A(G162gat), .B1(new_n915_), .B2(new_n710_), .ZN(new_n916_));
  OR2_X1    g715(.A1(new_n666_), .A2(G162gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n916_), .B1(new_n915_), .B2(new_n917_), .ZN(G1347gat));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n736_), .A2(new_n547_), .ZN(new_n920_));
  OAI211_X1 g719(.A(new_n835_), .B(new_n920_), .C1(new_n875_), .C2(new_n877_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n921_), .A2(new_n643_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n919_), .B1(new_n922_), .B2(new_n388_), .ZN(new_n923_));
  OAI211_X1 g722(.A(KEYINPUT62), .B(G169gat), .C1(new_n921_), .C2(new_n643_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n922_), .A2(new_n379_), .ZN(new_n925_));
  NAND3_X1  g724(.A1(new_n923_), .A2(new_n924_), .A3(new_n925_), .ZN(G1348gat));
  NOR2_X1   g725(.A1(new_n921_), .A2(new_n610_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n927_), .B1(KEYINPUT125), .B2(G176gat), .ZN(new_n928_));
  XOR2_X1   g727(.A(KEYINPUT125), .B(G176gat), .Z(new_n929_));
  NOR3_X1   g728(.A1(new_n921_), .A2(new_n610_), .A3(new_n929_), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n928_), .A2(new_n930_), .ZN(G1349gat));
  NOR2_X1   g730(.A1(new_n921_), .A2(new_n659_), .ZN(new_n932_));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933_));
  OAI211_X1 g732(.A(new_n932_), .B(new_n383_), .C1(new_n933_), .C2(G183gat), .ZN(new_n934_));
  NOR2_X1   g733(.A1(KEYINPUT126), .A2(G183gat), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n934_), .B1(new_n932_), .B2(new_n935_), .ZN(G1350gat));
  OAI21_X1  g735(.A(G190gat), .B1(new_n921_), .B2(new_n710_), .ZN(new_n937_));
  NAND3_X1  g736(.A1(new_n667_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n938_));
  OAI21_X1  g737(.A(new_n937_), .B1(new_n921_), .B2(new_n938_), .ZN(G1351gat));
  NAND3_X1  g738(.A1(new_n906_), .A2(new_n644_), .A3(new_n920_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g740(.A1(new_n906_), .A2(new_n609_), .A3(new_n920_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g742(.A(KEYINPUT63), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n805_), .B1(new_n944_), .B2(new_n652_), .ZN(new_n945_));
  XNOR2_X1  g744(.A(new_n945_), .B(KEYINPUT127), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n906_), .A2(new_n920_), .A3(new_n946_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n944_), .A2(new_n652_), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n947_), .B(new_n948_), .ZN(G1354gat));
  NAND2_X1  g748(.A1(new_n906_), .A2(new_n920_), .ZN(new_n950_));
  OAI21_X1  g749(.A(G218gat), .B1(new_n950_), .B2(new_n710_), .ZN(new_n951_));
  OR2_X1    g750(.A1(new_n666_), .A2(G218gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n950_), .B2(new_n952_), .ZN(G1355gat));
endmodule


