//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n760_, new_n761_, new_n762_, new_n763_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n872_, new_n873_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n906_, new_n907_, new_n909_, new_n910_, new_n912_, new_n913_,
    new_n915_, new_n916_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_;
  INV_X1    g000(.A(KEYINPUT38), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT75), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(KEYINPUT13), .ZN(new_n204_));
  OR2_X1    g003(.A1(new_n203_), .A2(KEYINPUT13), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT73), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT12), .ZN(new_n207_));
  XOR2_X1   g006(.A(KEYINPUT10), .B(G99gat), .Z(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  XOR2_X1   g009(.A(new_n210_), .B(KEYINPUT67), .Z(new_n211_));
  NOR2_X1   g010(.A1(KEYINPUT68), .A2(KEYINPUT9), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G85gat), .A3(G92gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT6), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n214_), .B1(G99gat), .B2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G99gat), .A2(G106gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(KEYINPUT68), .B(KEYINPUT9), .ZN(new_n220_));
  OAI221_X1 g019(.A(new_n213_), .B1(new_n215_), .B2(new_n217_), .C1(new_n219_), .C2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n211_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT71), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT70), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n224_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n216_), .A2(KEYINPUT6), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n214_), .A2(G99gat), .A3(G106gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n227_), .A3(KEYINPUT70), .ZN(new_n228_));
  NAND2_X1  g027(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  NOR2_X1   g029(.A1(KEYINPUT69), .A2(KEYINPUT7), .ZN(new_n231_));
  OAI22_X1  g030(.A1(new_n230_), .A2(new_n231_), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  INV_X1    g031(.A(G99gat), .ZN(new_n233_));
  INV_X1    g032(.A(G106gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n229_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  NAND4_X1  g034(.A1(new_n225_), .A2(new_n228_), .A3(new_n232_), .A4(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(new_n218_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n223_), .B1(new_n237_), .B2(KEYINPUT8), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT8), .ZN(new_n239_));
  AOI211_X1 g038(.A(KEYINPUT71), .B(new_n239_), .C1(new_n236_), .C2(new_n218_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n232_), .B(new_n235_), .C1(new_n215_), .C2(new_n217_), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n242_), .A2(new_n239_), .A3(new_n218_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n222_), .B1(new_n241_), .B2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G57gat), .B(G64gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(KEYINPUT11), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G71gat), .B(G78gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n246_), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n245_), .A2(KEYINPUT11), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n248_), .B1(new_n251_), .B2(new_n247_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n207_), .B1(new_n244_), .B2(new_n253_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G230gat), .A2(G233gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n257_), .B1(new_n244_), .B2(new_n253_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT70), .B1(new_n226_), .B2(new_n227_), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT69), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT7), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n262_), .A2(new_n229_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n235_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n259_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n219_), .B1(new_n265_), .B2(new_n228_), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT71), .B1(new_n266_), .B2(new_n239_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n237_), .A2(new_n223_), .A3(KEYINPUT8), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n267_), .A2(new_n268_), .A3(new_n243_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n222_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n253_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT12), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n254_), .A2(new_n258_), .A3(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n269_), .A2(new_n270_), .A3(new_n253_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n257_), .B1(new_n275_), .B2(new_n271_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n273_), .A2(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT5), .B(G176gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G204gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(G120gat), .B(G148gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(KEYINPUT72), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n206_), .B1(new_n277_), .B2(new_n283_), .ZN(new_n284_));
  AOI211_X1 g083(.A(KEYINPUT73), .B(new_n282_), .C1(new_n273_), .C2(new_n276_), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n257_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n269_), .A2(new_n270_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(new_n252_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n287_), .B1(new_n289_), .B2(new_n274_), .ZN(new_n290_));
  AOI21_X1  g089(.A(KEYINPUT12), .B1(new_n288_), .B2(new_n252_), .ZN(new_n291_));
  AOI211_X1 g090(.A(new_n207_), .B(new_n253_), .C1(new_n269_), .C2(new_n270_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n290_), .B1(new_n293_), .B2(new_n258_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n281_), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT74), .B1(new_n286_), .B2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT73), .B1(new_n294_), .B2(new_n282_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n277_), .A2(new_n206_), .A3(new_n283_), .ZN(new_n298_));
  AND4_X1   g097(.A1(KEYINPUT74), .A2(new_n297_), .A3(new_n295_), .A4(new_n298_), .ZN(new_n299_));
  OAI211_X1 g098(.A(new_n204_), .B(new_n205_), .C1(new_n296_), .C2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n297_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT74), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n297_), .A2(KEYINPUT74), .A3(new_n295_), .A4(new_n298_), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n303_), .A2(new_n203_), .A3(KEYINPUT13), .A4(new_n304_), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G15gat), .B(G22gat), .Z(new_n307_));
  NAND2_X1  g106(.A1(G1gat), .A2(G8gat), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n307_), .B1(KEYINPUT14), .B2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT80), .ZN(new_n310_));
  XOR2_X1   g109(.A(G1gat), .B(G8gat), .Z(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT80), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n309_), .B(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n311_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n312_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G231gat), .A2(G233gat), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n312_), .A2(new_n316_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(G231gat), .A3(G233gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n319_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n252_), .ZN(new_n323_));
  XOR2_X1   g122(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n324_));
  XNOR2_X1  g123(.A(G127gat), .B(G155gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G183gat), .B(G211gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT17), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n319_), .A2(new_n253_), .A3(new_n321_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n323_), .A2(new_n329_), .A3(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT82), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n323_), .A2(new_n330_), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT17), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n328_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT82), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n323_), .A2(new_n337_), .A3(new_n329_), .A4(new_n330_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n332_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n339_), .B(KEYINPUT83), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G232gat), .A2(G233gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT34), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G29gat), .B(G36gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(G50gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(KEYINPUT76), .B(G43gat), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n344_), .A2(new_n345_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(KEYINPUT15), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n344_), .B(new_n345_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT15), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n244_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n288_), .A2(new_n348_), .ZN(new_n355_));
  OAI211_X1 g154(.A(KEYINPUT35), .B(new_n342_), .C1(new_n354_), .C2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n353_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n288_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n244_), .A2(new_n350_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n342_), .A2(KEYINPUT35), .ZN(new_n360_));
  OR2_X1    g159(.A1(new_n342_), .A2(KEYINPUT35), .ZN(new_n361_));
  NAND4_X1  g160(.A1(new_n358_), .A2(new_n359_), .A3(new_n360_), .A4(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n356_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(G134gat), .B(G162gat), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(G218gat), .ZN(new_n365_));
  XOR2_X1   g164(.A(KEYINPUT77), .B(G190gat), .Z(new_n366_));
  XNOR2_X1  g165(.A(new_n365_), .B(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n368_), .A2(KEYINPUT36), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n368_), .A2(KEYINPUT36), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n363_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT79), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n356_), .A2(new_n369_), .A3(new_n362_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n374_), .A2(KEYINPUT78), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(KEYINPUT78), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT79), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n363_), .A2(new_n377_), .A3(new_n370_), .A4(new_n371_), .ZN(new_n378_));
  NAND4_X1  g177(.A1(new_n373_), .A2(new_n375_), .A3(new_n376_), .A4(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(KEYINPUT37), .ZN(new_n380_));
  AND3_X1   g179(.A1(new_n363_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n374_), .ZN(new_n382_));
  NOR3_X1   g181(.A1(new_n381_), .A2(KEYINPUT37), .A3(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n340_), .B1(new_n380_), .B2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n306_), .A2(new_n385_), .ZN(new_n386_));
  OR2_X1    g185(.A1(new_n386_), .A2(KEYINPUT84), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n317_), .A2(new_n348_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n320_), .A2(new_n350_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(G229gat), .A2(G233gat), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n357_), .A2(new_n317_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(new_n391_), .A3(new_n389_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n393_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G113gat), .B(G141gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(G169gat), .B(G197gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(KEYINPUT85), .A3(new_n400_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n393_), .A2(new_n395_), .A3(new_n400_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT85), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n405_), .B1(new_n396_), .B2(new_n400_), .ZN(new_n406_));
  AND2_X1   g205(.A1(new_n387_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(G1gat), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT102), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT4), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G127gat), .B(G134gat), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G113gat), .B(G120gat), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n412_), .A3(KEYINPUT92), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n411_), .A2(new_n412_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n411_), .A2(new_n412_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n413_), .B1(new_n416_), .B2(KEYINPUT92), .ZN(new_n417_));
  OR4_X1    g216(.A1(KEYINPUT93), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(G141gat), .A2(G148gat), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT2), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(G141gat), .ZN(new_n422_));
  INV_X1    g221(.A(G148gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n424_), .B1(KEYINPUT93), .B2(KEYINPUT3), .ZN(new_n425_));
  NAND3_X1  g224(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n426_));
  NAND4_X1  g225(.A1(new_n418_), .A2(new_n421_), .A3(new_n425_), .A4(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(G155gat), .A2(G162gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(G155gat), .A2(G162gat), .ZN(new_n429_));
  NOR2_X1   g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n427_), .A2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT1), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n429_), .B1(new_n428_), .B2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n433_), .B1(new_n432_), .B2(new_n428_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n434_), .A2(new_n424_), .A3(new_n419_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n431_), .A2(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n417_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n431_), .A2(new_n416_), .A3(new_n435_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n410_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT4), .B1(new_n417_), .B2(new_n436_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(G225gat), .A2(G233gat), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n409_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n437_), .A2(new_n438_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(new_n442_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n442_), .ZN(new_n446_));
  OAI211_X1 g245(.A(KEYINPUT102), .B(new_n446_), .C1(new_n439_), .C2(new_n440_), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n445_), .A3(new_n447_), .ZN(new_n448_));
  XOR2_X1   g247(.A(KEYINPUT103), .B(KEYINPUT0), .Z(new_n449_));
  XNOR2_X1  g248(.A(G1gat), .B(G29gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G57gat), .B(G85gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n448_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n453_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n443_), .A2(new_n455_), .A3(new_n445_), .A4(new_n447_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n454_), .A2(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(KEYINPUT95), .B(G204gat), .Z(new_n458_));
  NOR2_X1   g257(.A1(new_n458_), .A2(G197gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT94), .B(G197gat), .ZN(new_n460_));
  NOR2_X1   g259(.A1(new_n460_), .A2(G204gat), .ZN(new_n461_));
  OAI21_X1  g260(.A(KEYINPUT21), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  XOR2_X1   g261(.A(G211gat), .B(G218gat), .Z(new_n463_));
  INV_X1    g262(.A(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT96), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n458_), .A2(new_n465_), .A3(G197gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n460_), .A2(G204gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT95), .B(G204gat), .ZN(new_n468_));
  INV_X1    g267(.A(G197gat), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT96), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n466_), .A2(new_n467_), .A3(new_n470_), .ZN(new_n471_));
  OAI211_X1 g270(.A(new_n462_), .B(new_n464_), .C1(new_n471_), .C2(KEYINPUT21), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n471_), .A2(KEYINPUT21), .A3(new_n463_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n436_), .A2(KEYINPUT29), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G228gat), .A2(G233gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G50gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT28), .B1(new_n436_), .B2(KEYINPUT29), .ZN(new_n480_));
  INV_X1    g279(.A(G22gat), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT28), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT29), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n431_), .A2(new_n435_), .A3(new_n482_), .A4(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n480_), .A2(new_n481_), .A3(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n481_), .B1(new_n480_), .B2(new_n484_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n479_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n487_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(G50gat), .A3(new_n485_), .ZN(new_n490_));
  XOR2_X1   g289(.A(G78gat), .B(G106gat), .Z(new_n491_));
  OR2_X1    g290(.A1(new_n491_), .A2(KEYINPUT97), .ZN(new_n492_));
  AND3_X1   g291(.A1(new_n488_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n491_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n478_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n478_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n488_), .A2(new_n490_), .A3(new_n492_), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n488_), .A2(new_n490_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n496_), .B(new_n497_), .C1(new_n498_), .C2(new_n491_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G8gat), .B(G36gat), .ZN(new_n501_));
  INV_X1    g300(.A(G92gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  XNOR2_X1  g302(.A(KEYINPUT18), .B(G64gat), .ZN(new_n504_));
  XOR2_X1   g303(.A(new_n503_), .B(new_n504_), .Z(new_n505_));
  NAND2_X1  g304(.A1(G226gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT19), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT100), .ZN(new_n508_));
  XNOR2_X1  g307(.A(KEYINPUT90), .B(G176gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(KEYINPUT22), .B(G169gat), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G183gat), .A2(G190gat), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT23), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n515_), .B(new_n516_), .C1(G183gat), .C2(G190gat), .ZN(new_n517_));
  INV_X1    g316(.A(G169gat), .ZN(new_n518_));
  INV_X1    g317(.A(G176gat), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n517_), .A2(new_n521_), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n508_), .B1(new_n512_), .B2(new_n522_), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n510_), .A2(new_n511_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n524_), .A2(new_n517_), .A3(KEYINPUT100), .A4(new_n521_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT24), .ZN(new_n527_));
  NOR2_X1   g326(.A1(G169gat), .A2(G176gat), .ZN(new_n528_));
  NOR3_X1   g327(.A1(new_n520_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT25), .B(G183gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(KEYINPUT26), .B(G190gat), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n529_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n527_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n533_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n534_), .A2(KEYINPUT98), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n534_), .A2(KEYINPUT98), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n532_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT99), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n534_), .B(KEYINPUT98), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT99), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n539_), .A2(new_n540_), .A3(new_n532_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n526_), .B1(new_n538_), .B2(new_n541_), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n472_), .A2(new_n473_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n507_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT26), .ZN(new_n545_));
  OAI21_X1  g344(.A(KEYINPUT87), .B1(new_n545_), .B2(G190gat), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT87), .ZN(new_n547_));
  INV_X1    g346(.A(G190gat), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n547_), .A2(new_n548_), .A3(KEYINPUT26), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT25), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n546_), .A2(new_n549_), .B1(new_n550_), .B2(G183gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n545_), .A2(G190gat), .ZN(new_n552_));
  OAI21_X1  g351(.A(KEYINPUT86), .B1(new_n550_), .B2(G183gat), .ZN(new_n553_));
  OR3_X1    g352(.A1(new_n550_), .A2(KEYINPUT86), .A3(G183gat), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n551_), .A2(new_n552_), .A3(new_n553_), .A4(new_n554_), .ZN(new_n555_));
  OR2_X1    g354(.A1(new_n534_), .A2(KEYINPUT88), .ZN(new_n556_));
  INV_X1    g355(.A(new_n529_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n534_), .A2(KEYINPUT88), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n555_), .A2(new_n556_), .A3(new_n557_), .A4(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n560_));
  OAI21_X1  g359(.A(KEYINPUT22), .B1(new_n518_), .B2(KEYINPUT89), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n518_), .A2(KEYINPUT22), .ZN(new_n562_));
  OAI211_X1 g361(.A(new_n510_), .B(new_n561_), .C1(KEYINPUT89), .C2(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n563_), .A2(new_n521_), .A3(new_n517_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n559_), .A2(new_n560_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n560_), .B1(new_n559_), .B2(new_n564_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n474_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n544_), .A2(KEYINPUT20), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n507_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT20), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n523_), .A2(new_n525_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n541_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n540_), .B1(new_n539_), .B2(new_n532_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n571_), .B1(new_n575_), .B2(new_n474_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n559_), .A2(new_n564_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n577_), .A2(KEYINPUT91), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n543_), .A2(new_n578_), .A3(new_n565_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n570_), .B1(new_n576_), .B2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n505_), .B1(new_n569_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n579_), .ZN(new_n582_));
  OAI21_X1  g381(.A(KEYINPUT20), .B1(new_n542_), .B2(new_n543_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n507_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n505_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n578_), .A2(new_n565_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n571_), .B1(new_n586_), .B2(new_n474_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n544_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n584_), .A2(new_n585_), .A3(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n581_), .A2(KEYINPUT101), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT27), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT101), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n592_), .B(new_n505_), .C1(new_n569_), .C2(new_n580_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n590_), .A2(new_n591_), .A3(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n457_), .ZN(new_n595_));
  NOR3_X1   g394(.A1(new_n582_), .A2(new_n583_), .A3(new_n507_), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n543_), .B(new_n537_), .C1(new_n522_), .C2(new_n512_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n570_), .B1(new_n587_), .B2(new_n597_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n505_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(KEYINPUT27), .A3(new_n589_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n500_), .A2(new_n594_), .A3(new_n595_), .A4(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n444_), .A2(new_n446_), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n453_), .B(new_n602_), .C1(new_n441_), .C2(new_n446_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n604_), .B1(new_n590_), .B2(new_n593_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n456_), .B(KEYINPUT33), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n596_), .A2(new_n598_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n585_), .A2(KEYINPUT32), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  AOI22_X1  g408(.A1(new_n607_), .A2(new_n609_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n584_), .A2(new_n608_), .A3(new_n588_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT104), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  AOI22_X1  g412(.A1(new_n605_), .A2(new_n606_), .B1(new_n610_), .B2(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n601_), .B1(new_n614_), .B2(new_n500_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G227gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(KEYINPUT31), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n417_), .B(new_n617_), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n586_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G71gat), .B(G99gat), .ZN(new_n620_));
  INV_X1    g419(.A(G43gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XOR2_X1   g421(.A(KEYINPUT30), .B(G15gat), .Z(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(new_n619_), .B(new_n624_), .Z(new_n625_));
  NAND2_X1  g424(.A1(new_n495_), .A2(new_n499_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n594_), .A2(new_n626_), .A3(new_n600_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT105), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n594_), .A2(KEYINPUT105), .A3(new_n626_), .A4(new_n600_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n625_), .A2(new_n457_), .ZN(new_n632_));
  AOI22_X1  g431(.A1(new_n615_), .A2(new_n625_), .B1(new_n631_), .B2(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n386_), .B2(KEYINPUT84), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n407_), .A2(new_n408_), .A3(new_n457_), .A4(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT106), .ZN(new_n636_));
  INV_X1    g435(.A(new_n636_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n635_), .A2(KEYINPUT106), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n202_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  OR2_X1    g438(.A1(new_n635_), .A2(KEYINPUT106), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n640_), .A2(KEYINPUT38), .A3(new_n636_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n300_), .A2(new_n305_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n406_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n381_), .A2(KEYINPUT107), .A3(new_n382_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT107), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n646_), .B1(new_n372_), .B2(new_n374_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n645_), .A2(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n631_), .A2(new_n632_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n605_), .A2(new_n606_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n610_), .A2(new_n613_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n500_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n601_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n625_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n650_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n339_), .ZN(new_n657_));
  NAND4_X1  g456(.A1(new_n644_), .A2(new_n649_), .A3(new_n656_), .A4(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G1gat), .B1(new_n658_), .B2(new_n595_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n639_), .A2(new_n641_), .A3(new_n659_), .ZN(G1324gat));
  NAND2_X1  g459(.A1(new_n594_), .A2(new_n600_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n662_), .A2(G8gat), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n387_), .A2(new_n634_), .A3(new_n406_), .A4(new_n663_), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n664_), .B(KEYINPUT108), .ZN(new_n665_));
  INV_X1    g464(.A(G8gat), .ZN(new_n666_));
  INV_X1    g465(.A(new_n658_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n667_), .B2(new_n661_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT39), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n668_), .A2(new_n669_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n665_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(new_n665_), .B(KEYINPUT40), .C1(new_n670_), .C2(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1325gat));
  AND2_X1   g475(.A1(new_n407_), .A2(new_n634_), .ZN(new_n677_));
  INV_X1    g476(.A(G15gat), .ZN(new_n678_));
  INV_X1    g477(.A(new_n625_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G15gat), .B1(new_n658_), .B2(new_n625_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT41), .Z(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(G1326gat));
  NAND3_X1  g482(.A1(new_n677_), .A2(new_n481_), .A3(new_n500_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G22gat), .B1(new_n658_), .B2(new_n626_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT42), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1327gat));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n306_), .A2(new_n406_), .A3(new_n340_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n383_), .B1(new_n379_), .B2(KEYINPUT37), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT43), .B1(new_n633_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT43), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n656_), .A2(new_n693_), .A3(new_n690_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n689_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n688_), .B1(new_n695_), .B2(KEYINPUT109), .ZN(new_n696_));
  INV_X1    g495(.A(new_n340_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n642_), .A2(new_n643_), .A3(new_n697_), .ZN(new_n698_));
  NOR3_X1   g497(.A1(new_n633_), .A2(KEYINPUT43), .A3(new_n691_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n693_), .B1(new_n656_), .B2(new_n690_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT109), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n701_), .A2(new_n702_), .A3(KEYINPUT44), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n696_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G29gat), .B1(new_n704_), .B2(new_n595_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n633_), .A2(new_n649_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n698_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(G29gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n707_), .A2(new_n708_), .A3(new_n457_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n705_), .A2(new_n709_), .ZN(G1328gat));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT112), .ZN(new_n712_));
  INV_X1    g511(.A(G36gat), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n698_), .A2(new_n706_), .A3(new_n713_), .A4(new_n661_), .ZN(new_n714_));
  XOR2_X1   g513(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT110), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n714_), .B(new_n716_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n662_), .B1(new_n696_), .B2(new_n703_), .ZN(new_n718_));
  OAI211_X1 g517(.A(new_n712_), .B(new_n717_), .C1(new_n718_), .C2(new_n713_), .ZN(new_n719_));
  OR2_X1    g518(.A1(new_n711_), .A2(KEYINPUT112), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n719_), .B(new_n720_), .ZN(G1329gat));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722_));
  OAI21_X1  g521(.A(G43gat), .B1(new_n704_), .B2(new_n625_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n707_), .A2(new_n621_), .A3(new_n679_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n625_), .B1(new_n696_), .B2(new_n703_), .ZN(new_n726_));
  OAI211_X1 g525(.A(new_n722_), .B(new_n724_), .C1(new_n726_), .C2(new_n621_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n727_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n725_), .A2(new_n728_), .ZN(G1330gat));
  OAI21_X1  g528(.A(G50gat), .B1(new_n704_), .B2(new_n626_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n707_), .A2(new_n479_), .A3(new_n500_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1331gat));
  NOR3_X1   g531(.A1(new_n306_), .A2(new_n633_), .A3(new_n406_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(new_n385_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(G57gat), .B1(new_n736_), .B2(new_n457_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n733_), .A2(new_n649_), .A3(new_n697_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n738_), .A2(new_n595_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n737_), .B1(G57gat), .B2(new_n739_), .ZN(G1332gat));
  INV_X1    g539(.A(G64gat), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n736_), .A2(new_n741_), .A3(new_n661_), .ZN(new_n742_));
  OR2_X1    g541(.A1(new_n738_), .A2(new_n662_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT48), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(G64gat), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n744_), .B1(new_n743_), .B2(G64gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n742_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT114), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(new_n749_), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n742_), .B(KEYINPUT114), .C1(new_n746_), .C2(new_n747_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(G1333gat));
  OAI21_X1  g551(.A(G71gat), .B1(new_n738_), .B2(new_n625_), .ZN(new_n753_));
  XOR2_X1   g552(.A(KEYINPUT115), .B(KEYINPUT49), .Z(new_n754_));
  XNOR2_X1  g553(.A(new_n753_), .B(new_n754_), .ZN(new_n755_));
  NOR2_X1   g554(.A1(new_n625_), .A2(G71gat), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT116), .Z(new_n757_));
  NAND2_X1  g556(.A1(new_n736_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n755_), .A2(new_n758_), .ZN(G1334gat));
  OAI21_X1  g558(.A(G78gat), .B1(new_n738_), .B2(new_n626_), .ZN(new_n760_));
  XNOR2_X1  g559(.A(new_n760_), .B(KEYINPUT50), .ZN(new_n761_));
  INV_X1    g560(.A(G78gat), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n736_), .A2(new_n762_), .A3(new_n500_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(G1335gat));
  NOR3_X1   g563(.A1(new_n306_), .A2(new_n406_), .A3(new_n697_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n765_), .A2(new_n706_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n766_), .ZN(new_n767_));
  AOI21_X1  g566(.A(G85gat), .B1(new_n767_), .B2(new_n457_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n692_), .A2(new_n694_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n765_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT117), .Z(new_n771_));
  NAND2_X1  g570(.A1(new_n457_), .A2(G85gat), .ZN(new_n772_));
  XOR2_X1   g571(.A(new_n772_), .B(KEYINPUT118), .Z(new_n773_));
  AOI21_X1  g572(.A(new_n768_), .B1(new_n771_), .B2(new_n773_), .ZN(G1336gat));
  NAND3_X1  g573(.A1(new_n767_), .A2(new_n502_), .A3(new_n661_), .ZN(new_n775_));
  AND2_X1   g574(.A1(new_n771_), .A2(new_n661_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(new_n502_), .ZN(G1337gat));
  OAI21_X1  g576(.A(G99gat), .B1(new_n770_), .B2(new_n625_), .ZN(new_n778_));
  AND3_X1   g577(.A1(new_n765_), .A2(new_n208_), .A3(new_n706_), .ZN(new_n779_));
  AND3_X1   g578(.A1(new_n779_), .A2(KEYINPUT119), .A3(new_n679_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT119), .B1(new_n779_), .B2(new_n679_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n778_), .B1(new_n780_), .B2(new_n781_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n782_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g582(.A1(new_n767_), .A2(new_n209_), .A3(new_n500_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n769_), .A2(new_n500_), .A3(new_n765_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n785_), .A2(new_n786_), .A3(G106gat), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n785_), .B2(G106gat), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n784_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n789_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g589(.A1(new_n631_), .A2(new_n457_), .A3(new_n679_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n293_), .A2(KEYINPUT55), .A3(new_n258_), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n273_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n254_), .A2(new_n272_), .A3(new_n274_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n257_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n792_), .A2(new_n794_), .A3(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(new_n283_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n798_), .A2(KEYINPUT56), .B1(new_n294_), .B2(new_n281_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n390_), .A2(new_n391_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n394_), .A2(new_n392_), .A3(new_n389_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n800_), .A2(new_n801_), .A3(new_n399_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n803_), .B1(new_n401_), .B2(new_n404_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n797_), .A2(new_n805_), .A3(new_n283_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n799_), .A2(new_n804_), .A3(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT58), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n799_), .A2(KEYINPUT58), .A3(new_n804_), .A4(new_n806_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n690_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT57), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n804_), .B1(new_n296_), .B2(new_n299_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n799_), .A2(new_n406_), .A3(new_n806_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n812_), .B1(new_n815_), .B2(new_n649_), .ZN(new_n816_));
  AOI211_X1 g615(.A(KEYINPUT57), .B(new_n648_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n811_), .B1(new_n816_), .B2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n339_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT54), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n306_), .A2(new_n820_), .A3(new_n643_), .A4(new_n385_), .ZN(new_n821_));
  NAND4_X1  g620(.A1(new_n385_), .A2(new_n643_), .A3(new_n300_), .A4(new_n305_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(KEYINPUT54), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n791_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(G113gat), .B1(new_n825_), .B2(new_n406_), .ZN(new_n826_));
  AOI22_X1  g625(.A1(new_n818_), .A2(new_n340_), .B1(new_n823_), .B2(new_n821_), .ZN(new_n827_));
  NOR3_X1   g626(.A1(new_n827_), .A2(KEYINPUT59), .A3(new_n791_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT59), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n825_), .B2(new_n830_), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n809_), .A2(new_n690_), .A3(new_n810_), .ZN(new_n832_));
  AND3_X1   g631(.A1(new_n799_), .A2(new_n406_), .A3(new_n806_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n804_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n649_), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(KEYINPUT57), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n815_), .A2(new_n812_), .A3(new_n649_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n832_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n824_), .B1(new_n839_), .B2(new_n657_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n791_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n842_), .A2(KEYINPUT120), .A3(KEYINPUT59), .ZN(new_n843_));
  AOI211_X1 g642(.A(new_n643_), .B(new_n828_), .C1(new_n831_), .C2(new_n843_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n826_), .B1(new_n844_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g644(.A(G120gat), .ZN(new_n846_));
  OAI21_X1  g645(.A(new_n846_), .B1(new_n306_), .B2(KEYINPUT60), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n825_), .B(new_n847_), .C1(KEYINPUT60), .C2(new_n846_), .ZN(new_n848_));
  AOI211_X1 g647(.A(new_n306_), .B(new_n828_), .C1(new_n831_), .C2(new_n843_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n846_), .ZN(G1341gat));
  AOI21_X1  g649(.A(G127gat), .B1(new_n825_), .B2(new_n697_), .ZN(new_n851_));
  INV_X1    g650(.A(G127gat), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n852_), .B(new_n828_), .C1(new_n831_), .C2(new_n843_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n853_), .B2(new_n657_), .ZN(G1342gat));
  AOI21_X1  g653(.A(G134gat), .B1(new_n825_), .B2(new_n648_), .ZN(new_n855_));
  INV_X1    g654(.A(G134gat), .ZN(new_n856_));
  AOI211_X1 g655(.A(new_n856_), .B(new_n828_), .C1(new_n831_), .C2(new_n843_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n855_), .B1(new_n857_), .B2(new_n690_), .ZN(G1343gat));
  AOI21_X1  g657(.A(new_n679_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n859_));
  NOR3_X1   g658(.A1(new_n661_), .A2(new_n595_), .A3(new_n626_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n861_), .A2(new_n643_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(KEYINPUT121), .B(G141gat), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1344gat));
  OAI21_X1  g663(.A(KEYINPUT123), .B1(new_n861_), .B2(new_n306_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT123), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n859_), .A2(new_n866_), .A3(new_n642_), .A4(new_n860_), .ZN(new_n867_));
  XNOR2_X1  g666(.A(KEYINPUT122), .B(G148gat), .ZN(new_n868_));
  AND3_X1   g667(.A1(new_n865_), .A2(new_n867_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n868_), .B1(new_n865_), .B2(new_n867_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n869_), .A2(new_n870_), .ZN(G1345gat));
  NOR2_X1   g670(.A1(new_n861_), .A2(new_n340_), .ZN(new_n872_));
  XOR2_X1   g671(.A(KEYINPUT61), .B(G155gat), .Z(new_n873_));
  XNOR2_X1  g672(.A(new_n872_), .B(new_n873_), .ZN(G1346gat));
  INV_X1    g673(.A(G162gat), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n861_), .A2(new_n875_), .A3(new_n691_), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n861_), .B2(new_n649_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n877_), .A2(new_n878_), .ZN(new_n879_));
  OAI211_X1 g678(.A(KEYINPUT124), .B(new_n875_), .C1(new_n861_), .C2(new_n649_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n876_), .B1(new_n879_), .B2(new_n880_), .ZN(G1347gat));
  NOR2_X1   g680(.A1(new_n662_), .A2(new_n457_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(new_n626_), .A3(new_n679_), .ZN(new_n883_));
  OAI21_X1  g682(.A(KEYINPUT125), .B1(new_n827_), .B2(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT125), .ZN(new_n885_));
  INV_X1    g684(.A(new_n883_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n839_), .A2(new_n697_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n821_), .A2(new_n823_), .ZN(new_n888_));
  OAI211_X1 g687(.A(new_n885_), .B(new_n886_), .C1(new_n887_), .C2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n884_), .A2(new_n889_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n890_), .A2(new_n406_), .A3(new_n511_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n406_), .B(new_n886_), .C1(new_n887_), .C2(new_n888_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893_));
  AND3_X1   g692(.A1(new_n892_), .A2(new_n893_), .A3(G169gat), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n892_), .B2(G169gat), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n891_), .B1(new_n894_), .B2(new_n895_), .ZN(G1348gat));
  INV_X1    g695(.A(KEYINPUT126), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n509_), .B1(new_n890_), .B2(new_n642_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n883_), .B1(new_n819_), .B2(new_n824_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(G176gat), .A3(new_n642_), .ZN(new_n900_));
  INV_X1    g699(.A(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n897_), .B1(new_n898_), .B2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n306_), .B1(new_n884_), .B2(new_n889_), .ZN(new_n903_));
  OAI211_X1 g702(.A(KEYINPUT126), .B(new_n900_), .C1(new_n903_), .C2(new_n509_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n902_), .A2(new_n904_), .ZN(G1349gat));
  AOI21_X1  g704(.A(G183gat), .B1(new_n899_), .B2(new_n697_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n339_), .A2(new_n530_), .ZN(new_n907_));
  AOI21_X1  g706(.A(new_n906_), .B1(new_n890_), .B2(new_n907_), .ZN(G1350gat));
  NAND3_X1  g707(.A1(new_n890_), .A2(new_n648_), .A3(new_n531_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n691_), .B1(new_n884_), .B2(new_n889_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n548_), .ZN(G1351gat));
  NAND3_X1  g710(.A1(new_n859_), .A2(new_n500_), .A3(new_n882_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n643_), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n913_), .B(new_n469_), .ZN(G1352gat));
  INV_X1    g713(.A(new_n912_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n642_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(G204gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n917_), .B1(new_n916_), .B2(new_n468_), .ZN(G1353gat));
  NOR2_X1   g717(.A1(new_n912_), .A2(new_n339_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n920_));
  AND2_X1   g719(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n919_), .B1(new_n920_), .B2(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n922_), .B1(new_n919_), .B2(new_n920_), .ZN(G1354gat));
  XOR2_X1   g722(.A(KEYINPUT127), .B(G218gat), .Z(new_n924_));
  NOR3_X1   g723(.A1(new_n912_), .A2(new_n691_), .A3(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n915_), .A2(new_n648_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(new_n924_), .ZN(G1355gat));
endmodule


