//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n878_, new_n879_, new_n880_, new_n882_,
    new_n883_, new_n885_, new_n886_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n927_, new_n928_, new_n930_, new_n932_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_;
  XOR2_X1   g000(.A(KEYINPUT93), .B(KEYINPUT18), .Z(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT94), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G8gat), .B(G36gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G64gat), .B(G92gat), .ZN(new_n206_));
  XOR2_X1   g005(.A(new_n205_), .B(new_n206_), .Z(new_n207_));
  INV_X1    g006(.A(KEYINPUT81), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT26), .B(G190gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT80), .B(G183gat), .ZN(new_n210_));
  AND2_X1   g009(.A1(new_n210_), .A2(KEYINPUT25), .ZN(new_n211_));
  NOR2_X1   g010(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n208_), .B(new_n209_), .C1(new_n211_), .C2(new_n212_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n212_), .B1(new_n210_), .B2(KEYINPUT25), .ZN(new_n214_));
  INV_X1    g013(.A(new_n209_), .ZN(new_n215_));
  OAI21_X1  g014(.A(KEYINPUT81), .B1(new_n214_), .B2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217_));
  XNOR2_X1  g016(.A(new_n217_), .B(KEYINPUT82), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n220_));
  INV_X1    g019(.A(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n219_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G183gat), .A2(G190gat), .ZN(new_n223_));
  XOR2_X1   g022(.A(new_n223_), .B(KEYINPUT23), .Z(new_n224_));
  NOR3_X1   g023(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  NAND4_X1  g025(.A1(new_n213_), .A2(new_n216_), .A3(new_n222_), .A4(new_n226_), .ZN(new_n227_));
  XOR2_X1   g026(.A(KEYINPUT84), .B(G176gat), .Z(new_n228_));
  INV_X1    g027(.A(G169gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(KEYINPUT83), .A3(KEYINPUT22), .ZN(new_n230_));
  AND2_X1   g029(.A1(KEYINPUT83), .A2(KEYINPUT22), .ZN(new_n231_));
  OAI211_X1 g030(.A(new_n228_), .B(new_n230_), .C1(new_n229_), .C2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT85), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n233_), .B1(new_n223_), .B2(KEYINPUT23), .ZN(new_n234_));
  XNOR2_X1  g033(.A(new_n223_), .B(KEYINPUT23), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n234_), .B1(new_n235_), .B2(new_n233_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n210_), .A2(G190gat), .ZN(new_n237_));
  OAI211_X1 g036(.A(new_n232_), .B(new_n219_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n227_), .A2(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(G197gat), .B(G204gat), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT21), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G197gat), .B(G204gat), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT21), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G211gat), .B(G218gat), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n241_), .A2(new_n244_), .A3(new_n245_), .ZN(new_n246_));
  OR3_X1    g045(.A1(new_n242_), .A2(new_n245_), .A3(new_n243_), .ZN(new_n247_));
  AND2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n239_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n251_));
  NAND2_X1  g050(.A1(G226gat), .A2(G233gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(new_n251_), .B(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT20), .ZN(new_n254_));
  OR2_X1    g053(.A1(G183gat), .A2(G190gat), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n219_), .A2(KEYINPUT92), .B1(new_n235_), .B2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT92), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT22), .B(G169gat), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n218_), .A2(new_n257_), .B1(new_n228_), .B2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n234_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(new_n224_), .B2(KEYINPUT85), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n225_), .B1(new_n221_), .B2(new_n217_), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT25), .B(G183gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n209_), .A2(new_n263_), .ZN(new_n264_));
  AND2_X1   g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  AOI22_X1  g064(.A1(new_n256_), .A2(new_n259_), .B1(new_n261_), .B2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n254_), .B1(new_n266_), .B2(new_n248_), .ZN(new_n267_));
  AND3_X1   g066(.A1(new_n250_), .A2(new_n253_), .A3(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n256_), .A2(new_n259_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n261_), .A2(new_n265_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n254_), .B1(new_n271_), .B2(new_n249_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n227_), .A2(new_n248_), .A3(new_n238_), .ZN(new_n273_));
  AOI21_X1  g072(.A(new_n253_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n207_), .B1(new_n268_), .B2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n273_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n253_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n205_), .B(new_n206_), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n250_), .A2(new_n253_), .A3(new_n267_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n275_), .A2(new_n281_), .A3(KEYINPUT95), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT27), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT95), .ZN(new_n284_));
  NAND4_X1  g083(.A1(new_n278_), .A2(new_n284_), .A3(new_n279_), .A4(new_n280_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n282_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n272_), .A2(new_n253_), .A3(new_n273_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n250_), .A2(new_n267_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n287_), .B1(new_n288_), .B2(new_n253_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(new_n207_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n290_), .A2(KEYINPUT27), .A3(new_n281_), .ZN(new_n291_));
  AND2_X1   g090(.A1(new_n286_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G155gat), .B(G162gat), .ZN(new_n293_));
  OR2_X1    g092(.A1(new_n293_), .A2(KEYINPUT88), .ZN(new_n294_));
  OR3_X1    g093(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(G141gat), .A2(G148gat), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT2), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n295_), .A2(new_n298_), .A3(new_n299_), .A4(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n293_), .A2(KEYINPUT88), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n294_), .A2(new_n301_), .A3(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(G141gat), .A2(G148gat), .ZN(new_n304_));
  INV_X1    g103(.A(G155gat), .ZN(new_n305_));
  INV_X1    g104(.A(G162gat), .ZN(new_n306_));
  OAI21_X1  g105(.A(KEYINPUT1), .B1(new_n305_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n307_), .B1(G155gat), .B2(G162gat), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n305_), .A2(new_n306_), .A3(KEYINPUT1), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n296_), .B(new_n304_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n303_), .A2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(G127gat), .B(G134gat), .Z(new_n312_));
  XOR2_X1   g111(.A(G113gat), .B(G120gat), .Z(new_n313_));
  XOR2_X1   g112(.A(new_n312_), .B(new_n313_), .Z(new_n314_));
  NAND2_X1  g113(.A1(new_n311_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT96), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n312_), .B(new_n313_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n317_), .A2(new_n303_), .A3(new_n310_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n315_), .A2(new_n316_), .A3(new_n318_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n317_), .A2(KEYINPUT96), .A3(new_n303_), .A4(new_n310_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n320_), .A3(KEYINPUT4), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n315_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G225gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT97), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n319_), .A2(new_n320_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n328_), .A2(new_n325_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G1gat), .B(G29gat), .Z(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT98), .B(G85gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n330_), .B(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT0), .B(G57gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n327_), .A2(new_n329_), .A3(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n334_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n329_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n326_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n338_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n336_), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT99), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n335_), .A2(new_n340_), .A3(new_n341_), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n327_), .A2(KEYINPUT99), .A3(new_n329_), .A4(new_n334_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT100), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n342_), .A2(KEYINPUT100), .A3(new_n343_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n292_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT29), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n349_), .B1(new_n303_), .B2(new_n310_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(new_n248_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(KEYINPUT89), .A2(G233gat), .ZN(new_n354_));
  OAI21_X1  g153(.A(G228gat), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n355_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n357_), .B1(new_n350_), .B2(new_n248_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G78gat), .B(G106gat), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n356_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT90), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(new_n311_), .A2(KEYINPUT29), .ZN(new_n364_));
  XNOR2_X1  g163(.A(G22gat), .B(G50gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n365_), .B(KEYINPUT28), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n364_), .B(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n363_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n356_), .A2(new_n358_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n359_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n370_), .A2(new_n361_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  NAND4_X1  g171(.A1(new_n370_), .A2(new_n367_), .A3(KEYINPUT90), .A4(new_n361_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G15gat), .B(G43gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n375_), .B(KEYINPUT86), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT30), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G227gat), .A2(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(G71gat), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G99gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n227_), .A2(new_n238_), .A3(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n384_), .B1(new_n227_), .B2(new_n238_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n378_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT31), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n239_), .A2(new_n383_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n390_), .A2(new_n377_), .A3(new_n385_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n388_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n389_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n317_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n394_));
  NOR3_X1   g193(.A1(new_n386_), .A2(new_n387_), .A3(new_n378_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n377_), .B1(new_n390_), .B2(new_n385_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT31), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n388_), .A2(new_n389_), .A3(new_n391_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(new_n314_), .A3(new_n398_), .ZN(new_n399_));
  AND3_X1   g198(.A1(new_n394_), .A2(KEYINPUT87), .A3(new_n399_), .ZN(new_n400_));
  AOI21_X1  g199(.A(KEYINPUT87), .B1(new_n394_), .B2(new_n399_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n374_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n374_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n392_), .A2(new_n393_), .A3(new_n317_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n314_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n403_), .A2(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n402_), .A2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT33), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n335_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n282_), .A2(new_n285_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n324_), .A2(new_n325_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n334_), .B1(new_n328_), .B2(new_n326_), .ZN(new_n413_));
  AOI22_X1  g212(.A1(new_n335_), .A2(new_n409_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n410_), .A2(new_n411_), .A3(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n279_), .A2(KEYINPUT32), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(new_n274_), .B2(new_n268_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n417_), .B1(new_n289_), .B2(new_n416_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n342_), .A2(new_n418_), .A3(new_n343_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n415_), .A2(new_n419_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT87), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n421_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n394_), .A2(KEYINPUT87), .A3(new_n399_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n374_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  AOI22_X1  g223(.A1(new_n348_), .A2(new_n408_), .B1(new_n420_), .B2(new_n424_), .ZN(new_n425_));
  XOR2_X1   g224(.A(G29gat), .B(G36gat), .Z(new_n426_));
  XOR2_X1   g225(.A(G43gat), .B(G50gat), .Z(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G29gat), .B(G36gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G43gat), .B(G50gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n428_), .A2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT15), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  AOI21_X1  g233(.A(KEYINPUT15), .B1(new_n428_), .B2(new_n431_), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G15gat), .B(G22gat), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G1gat), .A2(G8gat), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT14), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(G1gat), .ZN(new_n441_));
  INV_X1    g240(.A(G8gat), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n443_), .A2(new_n438_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n440_), .A2(new_n444_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n437_), .A2(new_n438_), .A3(new_n443_), .A4(new_n439_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n436_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n432_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G229gat), .A2(G233gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n448_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n447_), .A2(new_n431_), .A3(new_n428_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n449_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n450_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n451_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G113gat), .B(G141gat), .Z(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT79), .ZN(new_n458_));
  XNOR2_X1  g257(.A(G169gat), .B(G197gat), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n456_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n460_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n451_), .A2(new_n455_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n461_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n425_), .A2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(G230gat), .A2(G233gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT64), .ZN(new_n468_));
  OR2_X1    g267(.A1(G85gat), .A2(G92gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G85gat), .A2(G92gat), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G99gat), .A2(G106gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(KEYINPUT6), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT6), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n474_), .A2(G99gat), .A3(G106gat), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT7), .ZN(new_n477_));
  INV_X1    g276(.A(G106gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n382_), .A3(new_n478_), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n471_), .B1(new_n476_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(KEYINPUT66), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n474_), .B1(G99gat), .B2(G106gat), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n472_), .A2(KEYINPUT6), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n480_), .B(new_n479_), .C1(new_n484_), .C2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT66), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n486_), .A2(new_n487_), .A3(new_n471_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n483_), .A2(KEYINPUT8), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n473_), .A2(new_n475_), .ZN(new_n490_));
  INV_X1    g289(.A(G85gat), .ZN(new_n491_));
  NOR2_X1   g290(.A1(new_n491_), .A2(KEYINPUT9), .ZN(new_n492_));
  AND2_X1   g291(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n492_), .B1(new_n493_), .B2(new_n494_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n469_), .A2(KEYINPUT9), .A3(new_n470_), .ZN(new_n496_));
  OR2_X1    g295(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n497_), .A2(new_n478_), .A3(new_n498_), .ZN(new_n499_));
  AND4_X1   g298(.A1(new_n490_), .A2(new_n495_), .A3(new_n496_), .A4(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n487_), .B1(new_n486_), .B2(new_n471_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT8), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n500_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n380_), .A2(KEYINPUT67), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT67), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(G71gat), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n504_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(G78gat), .ZN(new_n508_));
  INV_X1    g307(.A(G78gat), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n504_), .A2(new_n506_), .A3(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(G64gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(G57gat), .ZN(new_n512_));
  INV_X1    g311(.A(G57gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(G64gat), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n514_), .A3(KEYINPUT11), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT11), .B1(new_n512_), .B2(new_n514_), .ZN(new_n517_));
  OAI211_X1 g316(.A(new_n508_), .B(new_n510_), .C1(new_n516_), .C2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n510_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n509_), .B1(new_n504_), .B2(new_n506_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n515_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  AND2_X1   g320(.A1(new_n518_), .A2(new_n521_), .ZN(new_n522_));
  AND3_X1   g321(.A1(new_n489_), .A2(new_n503_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n522_), .B1(new_n489_), .B2(new_n503_), .ZN(new_n524_));
  OAI21_X1  g323(.A(new_n468_), .B1(new_n523_), .B2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT68), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(KEYINPUT68), .B(new_n468_), .C1(new_n523_), .C2(new_n524_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n522_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n486_), .A2(new_n487_), .A3(new_n471_), .ZN(new_n531_));
  NOR3_X1   g330(.A1(new_n531_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n482_), .A2(KEYINPUT66), .A3(new_n502_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n500_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n530_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n489_), .A2(new_n503_), .A3(new_n522_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(KEYINPUT12), .A3(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT12), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n524_), .A2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n538_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n468_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G120gat), .B(G148gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT70), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G176gat), .B(G204gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n545_), .B(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n529_), .A2(new_n543_), .A3(new_n549_), .ZN(new_n550_));
  AOI22_X1  g349(.A1(new_n527_), .A2(new_n528_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n549_), .B(KEYINPUT71), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n550_), .B(KEYINPUT72), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n529_), .A2(new_n543_), .ZN(new_n554_));
  XOR2_X1   g353(.A(new_n549_), .B(KEYINPUT71), .Z(new_n555_));
  INV_X1    g354(.A(KEYINPUT72), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n554_), .A2(new_n555_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n553_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n559_));
  NOR2_X1   g358(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n558_), .A2(new_n559_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT73), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT13), .ZN(new_n564_));
  NAND4_X1  g363(.A1(new_n553_), .A2(new_n563_), .A3(new_n564_), .A4(new_n557_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n562_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n436_), .B1(new_n532_), .B2(new_n535_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT34), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n570_), .A2(KEYINPUT35), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n489_), .A2(new_n503_), .A3(new_n432_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n568_), .A2(new_n571_), .A3(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n573_), .A2(KEYINPUT35), .A3(new_n570_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G190gat), .B(G218gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G134gat), .B(G162gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n577_), .A2(KEYINPUT36), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n570_), .A2(KEYINPUT35), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n568_), .A2(new_n579_), .A3(new_n571_), .A4(new_n572_), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n574_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n577_), .B(KEYINPUT36), .Z(new_n582_));
  INV_X1    g381(.A(KEYINPUT74), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n584_), .B1(new_n574_), .B2(new_n580_), .ZN(new_n585_));
  OAI21_X1  g384(.A(KEYINPUT37), .B1(new_n581_), .B2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n574_), .A2(new_n580_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n587_), .A2(new_n582_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT37), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n574_), .A2(new_n578_), .A3(new_n580_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n588_), .A2(new_n589_), .A3(new_n590_), .ZN(new_n591_));
  AND2_X1   g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n445_), .A2(KEYINPUT75), .A3(new_n446_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(KEYINPUT75), .B1(new_n445_), .B2(new_n446_), .ZN(new_n595_));
  INV_X1    g394(.A(G231gat), .ZN(new_n596_));
  INV_X1    g395(.A(G233gat), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NOR3_X1   g397(.A1(new_n594_), .A2(new_n595_), .A3(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  OAI21_X1  g399(.A(new_n598_), .B1(new_n594_), .B2(new_n595_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n601_), .A3(new_n522_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n598_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n595_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n604_), .B2(new_n593_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n530_), .B1(new_n605_), .B2(new_n599_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT17), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n608_), .B(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G183gat), .B(G211gat), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n610_), .A2(new_n611_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n602_), .A2(new_n606_), .A3(new_n607_), .A4(new_n614_), .ZN(new_n615_));
  OAI21_X1  g414(.A(KEYINPUT17), .B1(new_n612_), .B2(new_n613_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n602_), .A2(new_n606_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n617_), .B1(new_n618_), .B2(KEYINPUT77), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT77), .ZN(new_n620_));
  AOI211_X1 g419(.A(new_n620_), .B(new_n616_), .C1(new_n602_), .C2(new_n606_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n615_), .B1(new_n619_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(KEYINPUT78), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT78), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n615_), .B(new_n624_), .C1(new_n619_), .C2(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n592_), .A2(new_n626_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n466_), .A2(new_n567_), .A3(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n346_), .A2(new_n347_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n441_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT38), .ZN(new_n632_));
  OR2_X1    g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n631_), .A2(new_n632_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n562_), .A2(new_n464_), .A3(new_n565_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT101), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n636_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n420_), .A2(new_n424_), .ZN(new_n640_));
  NOR3_X1   g439(.A1(new_n374_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n422_), .A2(new_n423_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n642_), .B2(new_n374_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n292_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n640_), .B1(new_n643_), .B2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n588_), .A2(new_n590_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n626_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n630_), .ZN(new_n649_));
  NOR3_X1   g448(.A1(new_n639_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n633_), .B(new_n634_), .C1(new_n441_), .C2(new_n650_), .ZN(G1324gat));
  INV_X1    g450(.A(new_n292_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n629_), .A2(new_n442_), .A3(new_n652_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n639_), .A2(new_n648_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n654_), .A2(new_n652_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n656_), .A2(KEYINPUT39), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n442_), .B1(new_n656_), .B2(KEYINPUT39), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n655_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n657_), .B1(new_n655_), .B2(new_n658_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n653_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  XOR2_X1   g460(.A(new_n661_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g461(.A(new_n642_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n654_), .A2(new_n663_), .ZN(new_n664_));
  XOR2_X1   g463(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n665_));
  NAND3_X1  g464(.A1(new_n664_), .A2(G15gat), .A3(new_n665_), .ZN(new_n666_));
  OR3_X1    g465(.A1(new_n628_), .A2(G15gat), .A3(new_n642_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n665_), .B1(new_n664_), .B2(G15gat), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  XOR2_X1   g469(.A(new_n670_), .B(KEYINPUT104), .Z(G1326gat));
  INV_X1    g470(.A(G22gat), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n629_), .A2(new_n672_), .A3(new_n374_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n654_), .A2(new_n374_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n675_), .B2(G22gat), .ZN(new_n676_));
  AOI211_X1 g475(.A(KEYINPUT42), .B(new_n672_), .C1(new_n654_), .C2(new_n374_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n673_), .B1(new_n676_), .B2(new_n677_), .ZN(G1327gat));
  NOR2_X1   g477(.A1(new_n647_), .A2(new_n646_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n680_), .A2(new_n566_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n466_), .A2(new_n681_), .ZN(new_n682_));
  AOI21_X1  g481(.A(G29gat), .B1(new_n682_), .B2(new_n630_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT43), .ZN(new_n684_));
  INV_X1    g483(.A(new_n592_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n684_), .B1(new_n425_), .B2(new_n685_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n645_), .A2(KEYINPUT43), .A3(new_n592_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n686_), .A2(new_n626_), .A3(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT105), .B1(new_n688_), .B2(new_n639_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  OAI211_X1 g490(.A(KEYINPUT105), .B(KEYINPUT44), .C1(new_n688_), .C2(new_n639_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n630_), .A2(G29gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n683_), .B1(new_n693_), .B2(new_n694_), .ZN(G1328gat));
  NOR2_X1   g494(.A1(new_n292_), .A2(G36gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n466_), .A2(new_n681_), .A3(new_n696_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n697_), .A2(KEYINPUT106), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(KEYINPUT106), .ZN(new_n699_));
  AND3_X1   g498(.A1(new_n698_), .A2(KEYINPUT45), .A3(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(KEYINPUT45), .B1(new_n698_), .B2(new_n699_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n292_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n703_));
  INV_X1    g502(.A(G36gat), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n702_), .B1(new_n703_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT46), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n702_), .B(KEYINPUT46), .C1(new_n704_), .C2(new_n703_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(G1329gat));
  NAND2_X1  g508(.A1(new_n682_), .A2(new_n663_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT107), .B(G43gat), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n710_), .A2(KEYINPUT108), .A3(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT108), .B1(new_n710_), .B2(new_n711_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n406_), .A2(G43gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  XNOR2_X1  g516(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n718_), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n714_), .A2(new_n716_), .A3(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1330gat));
  AOI21_X1  g521(.A(G50gat), .B1(new_n682_), .B2(new_n374_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n374_), .A2(G50gat), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n723_), .B1(new_n693_), .B2(new_n724_), .ZN(G1331gat));
  NOR2_X1   g524(.A1(new_n567_), .A2(new_n464_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(new_n648_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n728_), .ZN(new_n729_));
  OAI21_X1  g528(.A(G57gat), .B1(new_n729_), .B2(new_n649_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n566_), .A2(KEYINPUT110), .A3(new_n627_), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT110), .B1(new_n566_), .B2(new_n627_), .ZN(new_n732_));
  NOR4_X1   g531(.A1(new_n731_), .A2(new_n425_), .A3(new_n732_), .A4(new_n464_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n733_), .A2(new_n513_), .A3(new_n630_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n730_), .A2(new_n734_), .ZN(G1332gat));
  NAND2_X1  g534(.A1(new_n728_), .A2(new_n652_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT111), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(new_n737_), .A3(G64gat), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT48), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n737_), .B1(new_n736_), .B2(G64gat), .ZN(new_n741_));
  OR3_X1    g540(.A1(new_n739_), .A2(new_n740_), .A3(new_n741_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n740_), .B1(new_n739_), .B2(new_n741_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n652_), .A2(new_n511_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT112), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n733_), .A2(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n742_), .A2(new_n743_), .A3(new_n746_), .ZN(G1333gat));
  NAND3_X1  g546(.A1(new_n733_), .A2(new_n380_), .A3(new_n663_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT49), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n728_), .A2(new_n663_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n749_), .B1(new_n750_), .B2(G71gat), .ZN(new_n751_));
  AOI211_X1 g550(.A(KEYINPUT49), .B(new_n380_), .C1(new_n728_), .C2(new_n663_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n748_), .B1(new_n751_), .B2(new_n752_), .ZN(G1334gat));
  NAND3_X1  g552(.A1(new_n733_), .A2(new_n509_), .A3(new_n374_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n728_), .A2(new_n374_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(G78gat), .A3(new_n756_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G78gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(G1335gat));
  NAND4_X1  g558(.A1(new_n686_), .A2(new_n626_), .A3(new_n687_), .A4(new_n726_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G85gat), .B1(new_n760_), .B2(new_n649_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n425_), .A2(new_n464_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n567_), .A2(new_n680_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n764_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n765_), .A2(new_n491_), .A3(new_n630_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n766_), .ZN(G1336gat));
  NOR2_X1   g566(.A1(new_n493_), .A2(new_n494_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n760_), .A2(new_n768_), .A3(new_n292_), .ZN(new_n769_));
  AOI21_X1  g568(.A(G92gat), .B1(new_n765_), .B2(new_n652_), .ZN(new_n770_));
  NOR2_X1   g569(.A1(new_n769_), .A2(new_n770_), .ZN(G1337gat));
  AND4_X1   g570(.A1(new_n497_), .A2(new_n765_), .A3(new_n498_), .A4(new_n406_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n687_), .A2(new_n626_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT43), .B1(new_n645_), .B2(new_n592_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n775_), .A2(new_n663_), .A3(new_n726_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n772_), .B1(new_n776_), .B2(G99gat), .ZN(new_n777_));
  XOR2_X1   g576(.A(new_n777_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g577(.A1(new_n765_), .A2(new_n478_), .A3(new_n374_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n760_), .A2(new_n403_), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n478_), .B1(new_n781_), .B2(KEYINPUT114), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT114), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n783_), .B1(new_n760_), .B2(new_n403_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n780_), .B1(new_n782_), .B2(new_n784_), .ZN(new_n785_));
  NAND4_X1  g584(.A1(new_n775_), .A2(KEYINPUT114), .A3(new_n374_), .A4(new_n726_), .ZN(new_n786_));
  AND4_X1   g585(.A1(new_n780_), .A2(new_n786_), .A3(G106gat), .A4(new_n784_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n779_), .B1(new_n785_), .B2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT53), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790_));
  OAI211_X1 g589(.A(new_n790_), .B(new_n779_), .C1(new_n785_), .C2(new_n787_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(G1339gat));
  NAND4_X1  g591(.A1(new_n627_), .A2(new_n562_), .A3(new_n465_), .A4(new_n565_), .ZN(new_n793_));
  OR2_X1    g592(.A1(KEYINPUT115), .A2(KEYINPUT54), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n793_), .A2(new_n794_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(KEYINPUT115), .A2(KEYINPUT54), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT116), .Z(new_n797_));
  INV_X1    g596(.A(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n795_), .A2(new_n798_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n793_), .A2(new_n794_), .A3(new_n797_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  AOI211_X1 g602(.A(KEYINPUT12), .B(new_n522_), .C1(new_n489_), .C2(new_n503_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n523_), .A2(new_n524_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(KEYINPUT12), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n803_), .B1(new_n806_), .B2(new_n468_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n541_), .A2(KEYINPUT55), .A3(new_n542_), .ZN(new_n808_));
  OAI21_X1  g607(.A(KEYINPUT117), .B1(new_n541_), .B2(new_n542_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n538_), .A2(new_n810_), .A3(new_n468_), .A4(new_n540_), .ZN(new_n811_));
  NAND4_X1  g610(.A1(new_n807_), .A2(new_n808_), .A3(new_n809_), .A4(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n812_), .A2(new_n555_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(KEYINPUT56), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n812_), .A2(new_n815_), .A3(new_n555_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n814_), .A2(new_n464_), .A3(new_n550_), .A4(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n448_), .A2(new_n449_), .A3(new_n454_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n453_), .A2(new_n450_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n460_), .A3(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n463_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823_));
  XNOR2_X1  g622(.A(new_n822_), .B(new_n823_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n553_), .A2(new_n818_), .A3(new_n557_), .A4(new_n824_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT72), .B1(new_n551_), .B2(new_n552_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n550_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n557_), .B(new_n824_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT119), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n817_), .A2(new_n825_), .A3(new_n829_), .ZN(new_n830_));
  AND3_X1   g629(.A1(new_n830_), .A2(KEYINPUT57), .A3(new_n646_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT57), .B1(new_n830_), .B2(new_n646_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n814_), .A2(new_n550_), .A3(new_n816_), .A4(new_n824_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(KEYINPUT120), .A2(KEYINPUT58), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n815_), .B1(new_n812_), .B2(new_n555_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n837_), .A2(new_n827_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n838_), .A2(new_n834_), .A3(new_n816_), .A4(new_n824_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n685_), .B1(new_n836_), .B2(new_n839_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n831_), .A2(new_n832_), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n802_), .B1(new_n841_), .B2(new_n647_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n649_), .A2(new_n652_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n842_), .A2(new_n843_), .A3(new_n641_), .A4(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n836_), .A2(new_n839_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n592_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT121), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n840_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n816_), .ZN(new_n851_));
  NOR4_X1   g650(.A1(new_n851_), .A2(new_n837_), .A3(new_n465_), .A4(new_n827_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n829_), .A2(new_n825_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n646_), .B1(new_n852_), .B2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n854_), .A2(new_n855_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n830_), .A2(KEYINPUT57), .A3(new_n646_), .ZN(new_n857_));
  NAND4_X1  g656(.A1(new_n848_), .A2(new_n850_), .A3(new_n856_), .A4(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n801_), .B1(new_n858_), .B2(new_n626_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n844_), .A2(new_n641_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n845_), .B1(new_n861_), .B2(new_n843_), .ZN(new_n862_));
  OAI21_X1  g661(.A(G113gat), .B1(new_n862_), .B2(new_n465_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n861_), .ZN(new_n864_));
  OR2_X1    g663(.A1(new_n465_), .A2(G113gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(G1340gat));
  OAI21_X1  g665(.A(G120gat), .B1(new_n862_), .B2(new_n567_), .ZN(new_n867_));
  INV_X1    g666(.A(G120gat), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n567_), .B2(KEYINPUT60), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n869_), .B1(KEYINPUT60), .B2(new_n868_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n867_), .B1(new_n864_), .B2(new_n870_), .ZN(G1341gat));
  OAI21_X1  g670(.A(G127gat), .B1(new_n862_), .B2(new_n626_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n626_), .A2(G127gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n864_), .B2(new_n873_), .ZN(G1342gat));
  OAI21_X1  g673(.A(G134gat), .B1(new_n862_), .B2(new_n685_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n646_), .A2(G134gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n875_), .B1(new_n864_), .B2(new_n876_), .ZN(G1343gat));
  NOR2_X1   g676(.A1(new_n859_), .A2(new_n402_), .ZN(new_n878_));
  NAND3_X1  g677(.A1(new_n878_), .A2(new_n464_), .A3(new_n844_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT122), .B(G141gat), .ZN(new_n880_));
  XOR2_X1   g679(.A(new_n879_), .B(new_n880_), .Z(G1344gat));
  NAND3_X1  g680(.A1(new_n878_), .A2(new_n566_), .A3(new_n844_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(KEYINPUT123), .B(G148gat), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n882_), .B(new_n883_), .ZN(G1345gat));
  NAND3_X1  g683(.A1(new_n878_), .A2(new_n647_), .A3(new_n844_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(KEYINPUT61), .B(G155gat), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n885_), .B(new_n886_), .ZN(G1346gat));
  NAND2_X1  g686(.A1(new_n878_), .A2(new_n844_), .ZN(new_n888_));
  OAI21_X1  g687(.A(G162gat), .B1(new_n888_), .B2(new_n685_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n646_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n306_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n888_), .B2(new_n891_), .ZN(G1347gat));
  AND2_X1   g691(.A1(new_n464_), .A2(new_n258_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n630_), .A2(new_n292_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n663_), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n895_), .A2(new_n374_), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT125), .B1(new_n842_), .B2(new_n896_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n856_), .A2(new_n847_), .A3(new_n857_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n801_), .B1(new_n898_), .B2(new_n626_), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n900_));
  INV_X1    g699(.A(new_n896_), .ZN(new_n901_));
  NOR3_X1   g700(.A1(new_n899_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n893_), .B1(new_n897_), .B2(new_n902_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n898_), .A2(new_n626_), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n901_), .B1(new_n906_), .B2(new_n802_), .ZN(new_n907_));
  AOI211_X1 g706(.A(new_n229_), .B(new_n905_), .C1(new_n907_), .C2(new_n464_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n842_), .A2(new_n464_), .A3(new_n896_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n904_), .B1(new_n909_), .B2(G169gat), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n903_), .B1(new_n908_), .B2(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n911_), .A2(KEYINPUT126), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913_));
  OAI211_X1 g712(.A(new_n903_), .B(new_n913_), .C1(new_n908_), .C2(new_n910_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n912_), .A2(new_n914_), .ZN(G1348gat));
  NOR2_X1   g714(.A1(new_n859_), .A2(new_n374_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n895_), .ZN(new_n917_));
  AND4_X1   g716(.A1(G176gat), .A2(new_n916_), .A3(new_n566_), .A4(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n897_), .A2(new_n902_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n919_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(new_n566_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n918_), .B1(new_n921_), .B2(new_n228_), .ZN(G1349gat));
  NOR3_X1   g721(.A1(new_n919_), .A2(new_n263_), .A3(new_n626_), .ZN(new_n923_));
  INV_X1    g722(.A(new_n210_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n916_), .A2(new_n647_), .A3(new_n917_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n923_), .B1(new_n924_), .B2(new_n925_), .ZN(G1350gat));
  OAI21_X1  g725(.A(G190gat), .B1(new_n919_), .B2(new_n685_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n890_), .A2(new_n209_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n919_), .B2(new_n928_), .ZN(G1351gat));
  NAND3_X1  g728(.A1(new_n878_), .A2(new_n464_), .A3(new_n894_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g730(.A1(new_n878_), .A2(new_n566_), .A3(new_n894_), .ZN(new_n932_));
  XNOR2_X1  g731(.A(new_n932_), .B(G204gat), .ZN(G1353gat));
  NAND3_X1  g732(.A1(new_n878_), .A2(new_n647_), .A3(new_n894_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(KEYINPUT63), .B(G211gat), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n934_), .A2(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n934_), .B2(new_n937_), .ZN(G1354gat));
  INV_X1    g737(.A(new_n859_), .ZN(new_n939_));
  INV_X1    g738(.A(new_n402_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n646_), .A2(G218gat), .ZN(new_n941_));
  NAND4_X1  g740(.A1(new_n939_), .A2(new_n940_), .A3(new_n894_), .A4(new_n941_), .ZN(new_n942_));
  INV_X1    g741(.A(new_n894_), .ZN(new_n943_));
  NOR4_X1   g742(.A1(new_n859_), .A2(new_n402_), .A3(new_n685_), .A4(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(G218gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n942_), .B1(new_n944_), .B2(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n946_), .A2(KEYINPUT127), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948_));
  OAI211_X1 g747(.A(new_n942_), .B(new_n948_), .C1(new_n944_), .C2(new_n945_), .ZN(new_n949_));
  NAND2_X1  g748(.A1(new_n947_), .A2(new_n949_), .ZN(G1355gat));
endmodule


