//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n782_, new_n783_, new_n784_,
    new_n786_, new_n787_, new_n788_, new_n789_, new_n790_, new_n791_,
    new_n792_, new_n793_, new_n794_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n893_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n933_, new_n934_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_;
  XNOR2_X1  g000(.A(KEYINPUT84), .B(G99gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT31), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G15gat), .B(G43gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  NAND2_X1  g004(.A1(G227gat), .A2(G233gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n205_), .B(new_n206_), .ZN(new_n207_));
  NOR2_X1   g006(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n208_), .B(G169gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT23), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n210_), .B1(G183gat), .B2(G190gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(KEYINPUT80), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT80), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT23), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(G183gat), .A2(G190gat), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n211_), .B1(new_n215_), .B2(new_n217_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n209_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n212_), .A2(new_n214_), .A3(new_n216_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT81), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n217_), .A2(new_n210_), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n212_), .A2(new_n214_), .A3(KEYINPUT81), .A4(new_n216_), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227_));
  INV_X1    g026(.A(G169gat), .ZN(new_n228_));
  INV_X1    g027(.A(G176gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n228_), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  OAI21_X1  g031(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n230_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT25), .B(G183gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT26), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n237_), .A2(G190gat), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n236_), .B1(KEYINPUT79), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT79), .ZN(new_n240_));
  INV_X1    g039(.A(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT26), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n237_), .A2(G190gat), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n240_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n235_), .B1(new_n239_), .B2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n220_), .B1(new_n226_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT82), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n249_));
  OR2_X1    g048(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n251_));
  AOI22_X1  g050(.A1(new_n250_), .A2(new_n251_), .B1(new_n242_), .B2(new_n240_), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n241_), .A2(KEYINPUT26), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT79), .B1(new_n238_), .B2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n234_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n249_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(KEYINPUT82), .A3(new_n220_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n248_), .A2(new_n257_), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n258_), .B(G71gat), .Z(new_n259_));
  INV_X1    g058(.A(G113gat), .ZN(new_n260_));
  INV_X1    g059(.A(G127gat), .ZN(new_n261_));
  INV_X1    g060(.A(G134gat), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G127gat), .A2(G134gat), .ZN(new_n264_));
  AOI21_X1  g063(.A(new_n260_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n263_), .A2(new_n260_), .A3(new_n264_), .ZN(new_n267_));
  AOI21_X1  g066(.A(G120gat), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n267_), .ZN(new_n269_));
  INV_X1    g068(.A(G120gat), .ZN(new_n270_));
  NOR3_X1   g069(.A1(new_n269_), .A2(new_n270_), .A3(new_n265_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT83), .B(KEYINPUT30), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n259_), .A2(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n259_), .A2(new_n274_), .ZN(new_n276_));
  OAI21_X1  g075(.A(new_n207_), .B1(new_n275_), .B2(new_n276_), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n259_), .A2(new_n274_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n207_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n259_), .A2(new_n274_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT27), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT94), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n284_), .B1(new_n226_), .B2(new_n219_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n249_), .B(KEYINPUT94), .C1(G183gat), .C2(G190gat), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n285_), .A2(new_n209_), .A3(new_n286_), .ZN(new_n287_));
  AND2_X1   g086(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(KEYINPUT89), .A2(G204gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(G197gat), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT90), .ZN(new_n291_));
  INV_X1    g090(.A(G204gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n291_), .B1(new_n292_), .B2(G197gat), .ZN(new_n293_));
  INV_X1    g092(.A(G197gat), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n295_));
  AND3_X1   g094(.A1(new_n290_), .A2(new_n293_), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT21), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G211gat), .A2(G218gat), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  NOR2_X1   g098(.A1(G211gat), .A2(G218gat), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT92), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(G211gat), .ZN(new_n302_));
  INV_X1    g101(.A(G218gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT92), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n305_), .A3(new_n298_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n301_), .A2(new_n306_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n296_), .A2(new_n297_), .A3(new_n307_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n301_), .A2(new_n306_), .ZN(new_n309_));
  NAND4_X1  g108(.A1(new_n290_), .A2(new_n297_), .A3(new_n293_), .A4(new_n295_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT91), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n293_), .A2(new_n295_), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n313_), .A2(KEYINPUT91), .A3(new_n297_), .A4(new_n290_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n309_), .B1(new_n312_), .B2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n294_), .A2(new_n292_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT89), .B(G204gat), .ZN(new_n317_));
  AOI211_X1 g116(.A(new_n297_), .B(new_n316_), .C1(new_n317_), .C2(new_n294_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n308_), .B1(new_n315_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n218_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(new_n238_), .A2(new_n253_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(new_n236_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n235_), .A3(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n287_), .A2(new_n320_), .A3(new_n324_), .ZN(new_n325_));
  AND3_X1   g124(.A1(new_n256_), .A2(KEYINPUT82), .A3(new_n220_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT82), .B1(new_n256_), .B2(new_n220_), .ZN(new_n327_));
  AOI211_X1 g126(.A(new_n309_), .B(new_n318_), .C1(new_n312_), .C2(new_n314_), .ZN(new_n328_));
  OAI22_X1  g127(.A1(new_n326_), .A2(new_n327_), .B1(new_n328_), .B2(new_n308_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n325_), .A2(new_n329_), .A3(KEYINPUT20), .ZN(new_n330_));
  NAND2_X1  g129(.A1(G226gat), .A2(G233gat), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT19), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n287_), .A2(new_n324_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n315_), .A2(new_n319_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n308_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n335_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n320_), .A2(new_n248_), .A3(new_n257_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n339_), .A2(KEYINPUT20), .A3(new_n332_), .A4(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(G8gat), .B(G36gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(KEYINPUT18), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(G64gat), .ZN(new_n344_));
  INV_X1    g143(.A(G92gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n344_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  AND3_X1   g146(.A1(new_n334_), .A2(new_n341_), .A3(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n347_), .B1(new_n334_), .B2(new_n341_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n283_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n340_), .A2(KEYINPUT20), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n320_), .B1(new_n287_), .B2(new_n324_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n351_), .A2(new_n333_), .A3(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT20), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n354_), .B1(new_n258_), .B2(new_n338_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n332_), .B1(new_n355_), .B2(new_n325_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n346_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n357_));
  NOR3_X1   g156(.A1(new_n351_), .A2(new_n332_), .A3(new_n352_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n333_), .B1(new_n355_), .B2(new_n325_), .ZN(new_n359_));
  OAI21_X1  g158(.A(new_n347_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n357_), .A2(new_n360_), .A3(KEYINPUT27), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G78gat), .B(G106gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  XNOR2_X1  g163(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n365_));
  NOR2_X1   g164(.A1(G155gat), .A2(G162gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  OR2_X1    g166(.A1(new_n365_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n365_), .A2(new_n367_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G155gat), .A2(G162gat), .ZN(new_n370_));
  XOR2_X1   g169(.A(new_n370_), .B(KEYINPUT1), .Z(new_n371_));
  NAND3_X1  g170(.A1(new_n368_), .A2(new_n369_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G141gat), .A2(G148gat), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(G141gat), .A2(G148gat), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n372_), .A2(new_n376_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n365_), .B(new_n366_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n375_), .A2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT2), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n373_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n383_));
  OAI21_X1  g182(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n380_), .A2(new_n382_), .A3(new_n383_), .A4(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n378_), .A2(new_n370_), .A3(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n377_), .A2(new_n386_), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT88), .B1(new_n387_), .B2(KEYINPUT29), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n364_), .B1(new_n388_), .B2(new_n338_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n388_), .A2(new_n338_), .A3(new_n364_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n390_), .A2(KEYINPUT93), .A3(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT93), .ZN(new_n393_));
  INV_X1    g192(.A(new_n391_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n393_), .B1(new_n394_), .B2(new_n389_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n376_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n396_), .B1(new_n378_), .B2(new_n371_), .ZN(new_n397_));
  AND4_X1   g196(.A1(new_n368_), .A2(new_n369_), .A3(new_n370_), .A4(new_n385_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G22gat), .B(G50gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n399_), .A2(new_n400_), .A3(new_n402_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n401_), .B1(new_n387_), .B2(KEYINPUT29), .ZN(new_n404_));
  XNOR2_X1  g203(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n403_), .A2(new_n404_), .A3(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n406_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n392_), .A2(new_n395_), .A3(new_n410_), .ZN(new_n411_));
  OAI221_X1 g210(.A(new_n393_), .B1(new_n394_), .B2(new_n389_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n350_), .A2(new_n361_), .A3(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT99), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n350_), .A2(new_n361_), .A3(KEYINPUT99), .A4(new_n413_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n282_), .B1(new_n416_), .B2(new_n417_), .ZN(new_n418_));
  OAI22_X1  g217(.A1(new_n397_), .A2(new_n398_), .B1(new_n271_), .B2(new_n268_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n272_), .A2(new_n377_), .A3(new_n386_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(KEYINPUT95), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT95), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n399_), .A2(new_n422_), .A3(new_n272_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n421_), .A2(KEYINPUT4), .A3(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G225gat), .A2(G233gat), .ZN(new_n425_));
  XOR2_X1   g224(.A(new_n425_), .B(KEYINPUT96), .Z(new_n426_));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n419_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n424_), .A2(new_n426_), .A3(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G1gat), .B(G29gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(G85gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n431_), .B(KEYINPUT0), .ZN(new_n432_));
  INV_X1    g231(.A(G57gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n432_), .B(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n426_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n421_), .A2(new_n436_), .A3(new_n423_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n429_), .A2(new_n435_), .A3(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT98), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n435_), .B1(new_n429_), .B2(new_n437_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  AOI211_X1 g241(.A(new_n439_), .B(new_n435_), .C1(new_n429_), .C2(new_n437_), .ZN(new_n443_));
  NOR2_X1   g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n277_), .A2(new_n281_), .ZN(new_n446_));
  OAI211_X1 g245(.A(new_n350_), .B(new_n361_), .C1(new_n442_), .C2(new_n443_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n413_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n446_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(new_n441_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n450_), .A2(new_n439_), .A3(new_n438_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n346_), .A2(KEYINPUT32), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT97), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n453_), .B1(new_n334_), .B2(new_n341_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n330_), .A2(new_n332_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n339_), .A2(KEYINPUT20), .A3(new_n340_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n455_), .B1(new_n332_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n452_), .B1(new_n454_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n443_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n452_), .A2(KEYINPUT97), .ZN(new_n460_));
  OAI21_X1  g259(.A(new_n460_), .B1(new_n356_), .B2(new_n353_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n451_), .A2(new_n458_), .A3(new_n459_), .A4(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n441_), .A2(KEYINPUT33), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n348_), .A2(new_n349_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n424_), .A2(new_n428_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n434_), .B1(new_n465_), .B2(new_n436_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n421_), .A2(new_n423_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n466_), .B1(new_n436_), .B2(new_n467_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n441_), .A2(KEYINPUT33), .ZN(new_n469_));
  NAND4_X1  g268(.A1(new_n463_), .A2(new_n464_), .A3(new_n468_), .A4(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n462_), .A2(new_n470_), .A3(new_n413_), .ZN(new_n471_));
  AOI22_X1  g270(.A1(new_n418_), .A2(new_n445_), .B1(new_n449_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT78), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G29gat), .B(G36gat), .ZN(new_n474_));
  INV_X1    g273(.A(G43gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n474_), .B(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(G50gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n474_), .B(G43gat), .ZN(new_n478_));
  INV_X1    g277(.A(G50gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  AND2_X1   g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G15gat), .B(G22gat), .ZN(new_n482_));
  INV_X1    g281(.A(G1gat), .ZN(new_n483_));
  INV_X1    g282(.A(G8gat), .ZN(new_n484_));
  OAI21_X1  g283(.A(KEYINPUT14), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G1gat), .B(G8gat), .ZN(new_n487_));
  XOR2_X1   g286(.A(new_n486_), .B(new_n487_), .Z(new_n488_));
  NAND2_X1  g287(.A1(new_n481_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT77), .ZN(new_n490_));
  INV_X1    g289(.A(new_n488_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n477_), .A2(new_n480_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n489_), .A2(new_n490_), .A3(new_n493_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n491_), .A2(new_n492_), .A3(KEYINPUT77), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G229gat), .A2(G233gat), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT15), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n492_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n477_), .A2(new_n480_), .A3(KEYINPUT15), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n488_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n497_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n491_), .A2(new_n492_), .ZN(new_n504_));
  NOR3_X1   g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n473_), .B1(new_n498_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G113gat), .B(G141gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(new_n228_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(new_n508_), .B(new_n294_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n506_), .B(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G120gat), .B(G148gat), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n513_), .B(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G176gat), .B(G204gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  NAND2_X1  g316(.A1(G230gat), .A2(G233gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT65), .ZN(new_n519_));
  OAI22_X1  g318(.A1(new_n519_), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT7), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n520_), .B1(KEYINPUT65), .B2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G99gat), .A2(G106gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT6), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n519_), .B(KEYINPUT7), .C1(G99gat), .C2(G106gat), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n522_), .A2(new_n524_), .A3(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G85gat), .B(G92gat), .Z(new_n527_));
  INV_X1    g326(.A(KEYINPUT8), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n528_), .A2(KEYINPUT66), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n527_), .A2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n526_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT67), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n531_), .B(KEYINPUT66), .C1(new_n532_), .C2(new_n528_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n527_), .A2(KEYINPUT9), .ZN(new_n534_));
  AND2_X1   g333(.A1(new_n534_), .A2(new_n524_), .ZN(new_n535_));
  INV_X1    g334(.A(G85gat), .ZN(new_n536_));
  OR3_X1    g335(.A1(new_n536_), .A2(new_n345_), .A3(KEYINPUT9), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT64), .ZN(new_n538_));
  XNOR2_X1  g337(.A(KEYINPUT10), .B(G99gat), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n538_), .B1(new_n539_), .B2(G106gat), .ZN(new_n540_));
  OR3_X1    g339(.A1(new_n539_), .A2(new_n538_), .A3(G106gat), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n535_), .A2(new_n537_), .A3(new_n540_), .A4(new_n541_), .ZN(new_n542_));
  OAI21_X1  g341(.A(KEYINPUT66), .B1(new_n532_), .B2(new_n528_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n526_), .A2(new_n543_), .A3(new_n530_), .ZN(new_n544_));
  XOR2_X1   g343(.A(G71gat), .B(G78gat), .Z(new_n545_));
  INV_X1    g344(.A(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G57gat), .B(G64gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(KEYINPUT11), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  OR2_X1    g348(.A1(new_n547_), .A2(KEYINPUT11), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n545_), .A2(KEYINPUT11), .A3(new_n547_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n549_), .A2(new_n550_), .A3(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n533_), .A2(new_n542_), .A3(new_n544_), .A4(new_n553_), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT68), .ZN(new_n555_));
  NAND3_X1  g354(.A1(new_n533_), .A2(new_n542_), .A3(new_n544_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n556_), .A2(new_n552_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n518_), .B1(new_n555_), .B2(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT12), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n557_), .A2(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n556_), .A2(KEYINPUT12), .A3(new_n552_), .ZN(new_n561_));
  NAND4_X1  g360(.A1(new_n560_), .A2(new_n518_), .A3(new_n554_), .A4(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n517_), .B1(new_n558_), .B2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n518_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT68), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n554_), .B(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n557_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n565_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n517_), .ZN(new_n570_));
  NAND3_X1  g369(.A1(new_n569_), .A2(new_n562_), .A3(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n564_), .A2(KEYINPUT13), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(KEYINPUT13), .B1(new_n564_), .B2(new_n571_), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n472_), .A2(new_n512_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT70), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT34), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n531_), .B(new_n543_), .ZN(new_n581_));
  AOI22_X1  g380(.A1(new_n581_), .A2(new_n542_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n556_), .A2(new_n492_), .ZN(new_n583_));
  OAI211_X1 g382(.A(KEYINPUT35), .B(new_n580_), .C1(new_n582_), .C2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n500_), .A2(new_n501_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n556_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n587_));
  OR2_X1    g386(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n581_), .A2(new_n481_), .A3(new_n542_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n586_), .A2(new_n587_), .A3(new_n588_), .A4(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(G162gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(G190gat), .B(G218gat), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT71), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(G134gat), .ZN(new_n594_));
  INV_X1    g393(.A(new_n594_), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n593_), .A2(G134gat), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n591_), .B1(new_n595_), .B2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT36), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n593_), .A2(G134gat), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n599_), .A2(G162gat), .A3(new_n594_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n597_), .A2(new_n598_), .A3(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(KEYINPUT72), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND4_X1  g402(.A1(new_n597_), .A2(new_n600_), .A3(KEYINPUT72), .A4(new_n598_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n584_), .A2(new_n590_), .A3(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT73), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n584_), .A2(KEYINPUT73), .A3(new_n590_), .A4(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n584_), .A2(new_n590_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n597_), .A2(new_n600_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT36), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(new_n601_), .A3(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT74), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n615_), .A2(new_n616_), .A3(KEYINPUT37), .ZN(new_n617_));
  INV_X1    g416(.A(new_n601_), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n584_), .B2(new_n590_), .ZN(new_n619_));
  AOI22_X1  g418(.A1(new_n608_), .A2(new_n609_), .B1(new_n613_), .B2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT37), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT74), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n619_), .A2(KEYINPUT75), .A3(new_n613_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT75), .B1(new_n619_), .B2(new_n613_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n621_), .B(new_n610_), .C1(new_n624_), .C2(new_n625_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n617_), .A2(new_n622_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n488_), .B(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(new_n553_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT17), .ZN(new_n632_));
  XNOR2_X1  g431(.A(G127gat), .B(G155gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT16), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(G183gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(new_n302_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n631_), .B1(new_n632_), .B2(new_n636_), .ZN(new_n637_));
  NOR3_X1   g436(.A1(new_n636_), .A2(KEYINPUT76), .A3(new_n632_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n638_), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n640_), .A2(new_n631_), .ZN(new_n641_));
  OR2_X1    g440(.A1(new_n639_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n628_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n577_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n646_), .A2(new_n483_), .A3(new_n444_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT38), .ZN(new_n648_));
  INV_X1    g447(.A(new_n625_), .ZN(new_n649_));
  AOI22_X1  g448(.A1(new_n649_), .A2(new_n623_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n650_), .A2(new_n643_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n577_), .A2(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n652_), .A2(new_n444_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n648_), .B1(new_n483_), .B2(new_n653_), .ZN(G1324gat));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n350_), .A2(new_n361_), .ZN(new_n658_));
  AOI211_X1 g457(.A(new_n484_), .B(new_n657_), .C1(new_n652_), .C2(new_n658_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n659_), .B1(KEYINPUT100), .B2(KEYINPUT39), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n646_), .A2(new_n484_), .A3(new_n658_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n652_), .A2(new_n658_), .ZN(new_n662_));
  OAI211_X1 g461(.A(new_n655_), .B(new_n656_), .C1(new_n662_), .C2(new_n484_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n660_), .A2(new_n661_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  NAND4_X1  g465(.A1(new_n660_), .A2(KEYINPUT40), .A3(new_n661_), .A4(new_n663_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(G1325gat));
  OR3_X1    g467(.A1(new_n645_), .A2(G15gat), .A3(new_n282_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n416_), .A2(new_n417_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(new_n445_), .A3(new_n446_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n449_), .A2(new_n471_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n576_), .A2(new_n512_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(new_n446_), .A4(new_n651_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(new_n676_), .A3(G15gat), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n676_), .B1(new_n675_), .B2(G15gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT101), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n675_), .A2(G15gat), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n681_), .A2(KEYINPUT102), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n682_), .A2(new_n683_), .A3(new_n677_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n680_), .A2(new_n684_), .A3(KEYINPUT41), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT41), .B1(new_n680_), .B2(new_n684_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n669_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT103), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n689_));
  OAI211_X1 g488(.A(new_n689_), .B(new_n669_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n688_), .A2(new_n690_), .ZN(G1326gat));
  INV_X1    g490(.A(G22gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n692_), .B1(new_n652_), .B2(new_n448_), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT42), .Z(new_n694_));
  NAND3_X1  g493(.A1(new_n646_), .A2(new_n692_), .A3(new_n448_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(G1327gat));
  INV_X1    g495(.A(new_n650_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n697_), .A2(new_n642_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n577_), .A2(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(G29gat), .B1(new_n700_), .B2(new_n444_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n674_), .A2(new_n643_), .ZN(new_n703_));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n472_), .B2(new_n627_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n449_), .A2(new_n471_), .ZN(new_n706_));
  AOI211_X1 g505(.A(new_n444_), .B(new_n282_), .C1(new_n416_), .C2(new_n417_), .ZN(new_n707_));
  OAI211_X1 g506(.A(new_n705_), .B(new_n628_), .C1(new_n706_), .C2(new_n707_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n703_), .B1(new_n704_), .B2(new_n708_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n702_), .B1(new_n709_), .B2(KEYINPUT104), .ZN(new_n710_));
  INV_X1    g509(.A(new_n703_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n705_), .B1(new_n673_), .B2(new_n628_), .ZN(new_n712_));
  AOI211_X1 g511(.A(KEYINPUT43), .B(new_n627_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n711_), .B1(new_n712_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n714_), .A2(new_n715_), .A3(KEYINPUT44), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n710_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n718_), .A2(new_n445_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n701_), .B1(new_n719_), .B2(G29gat), .ZN(G1328gat));
  AOI21_X1  g519(.A(KEYINPUT44), .B1(new_n714_), .B2(new_n715_), .ZN(new_n721_));
  NOR3_X1   g520(.A1(new_n709_), .A2(KEYINPUT104), .A3(new_n702_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n658_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G36gat), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT46), .ZN(new_n726_));
  INV_X1    g525(.A(G36gat), .ZN(new_n727_));
  NAND4_X1  g526(.A1(new_n577_), .A2(new_n727_), .A3(new_n658_), .A4(new_n698_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND4_X1  g530(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .A4(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n725_), .A2(new_n726_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n727_), .B1(new_n717_), .B2(new_n658_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n733_), .B(new_n734_), .C1(new_n735_), .C2(new_n730_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n732_), .A2(new_n736_), .ZN(G1329gat));
  AOI21_X1  g536(.A(new_n475_), .B1(new_n717_), .B2(new_n446_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT47), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n699_), .A2(G43gat), .A3(new_n282_), .ZN(new_n740_));
  OR3_X1    g539(.A1(new_n738_), .A2(new_n739_), .A3(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n738_), .B2(new_n740_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1330gat));
  OAI21_X1  g542(.A(G50gat), .B1(new_n718_), .B2(new_n413_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n700_), .A2(new_n479_), .A3(new_n448_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n744_), .A2(new_n745_), .ZN(G1331gat));
  NOR2_X1   g545(.A1(new_n575_), .A2(new_n511_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n673_), .A2(new_n651_), .A3(new_n747_), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n748_), .A2(new_n433_), .A3(new_n445_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n472_), .A2(new_n511_), .A3(new_n575_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n750_), .A2(new_n444_), .A3(new_n644_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n749_), .B1(new_n433_), .B2(new_n751_), .ZN(G1332gat));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n644_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n658_), .ZN(new_n754_));
  OR3_X1    g553(.A1(new_n753_), .A2(G64gat), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(G64gat), .B1(new_n748_), .B2(new_n754_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n756_), .A2(KEYINPUT107), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(KEYINPUT107), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n757_), .A2(KEYINPUT48), .A3(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT48), .B1(new_n757_), .B2(new_n758_), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n755_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT108), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT108), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n763_), .B(new_n755_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1333gat));
  OAI21_X1  g564(.A(G71gat), .B1(new_n748_), .B2(new_n282_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT49), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n282_), .A2(G71gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n753_), .B2(new_n768_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT109), .Z(G1334gat));
  OAI21_X1  g569(.A(G78gat), .B1(new_n748_), .B2(new_n413_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT50), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n413_), .A2(G78gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n753_), .B2(new_n773_), .ZN(G1335gat));
  NAND2_X1  g573(.A1(new_n750_), .A2(new_n698_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n536_), .B1(new_n775_), .B2(new_n445_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT110), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n704_), .A2(new_n708_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n778_), .A2(new_n643_), .A3(new_n747_), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n779_), .A2(new_n536_), .A3(new_n445_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n777_), .A2(new_n780_), .ZN(G1336gat));
  NOR3_X1   g580(.A1(new_n779_), .A2(new_n345_), .A3(new_n754_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n775_), .ZN(new_n783_));
  AOI21_X1  g582(.A(G92gat), .B1(new_n783_), .B2(new_n658_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1337gat));
  NAND4_X1  g584(.A1(new_n778_), .A2(new_n446_), .A3(new_n643_), .A4(new_n747_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(G99gat), .ZN(new_n787_));
  OR3_X1    g586(.A1(new_n775_), .A2(new_n539_), .A3(new_n282_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT112), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n787_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT51), .ZN(new_n791_));
  OR3_X1    g590(.A1(new_n790_), .A2(KEYINPUT111), .A3(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n787_), .A2(new_n788_), .A3(KEYINPUT111), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n791_), .B1(new_n790_), .B2(KEYINPUT111), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n792_), .A2(new_n793_), .A3(new_n794_), .ZN(G1338gat));
  OR3_X1    g594(.A1(new_n775_), .A2(G106gat), .A3(new_n413_), .ZN(new_n796_));
  NAND4_X1  g595(.A1(new_n778_), .A2(new_n448_), .A3(new_n643_), .A4(new_n747_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT52), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n797_), .A2(new_n798_), .A3(G106gat), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n798_), .B1(new_n797_), .B2(G106gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n573_), .A2(new_n511_), .A3(new_n574_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n627_), .A2(new_n803_), .A3(new_n804_), .A4(new_n642_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT54), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n627_), .A2(new_n642_), .A3(new_n804_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n807_), .A2(KEYINPUT113), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n806_), .B(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n560_), .A2(new_n561_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n565_), .B1(new_n810_), .B2(new_n567_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n556_), .A2(KEYINPUT12), .A3(new_n552_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT12), .B1(new_n556_), .B2(new_n552_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND4_X1  g613(.A1(new_n814_), .A2(KEYINPUT55), .A3(new_n518_), .A4(new_n554_), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT55), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n562_), .A2(new_n816_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n811_), .A2(new_n815_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT56), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n819_), .A3(new_n517_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n819_), .B1(new_n818_), .B2(new_n517_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n571_), .ZN(new_n823_));
  NOR3_X1   g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n498_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n496_), .A2(new_n497_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n503_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n510_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n825_), .A2(new_n828_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n824_), .A2(KEYINPUT115), .A3(KEYINPUT58), .A4(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT115), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n818_), .A2(new_n517_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n832_), .A2(KEYINPUT56), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n833_), .A2(new_n571_), .A3(new_n829_), .A4(new_n820_), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n831_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  XNOR2_X1  g635(.A(KEYINPUT114), .B(KEYINPUT58), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n834_), .A2(new_n837_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n830_), .A2(new_n836_), .A3(new_n628_), .A4(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n833_), .A2(new_n511_), .A3(new_n571_), .A4(new_n820_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n564_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n829_), .B1(new_n841_), .B2(new_n823_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n843_), .A2(new_n697_), .ZN(new_n844_));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n843_), .A2(KEYINPUT57), .A3(new_n697_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n839_), .A2(new_n846_), .A3(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(new_n643_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n809_), .A2(KEYINPUT116), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT57), .B1(new_n843_), .B2(new_n697_), .ZN(new_n852_));
  AOI211_X1 g651(.A(new_n845_), .B(new_n650_), .C1(new_n840_), .C2(new_n842_), .ZN(new_n853_));
  NOR2_X1   g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n642_), .B1(new_n854_), .B2(new_n839_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n808_), .A2(KEYINPUT54), .A3(new_n805_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT54), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n807_), .A2(KEYINPUT113), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n856_), .A2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n851_), .B1(new_n855_), .B2(new_n859_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n418_), .A2(new_n444_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n850_), .A2(new_n860_), .A3(new_n861_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n260_), .B1(new_n862_), .B2(new_n512_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT117), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(KEYINPUT59), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n809_), .A2(new_n849_), .ZN(new_n866_));
  XOR2_X1   g665(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n861_), .A3(new_n867_), .ZN(new_n868_));
  NAND4_X1  g667(.A1(new_n865_), .A2(G113gat), .A3(new_n511_), .A4(new_n868_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n870_));
  OAI211_X1 g669(.A(new_n870_), .B(new_n260_), .C1(new_n862_), .C2(new_n512_), .ZN(new_n871_));
  AND3_X1   g670(.A1(new_n864_), .A2(new_n869_), .A3(new_n871_), .ZN(G1340gat));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n575_), .B2(G120gat), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n850_), .A2(new_n860_), .A3(new_n861_), .A4(new_n874_), .ZN(new_n875_));
  NAND4_X1  g674(.A1(new_n865_), .A2(new_n576_), .A3(new_n868_), .A4(new_n875_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(G120gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(KEYINPUT60), .B2(new_n875_), .ZN(G1341gat));
  AND2_X1   g677(.A1(new_n865_), .A2(new_n868_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n643_), .A2(new_n261_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n850_), .A2(new_n860_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n881_), .A2(new_n642_), .A3(new_n861_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n879_), .A2(new_n880_), .B1(new_n261_), .B2(new_n882_), .ZN(G1342gat));
  NOR2_X1   g682(.A1(new_n627_), .A2(new_n262_), .ZN(new_n884_));
  NAND3_X1  g683(.A1(new_n881_), .A2(new_n650_), .A3(new_n861_), .ZN(new_n885_));
  AOI22_X1  g684(.A1(new_n879_), .A2(new_n884_), .B1(new_n262_), .B2(new_n885_), .ZN(G1343gat));
  NOR2_X1   g685(.A1(new_n446_), .A2(new_n413_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n445_), .A2(new_n658_), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n850_), .A2(new_n860_), .A3(new_n887_), .A4(new_n888_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n889_), .A2(new_n512_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT119), .B(G141gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1344gat));
  NOR2_X1   g691(.A1(new_n889_), .A2(new_n575_), .ZN(new_n893_));
  XOR2_X1   g692(.A(new_n893_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g693(.A1(new_n889_), .A2(new_n643_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT61), .B(G155gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(KEYINPUT120), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n895_), .B(new_n897_), .ZN(G1346gat));
  NAND2_X1  g697(.A1(new_n628_), .A2(G162gat), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(KEYINPUT122), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n889_), .A2(new_n900_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n591_), .B1(new_n889_), .B2(new_n697_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(KEYINPUT121), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n904_), .B(new_n591_), .C1(new_n889_), .C2(new_n697_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n901_), .B1(new_n903_), .B2(new_n905_), .ZN(G1347gat));
  XNOR2_X1  g705(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NOR2_X1   g707(.A1(new_n754_), .A2(new_n444_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(new_n446_), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(KEYINPUT123), .Z(new_n911_));
  NAND3_X1  g710(.A1(new_n866_), .A2(new_n413_), .A3(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n511_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n908_), .B1(new_n914_), .B2(G169gat), .ZN(new_n915_));
  OAI211_X1 g714(.A(G169gat), .B(new_n908_), .C1(new_n912_), .C2(new_n512_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(KEYINPUT22), .B(G169gat), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n511_), .A2(new_n918_), .ZN(new_n919_));
  XOR2_X1   g718(.A(new_n919_), .B(KEYINPUT125), .Z(new_n920_));
  OAI22_X1  g719(.A1(new_n915_), .A2(new_n917_), .B1(new_n912_), .B2(new_n920_), .ZN(G1348gat));
  AOI21_X1  g720(.A(G176gat), .B1(new_n913_), .B2(new_n576_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n881_), .A2(new_n413_), .ZN(new_n923_));
  AND3_X1   g722(.A1(new_n911_), .A2(G176gat), .A3(new_n576_), .ZN(new_n924_));
  AOI21_X1  g723(.A(new_n922_), .B1(new_n923_), .B2(new_n924_), .ZN(G1349gat));
  NOR3_X1   g724(.A1(new_n912_), .A2(new_n236_), .A3(new_n643_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n923_), .A2(new_n642_), .A3(new_n911_), .ZN(new_n927_));
  INV_X1    g726(.A(G183gat), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n926_), .B1(new_n927_), .B2(new_n928_), .ZN(G1350gat));
  OAI21_X1  g728(.A(G190gat), .B1(new_n912_), .B2(new_n627_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n650_), .A2(new_n322_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n912_), .B2(new_n931_), .ZN(G1351gat));
  NAND4_X1  g731(.A1(new_n850_), .A2(new_n860_), .A3(new_n887_), .A4(new_n909_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(new_n512_), .ZN(new_n934_));
  XNOR2_X1  g733(.A(new_n934_), .B(new_n294_), .ZN(G1352gat));
  NOR2_X1   g734(.A1(new_n933_), .A2(new_n575_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(new_n317_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n937_), .B1(new_n292_), .B2(new_n936_), .ZN(G1353gat));
  NOR2_X1   g737(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n939_));
  AND4_X1   g738(.A1(new_n860_), .A2(new_n850_), .A3(new_n887_), .A4(new_n909_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n939_), .B1(new_n940_), .B2(new_n642_), .ZN(new_n941_));
  XOR2_X1   g740(.A(KEYINPUT63), .B(G211gat), .Z(new_n942_));
  NOR3_X1   g741(.A1(new_n933_), .A2(new_n643_), .A3(new_n942_), .ZN(new_n943_));
  OAI21_X1  g742(.A(KEYINPUT126), .B1(new_n941_), .B2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n945_));
  OAI22_X1  g744(.A1(new_n933_), .A2(new_n643_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n940_), .A2(new_n642_), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n945_), .B(new_n946_), .C1(new_n947_), .C2(new_n942_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n944_), .A2(new_n948_), .ZN(G1354gat));
  AOI21_X1  g748(.A(G218gat), .B1(new_n940_), .B2(new_n650_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n628_), .A2(G218gat), .ZN(new_n951_));
  XNOR2_X1  g750(.A(new_n951_), .B(KEYINPUT127), .ZN(new_n952_));
  AOI21_X1  g751(.A(new_n950_), .B1(new_n940_), .B2(new_n952_), .ZN(G1355gat));
endmodule


