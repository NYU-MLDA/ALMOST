//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n768_, new_n769_, new_n770_, new_n772_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n876_, new_n877_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n921_, new_n922_, new_n924_,
    new_n925_, new_n926_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_;
  INV_X1    g000(.A(G50gat), .ZN(new_n202_));
  INV_X1    g001(.A(G29gat), .ZN(new_n203_));
  INV_X1    g002(.A(G36gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G43gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n205_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n206_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n202_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n210_), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G50gat), .A3(new_n208_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215_));
  INV_X1    g014(.A(G1gat), .ZN(new_n216_));
  INV_X1    g015(.A(G8gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT14), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n215_), .A2(new_n218_), .ZN(new_n219_));
  XNOR2_X1  g018(.A(G1gat), .B(G8gat), .ZN(new_n220_));
  XNOR2_X1  g019(.A(new_n219_), .B(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n214_), .A2(new_n221_), .ZN(new_n222_));
  AND3_X1   g021(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT15), .ZN(new_n223_));
  AOI21_X1  g022(.A(KEYINPUT15), .B1(new_n211_), .B2(new_n213_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n222_), .B1(new_n226_), .B2(new_n221_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(G229gat), .A2(G233gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n214_), .B(new_n221_), .ZN(new_n230_));
  INV_X1    g029(.A(new_n228_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G113gat), .B(G141gat), .ZN(new_n234_));
  INV_X1    g033(.A(G169gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(G197gat), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n233_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n233_), .A2(new_n238_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT12), .ZN(new_n243_));
  XOR2_X1   g042(.A(KEYINPUT10), .B(G99gat), .Z(new_n244_));
  INV_X1    g043(.A(G106gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT65), .ZN(new_n247_));
  AND3_X1   g046(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G99gat), .A2(G106gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT6), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n253_), .A2(KEYINPUT65), .A3(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(G85gat), .ZN(new_n256_));
  INV_X1    g055(.A(G92gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(G85gat), .A2(G92gat), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n258_), .A2(KEYINPUT9), .A3(new_n259_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n246_), .A2(new_n250_), .A3(new_n255_), .A4(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n259_), .A2(KEYINPUT9), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  NOR3_X1   g064(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n268_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n253_), .A2(KEYINPUT66), .A3(new_n254_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n267_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  AND2_X1   g070(.A1(new_n258_), .A2(new_n259_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT8), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n267_), .A2(new_n250_), .A3(new_n255_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT8), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(new_n272_), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n263_), .B1(new_n274_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT11), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT67), .B(G71gat), .ZN(new_n280_));
  INV_X1    g079(.A(G78gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(G71gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT67), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT67), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(G71gat), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n284_), .A2(new_n286_), .A3(new_n281_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n279_), .B1(new_n282_), .B2(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n284_), .A2(new_n286_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G78gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n280_), .A2(new_n281_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n290_), .A2(new_n291_), .A3(KEYINPUT11), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G57gat), .B(G64gat), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n288_), .A2(new_n292_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n293_), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n290_), .A2(new_n291_), .A3(KEYINPUT11), .A4(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n294_), .A2(new_n296_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n243_), .B1(new_n278_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n278_), .A2(new_n297_), .ZN(new_n299_));
  AND2_X1   g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(G230gat), .A2(G233gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n301_), .B(KEYINPUT64), .Z(new_n302_));
  OR2_X1    g101(.A1(new_n261_), .A2(new_n262_), .ZN(new_n303_));
  AND2_X1   g102(.A1(new_n272_), .A2(new_n276_), .ZN(new_n304_));
  AND2_X1   g103(.A1(new_n304_), .A2(new_n275_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n276_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n307_));
  NOR3_X1   g106(.A1(new_n305_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(KEYINPUT68), .B1(new_n274_), .B2(new_n277_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n303_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n297_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(KEYINPUT12), .A3(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n300_), .A2(new_n302_), .A3(new_n312_), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n278_), .A2(new_n297_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(new_n299_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n302_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G120gat), .B(G148gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT5), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(G176gat), .ZN(new_n320_));
  INV_X1    g119(.A(G204gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n320_), .B(new_n321_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n313_), .A2(new_n317_), .A3(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n324_), .B(KEYINPUT69), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n313_), .A2(new_n317_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(new_n322_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n325_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT70), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT13), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n328_), .A2(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(new_n325_), .B2(new_n327_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT71), .B1(new_n332_), .B2(new_n334_), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n325_), .B(new_n327_), .C1(new_n329_), .C2(new_n330_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT71), .ZN(new_n337_));
  INV_X1    g136(.A(new_n328_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n336_), .B(new_n337_), .C1(new_n338_), .C2(new_n333_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n242_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G225gat), .A2(G233gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT4), .ZN(new_n344_));
  OR2_X1    g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT1), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n345_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G141gat), .A2(G148gat), .ZN(new_n351_));
  OAI21_X1  g150(.A(KEYINPUT84), .B1(G141gat), .B2(G148gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(G141gat), .A2(G148gat), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT84), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n350_), .A2(new_n351_), .A3(new_n352_), .A4(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT85), .ZN(new_n357_));
  INV_X1    g156(.A(G141gat), .ZN(new_n358_));
  INV_X1    g157(.A(G148gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n353_), .A2(new_n357_), .A3(KEYINPUT3), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n351_), .A2(KEYINPUT2), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT2), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n365_), .A2(G141gat), .A3(G148gat), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n362_), .A2(new_n363_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT86), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n346_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n364_), .A2(new_n366_), .ZN(new_n370_));
  NOR4_X1   g169(.A1(new_n361_), .A2(KEYINPUT85), .A3(G141gat), .A4(G148gat), .ZN(new_n371_));
  AOI21_X1  g170(.A(KEYINPUT3), .B1(new_n353_), .B2(new_n357_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n368_), .B(new_n370_), .C1(new_n371_), .C2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n345_), .ZN(new_n374_));
  OAI21_X1  g173(.A(new_n356_), .B1(new_n369_), .B2(new_n374_), .ZN(new_n375_));
  OR2_X1    g174(.A1(G127gat), .A2(G134gat), .ZN(new_n376_));
  NAND2_X1  g175(.A1(G127gat), .A2(G134gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(G113gat), .ZN(new_n379_));
  INV_X1    g178(.A(G113gat), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n376_), .A2(new_n380_), .A3(new_n377_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n379_), .A2(G120gat), .A3(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(G120gat), .B1(new_n379_), .B2(new_n381_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT93), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n375_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n356_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n373_), .A2(new_n345_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n370_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n390_));
  AOI22_X1  g189(.A1(new_n390_), .A2(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n388_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(new_n384_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n344_), .B1(new_n387_), .B2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n389_), .A2(new_n391_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n384_), .B1(new_n395_), .B2(new_n356_), .ZN(new_n396_));
  AOI21_X1  g195(.A(KEYINPUT4), .B1(new_n396_), .B2(new_n386_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n343_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(new_n396_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n399_), .A2(new_n342_), .A3(new_n393_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n398_), .A2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G1gat), .B(G29gat), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n402_), .B(G85gat), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT0), .ZN(new_n404_));
  XOR2_X1   g203(.A(new_n404_), .B(G57gat), .Z(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n401_), .A2(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n398_), .A2(new_n400_), .A3(new_n405_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n409_), .ZN(new_n410_));
  NOR3_X1   g209(.A1(new_n375_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT28), .ZN(new_n413_));
  INV_X1    g212(.A(KEYINPUT29), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n392_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(G228gat), .A2(G233gat), .ZN(new_n417_));
  INV_X1    g216(.A(G22gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n412_), .A2(new_n416_), .A3(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n419_), .B1(new_n411_), .B2(new_n415_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n421_), .A2(new_n422_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n392_), .A2(new_n414_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n321_), .A2(KEYINPUT88), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT88), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(G204gat), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n425_), .A2(new_n427_), .A3(new_n237_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT87), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n429_), .B1(new_n237_), .B2(G204gat), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n321_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  OAI21_X1  g231(.A(KEYINPUT21), .B1(new_n428_), .B2(new_n432_), .ZN(new_n433_));
  XOR2_X1   g232(.A(G211gat), .B(G218gat), .Z(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n237_), .A2(G204gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT88), .B(G204gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n436_), .B1(new_n437_), .B2(new_n237_), .ZN(new_n438_));
  OAI211_X1 g237(.A(new_n433_), .B(new_n435_), .C1(KEYINPUT21), .C2(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n438_), .A2(KEYINPUT21), .A3(new_n434_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n438_), .A2(KEYINPUT89), .A3(KEYINPUT21), .A4(new_n434_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(new_n442_), .A3(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  OAI21_X1  g244(.A(G50gat), .B1(new_n424_), .B2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G78gat), .B(G106gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n375_), .A2(KEYINPUT29), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n449_), .A2(new_n202_), .A3(new_n444_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n448_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n448_), .B1(new_n446_), .B2(new_n450_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n423_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(G227gat), .A2(G233gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n455_), .B(KEYINPUT30), .ZN(new_n456_));
  XOR2_X1   g255(.A(KEYINPUT80), .B(KEYINPUT81), .Z(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G15gat), .B(G43gat), .Z(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(new_n384_), .ZN(new_n461_));
  INV_X1    g260(.A(G176gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n235_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G169gat), .A2(G176gat), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(KEYINPUT24), .A3(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(KEYINPUT76), .A2(G190gat), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT26), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT26), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n468_), .A2(KEYINPUT76), .A3(G190gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n467_), .A2(new_n469_), .ZN(new_n470_));
  AND2_X1   g269(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n471_));
  NOR2_X1   g270(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n465_), .B1(new_n470_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT77), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  OR2_X1    g275(.A1(new_n463_), .A2(KEYINPUT24), .ZN(new_n477_));
  OAI211_X1 g276(.A(KEYINPUT77), .B(new_n465_), .C1(new_n470_), .C2(new_n473_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(G183gat), .A2(G190gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n479_), .B(KEYINPUT23), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .A4(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT79), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(G183gat), .B2(G190gat), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT78), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n484_), .B1(new_n235_), .B2(KEYINPUT22), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT22), .B(G169gat), .ZN(new_n486_));
  OAI211_X1 g285(.A(new_n462_), .B(new_n485_), .C1(new_n486_), .C2(new_n484_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n483_), .A2(new_n487_), .A3(new_n464_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n481_), .A2(new_n482_), .A3(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n482_), .B1(new_n481_), .B2(new_n488_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(KEYINPUT82), .B(KEYINPUT31), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT83), .ZN(new_n492_));
  XOR2_X1   g291(.A(G71gat), .B(G99gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n489_), .A2(new_n490_), .A3(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n461_), .A2(new_n496_), .A3(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n460_), .B(new_n385_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n497_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n499_), .B1(new_n500_), .B2(new_n495_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n498_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n450_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n202_), .B1(new_n449_), .B2(new_n444_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n447_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n505_), .A2(new_n421_), .A3(new_n422_), .A4(new_n451_), .ZN(new_n506_));
  AND3_X1   g305(.A1(new_n454_), .A2(new_n502_), .A3(new_n506_), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n502_), .B1(new_n454_), .B2(new_n506_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n481_), .A2(new_n488_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT79), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n481_), .A2(new_n482_), .A3(new_n488_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n511_), .A2(new_n512_), .A3(new_n445_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT92), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n483_), .A2(new_n514_), .ZN(new_n515_));
  OAI211_X1 g314(.A(new_n480_), .B(KEYINPUT92), .C1(G183gat), .C2(G190gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n486_), .A2(new_n462_), .ZN(new_n517_));
  NAND4_X1  g316(.A1(new_n515_), .A2(new_n464_), .A3(new_n516_), .A4(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n463_), .A2(new_n464_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n520_));
  OR2_X1    g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT26), .B(G190gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(new_n522_), .B1(new_n472_), .B2(new_n471_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n520_), .A2(new_n235_), .A3(new_n462_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n521_), .A2(new_n480_), .A3(new_n523_), .A4(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n518_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(new_n444_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n513_), .A2(KEYINPUT20), .A3(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G226gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT19), .ZN(new_n530_));
  XOR2_X1   g329(.A(new_n530_), .B(KEYINPUT90), .Z(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n528_), .A2(new_n532_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n444_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n445_), .A2(new_n525_), .A3(new_n518_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n530_), .ZN(new_n536_));
  NAND4_X1  g335(.A1(new_n534_), .A2(KEYINPUT20), .A3(new_n535_), .A4(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G8gat), .B(G36gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT18), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(G92gat), .ZN(new_n541_));
  INV_X1    g340(.A(G64gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n539_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n257_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n533_), .A2(new_n537_), .A3(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n534_), .A2(KEYINPUT20), .A3(new_n535_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n530_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n513_), .A2(KEYINPUT20), .A3(new_n531_), .A4(new_n527_), .ZN(new_n549_));
  AND2_X1   g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  OAI211_X1 g349(.A(KEYINPUT27), .B(new_n546_), .C1(new_n550_), .C2(new_n545_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT99), .B(KEYINPUT27), .ZN(new_n552_));
  AND3_X1   g351(.A1(new_n533_), .A2(new_n537_), .A3(new_n545_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n545_), .B1(new_n533_), .B2(new_n537_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n552_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n509_), .A2(new_n556_), .ZN(new_n557_));
  NAND3_X1  g356(.A1(new_n541_), .A2(new_n544_), .A3(KEYINPUT32), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT98), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n558_), .A2(KEYINPUT96), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT96), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n541_), .A2(new_n544_), .A3(new_n563_), .A4(KEYINPUT32), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT97), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n533_), .A2(new_n565_), .A3(new_n566_), .A4(new_n537_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n533_), .A2(new_n537_), .A3(new_n565_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n568_), .A2(KEYINPUT97), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n409_), .A2(new_n567_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT33), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n408_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(KEYINPUT94), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT94), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n408_), .A2(new_n574_), .A3(new_n571_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n533_), .A2(new_n537_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n545_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT95), .ZN(new_n580_));
  INV_X1    g379(.A(new_n393_), .ZN(new_n581_));
  OAI21_X1  g380(.A(new_n580_), .B1(new_n581_), .B2(new_n396_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n399_), .A2(KEYINPUT95), .A3(new_n393_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n343_), .A3(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n342_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n584_), .A2(new_n406_), .A3(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n398_), .A2(new_n400_), .A3(KEYINPUT33), .A4(new_n405_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n579_), .A2(new_n586_), .A3(new_n546_), .A4(new_n587_), .ZN(new_n588_));
  OAI22_X1  g387(.A1(new_n561_), .A2(new_n570_), .B1(new_n576_), .B2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n454_), .A2(new_n506_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n502_), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n410_), .A2(new_n557_), .B1(new_n589_), .B2(new_n593_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n341_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT74), .ZN(new_n596_));
  NAND2_X1  g395(.A1(G232gat), .A2(G233gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n597_), .B(KEYINPUT34), .ZN(new_n598_));
  XNOR2_X1  g397(.A(KEYINPUT72), .B(KEYINPUT35), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n274_), .A2(KEYINPUT68), .A3(new_n277_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n307_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n225_), .B1(new_n604_), .B2(new_n303_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n214_), .ZN(new_n606_));
  OAI211_X1 g405(.A(new_n303_), .B(new_n606_), .C1(new_n306_), .C2(new_n305_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n601_), .B1(new_n605_), .B2(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n598_), .A2(new_n599_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n601_), .A2(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(new_n263_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n612_));
  OAI211_X1 g411(.A(new_n607_), .B(new_n611_), .C1(new_n612_), .C2(new_n225_), .ZN(new_n613_));
  AOI21_X1  g412(.A(new_n596_), .B1(new_n609_), .B2(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n613_), .A2(new_n596_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n614_), .A2(KEYINPUT73), .A3(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G190gat), .B(G218gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(G134gat), .ZN(new_n618_));
  INV_X1    g417(.A(G162gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(KEYINPUT36), .B1(new_n616_), .B2(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n608_), .B1(new_n310_), .B2(new_n226_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n613_), .B1(new_n623_), .B2(new_n600_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT74), .ZN(new_n625_));
  INV_X1    g424(.A(new_n615_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(new_n626_), .A3(new_n621_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT73), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n625_), .A2(new_n628_), .A3(new_n626_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT36), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n630_), .A3(new_n620_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n622_), .A2(new_n627_), .A3(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n632_), .A2(KEYINPUT37), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT37), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n622_), .A2(new_n631_), .A3(new_n634_), .A4(new_n627_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n633_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n297_), .B(new_n221_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n637_), .B(new_n638_), .Z(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT75), .ZN(new_n640_));
  XNOR2_X1  g439(.A(G127gat), .B(G155gat), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT16), .ZN(new_n642_));
  INV_X1    g441(.A(G183gat), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n642_), .B(new_n643_), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n644_), .B(G211gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n646_), .A2(KEYINPUT17), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n640_), .B(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n639_), .A2(KEYINPUT17), .A3(new_n646_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n636_), .A2(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n595_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n652_), .A2(new_n216_), .A3(new_n409_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT38), .ZN(new_n654_));
  OR3_X1    g453(.A1(new_n341_), .A2(KEYINPUT100), .A3(new_n650_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n594_), .A2(new_n632_), .ZN(new_n656_));
  OAI21_X1  g455(.A(KEYINPUT100), .B1(new_n341_), .B2(new_n650_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n655_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G1gat), .B1(new_n658_), .B2(new_n410_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n654_), .A2(new_n659_), .ZN(G1324gat));
  NAND3_X1  g459(.A1(new_n652_), .A2(new_n217_), .A3(new_n556_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT39), .ZN(new_n662_));
  INV_X1    g461(.A(new_n658_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(new_n556_), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n662_), .B1(new_n664_), .B2(G8gat), .ZN(new_n665_));
  AOI211_X1 g464(.A(KEYINPUT39), .B(new_n217_), .C1(new_n663_), .C2(new_n556_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n661_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g467(.A(G15gat), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n652_), .A2(new_n669_), .A3(new_n592_), .ZN(new_n670_));
  OAI21_X1  g469(.A(G15gat), .B1(new_n658_), .B2(new_n502_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT41), .ZN(new_n672_));
  AND2_X1   g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n671_), .A2(new_n672_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n670_), .B1(new_n673_), .B2(new_n674_), .ZN(G1326gat));
  NAND3_X1  g474(.A1(new_n652_), .A2(new_n418_), .A3(new_n591_), .ZN(new_n676_));
  OAI21_X1  g475(.A(G22gat), .B1(new_n658_), .B2(new_n590_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n677_), .A2(new_n678_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n676_), .B1(new_n679_), .B2(new_n680_), .ZN(G1327gat));
  NAND2_X1  g480(.A1(new_n589_), .A2(new_n593_), .ZN(new_n682_));
  AND2_X1   g481(.A1(new_n551_), .A2(new_n555_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n683_), .B(new_n410_), .C1(new_n507_), .C2(new_n508_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n685_), .A2(new_n636_), .A3(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n686_), .B1(new_n685_), .B2(new_n636_), .ZN(new_n688_));
  OAI211_X1 g487(.A(new_n340_), .B(new_n650_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  AND2_X1   g490(.A1(new_n633_), .A2(new_n635_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT43), .B1(new_n692_), .B2(new_n594_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n685_), .A2(new_n636_), .A3(new_n686_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  NAND4_X1  g494(.A1(new_n695_), .A2(KEYINPUT44), .A3(new_n340_), .A4(new_n650_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n691_), .A2(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G29gat), .B1(new_n697_), .B2(new_n410_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n650_), .ZN(new_n699_));
  INV_X1    g498(.A(new_n632_), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n595_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n702_), .A2(new_n203_), .A3(new_n409_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n698_), .A2(new_n703_), .ZN(G1328gat));
  NAND3_X1  g503(.A1(new_n702_), .A2(new_n204_), .A3(new_n556_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT45), .ZN(new_n706_));
  OAI21_X1  g505(.A(G36gat), .B1(new_n697_), .B2(new_n683_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT102), .B1(new_n706_), .B2(new_n707_), .ZN(new_n708_));
  XOR2_X1   g507(.A(new_n708_), .B(KEYINPUT46), .Z(G1329gat));
  INV_X1    g508(.A(KEYINPUT47), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n340_), .A2(new_n592_), .A3(new_n685_), .A4(new_n701_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(new_n206_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT104), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n691_), .A2(new_n696_), .A3(G43gat), .A4(new_n592_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n714_), .A2(KEYINPUT103), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n714_), .A2(KEYINPUT103), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n713_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(KEYINPUT106), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT105), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n714_), .B(KEYINPUT103), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n721_), .A3(new_n713_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n718_), .A2(new_n719_), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n719_), .B1(new_n718_), .B2(new_n722_), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n710_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  NOR2_X1   g524(.A1(new_n717_), .A2(KEYINPUT106), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n721_), .B1(new_n720_), .B2(new_n713_), .ZN(new_n727_));
  OAI21_X1  g526(.A(KEYINPUT105), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n718_), .A2(new_n719_), .A3(new_n722_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n728_), .A2(KEYINPUT47), .A3(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n725_), .A2(new_n730_), .ZN(G1330gat));
  OAI21_X1  g530(.A(G50gat), .B1(new_n697_), .B2(new_n590_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n702_), .A2(new_n202_), .A3(new_n591_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1331gat));
  NAND2_X1  g533(.A1(new_n335_), .A2(new_n339_), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n735_), .A2(new_n241_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n736_), .A2(new_n656_), .A3(new_n699_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n737_), .A2(G57gat), .A3(new_n409_), .ZN(new_n738_));
  XOR2_X1   g537(.A(new_n738_), .B(KEYINPUT108), .Z(new_n739_));
  NOR3_X1   g538(.A1(new_n735_), .A2(new_n594_), .A3(new_n241_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(new_n651_), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n741_), .A2(KEYINPUT107), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n410_), .B1(new_n741_), .B2(KEYINPUT107), .ZN(new_n743_));
  AOI21_X1  g542(.A(G57gat), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n739_), .A2(new_n744_), .ZN(G1332gat));
  AOI21_X1  g544(.A(new_n542_), .B1(new_n737_), .B2(new_n556_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT48), .Z(new_n747_));
  INV_X1    g546(.A(new_n741_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n748_), .A2(new_n542_), .A3(new_n556_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n747_), .A2(new_n749_), .ZN(G1333gat));
  AOI21_X1  g549(.A(new_n283_), .B1(new_n737_), .B2(new_n592_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT49), .Z(new_n752_));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n283_), .A3(new_n592_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(G1334gat));
  AOI21_X1  g553(.A(new_n281_), .B1(new_n737_), .B2(new_n591_), .ZN(new_n755_));
  XOR2_X1   g554(.A(new_n755_), .B(KEYINPUT50), .Z(new_n756_));
  NAND3_X1  g555(.A1(new_n748_), .A2(new_n281_), .A3(new_n591_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(G1335gat));
  NAND2_X1  g557(.A1(new_n740_), .A2(new_n701_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n256_), .B1(new_n759_), .B2(new_n410_), .ZN(new_n760_));
  XOR2_X1   g559(.A(new_n760_), .B(KEYINPUT109), .Z(new_n761_));
  AND3_X1   g560(.A1(new_n695_), .A2(new_n650_), .A3(new_n736_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT110), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT110), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n410_), .A2(new_n256_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n761_), .B1(new_n765_), .B2(new_n766_), .ZN(G1336gat));
  OAI21_X1  g566(.A(new_n257_), .B1(new_n759_), .B2(new_n683_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT111), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n683_), .A2(new_n257_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n769_), .B1(new_n765_), .B2(new_n770_), .ZN(G1337gat));
  NAND3_X1  g570(.A1(new_n763_), .A2(new_n592_), .A3(new_n764_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n772_), .A2(G99gat), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n740_), .A2(new_n244_), .A3(new_n592_), .A4(new_n701_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(KEYINPUT112), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n773_), .A2(new_n777_), .A3(new_n774_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n779_), .B(KEYINPUT51), .ZN(G1338gat));
  AOI21_X1  g579(.A(new_n245_), .B1(new_n762_), .B2(new_n591_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  XNOR2_X1  g581(.A(new_n781_), .B(new_n782_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n759_), .A2(G106gat), .A3(new_n590_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT113), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n783_), .A2(new_n788_), .A3(new_n785_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT53), .ZN(new_n791_));
  XNOR2_X1  g590(.A(new_n790_), .B(new_n791_), .ZN(G1339gat));
  NAND2_X1  g591(.A1(new_n311_), .A2(KEYINPUT12), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n298_), .B(new_n299_), .C1(new_n612_), .C2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(KEYINPUT115), .B1(new_n794_), .B2(new_n316_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796_));
  AOI21_X1  g595(.A(new_n796_), .B1(new_n794_), .B2(new_n316_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n300_), .A2(new_n312_), .A3(new_n798_), .A4(new_n302_), .ZN(new_n799_));
  AND3_X1   g598(.A1(new_n795_), .A2(new_n797_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n794_), .A2(new_n316_), .ZN(new_n801_));
  AOI22_X1  g600(.A1(new_n795_), .A2(new_n799_), .B1(new_n801_), .B2(KEYINPUT55), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n322_), .B1(new_n800_), .B2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT56), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT56), .ZN(new_n805_));
  OAI211_X1 g604(.A(new_n805_), .B(new_n322_), .C1(new_n800_), .C2(new_n802_), .ZN(new_n806_));
  NAND4_X1  g605(.A1(new_n804_), .A2(new_n241_), .A3(new_n325_), .A4(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n227_), .A2(new_n231_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n230_), .A2(new_n228_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n808_), .A2(new_n238_), .A3(new_n809_), .ZN(new_n810_));
  AND2_X1   g609(.A1(new_n239_), .A2(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n328_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n807_), .A2(new_n812_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT57), .B1(new_n813_), .B2(new_n700_), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n814_), .A2(KEYINPUT116), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(KEYINPUT116), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n804_), .A2(new_n325_), .A3(new_n811_), .A4(new_n806_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n818_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n819_), .A2(new_n636_), .A3(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n813_), .A2(KEYINPUT57), .A3(new_n700_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n815_), .A2(new_n816_), .A3(new_n821_), .A4(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n650_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT114), .B1(new_n699_), .B2(new_n242_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n826_));
  NOR3_X1   g625(.A1(new_n650_), .A2(new_n826_), .A3(new_n241_), .ZN(new_n827_));
  OAI221_X1 g626(.A(new_n692_), .B1(new_n334_), .B2(new_n332_), .C1(new_n825_), .C2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT54), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n824_), .A2(new_n829_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n556_), .A2(new_n410_), .ZN(new_n831_));
  AND2_X1   g630(.A1(new_n831_), .A2(new_n508_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(G113gat), .B1(new_n834_), .B2(new_n241_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n833_), .A2(KEYINPUT59), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n817_), .B(KEYINPUT58), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n814_), .B1(new_n636_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n813_), .A2(new_n700_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT57), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n821_), .A2(new_n843_), .A3(new_n839_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n822_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n650_), .B1(new_n840_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n829_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT59), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n848_), .A3(new_n832_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n836_), .A2(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n242_), .A2(new_n380_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n835_), .B1(new_n851_), .B2(new_n852_), .ZN(G1340gat));
  INV_X1    g652(.A(new_n735_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n851_), .A2(KEYINPUT118), .A3(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT118), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n856_), .B1(new_n850_), .B2(new_n735_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n855_), .A2(G120gat), .A3(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(G120gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(new_n735_), .B2(KEYINPUT60), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n834_), .B(new_n860_), .C1(KEYINPUT60), .C2(new_n859_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n861_), .ZN(G1341gat));
  AOI21_X1  g661(.A(G127gat), .B1(new_n834_), .B2(new_n699_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(KEYINPUT119), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n851_), .A2(G127gat), .A3(new_n699_), .ZN(new_n865_));
  AND2_X1   g664(.A1(new_n864_), .A2(new_n865_), .ZN(G1342gat));
  AOI21_X1  g665(.A(G134gat), .B1(new_n834_), .B2(new_n632_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n636_), .A2(G134gat), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n867_), .B1(new_n851_), .B2(new_n868_), .ZN(G1343gat));
  AND2_X1   g668(.A1(new_n830_), .A2(new_n507_), .ZN(new_n870_));
  AND2_X1   g669(.A1(new_n870_), .A2(new_n831_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n241_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g672(.A1(new_n871_), .A2(new_n854_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g674(.A1(new_n871_), .A2(new_n699_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT61), .B(G155gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n876_), .B(new_n877_), .ZN(G1346gat));
  AOI21_X1  g677(.A(G162gat), .B1(new_n871_), .B2(new_n632_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n692_), .A2(new_n619_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n871_), .B2(new_n880_), .ZN(G1347gat));
  NOR2_X1   g680(.A1(new_n683_), .A2(new_n409_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n508_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n822_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n885_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n821_), .A2(new_n843_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(KEYINPUT117), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n699_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n828_), .B(new_n890_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n241_), .B(new_n884_), .C1(new_n889_), .C2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n892_), .A2(KEYINPUT120), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT120), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n847_), .A2(new_n894_), .A3(new_n241_), .A4(new_n884_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n893_), .A2(G169gat), .A3(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n883_), .B1(new_n846_), .B2(new_n829_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n899_), .A2(new_n486_), .A3(new_n241_), .ZN(new_n900_));
  NAND4_X1  g699(.A1(new_n893_), .A2(KEYINPUT62), .A3(new_n895_), .A4(G169gat), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n898_), .A2(new_n900_), .A3(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  NAND4_X1  g703(.A1(new_n898_), .A2(KEYINPUT121), .A3(new_n900_), .A4(new_n901_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1348gat));
  AOI21_X1  g705(.A(G176gat), .B1(new_n899_), .B2(new_n854_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(KEYINPUT122), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n891_), .B1(new_n823_), .B2(new_n650_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n909_), .B1(new_n910_), .B2(new_n591_), .ZN(new_n911_));
  NAND3_X1  g710(.A1(new_n830_), .A2(KEYINPUT123), .A3(new_n590_), .ZN(new_n912_));
  NAND4_X1  g711(.A1(new_n911_), .A2(new_n912_), .A3(new_n592_), .A4(new_n882_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n913_), .A2(new_n462_), .A3(new_n735_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n908_), .A2(new_n914_), .ZN(G1349gat));
  AND2_X1   g714(.A1(new_n911_), .A2(new_n882_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n912_), .A2(new_n592_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT124), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n916_), .A2(new_n917_), .A3(new_n918_), .A4(new_n699_), .ZN(new_n919_));
  OAI21_X1  g718(.A(KEYINPUT124), .B1(new_n913_), .B2(new_n650_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n919_), .A2(new_n920_), .A3(new_n643_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n899_), .A2(new_n473_), .A3(new_n699_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1350gat));
  NAND3_X1  g722(.A1(new_n899_), .A2(new_n632_), .A3(new_n522_), .ZN(new_n924_));
  AND2_X1   g723(.A1(new_n899_), .A2(new_n636_), .ZN(new_n925_));
  INV_X1    g724(.A(G190gat), .ZN(new_n926_));
  OAI21_X1  g725(.A(new_n924_), .B1(new_n925_), .B2(new_n926_), .ZN(G1351gat));
  AND2_X1   g726(.A1(new_n870_), .A2(new_n882_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n928_), .A2(new_n241_), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n929_), .B(G197gat), .ZN(G1352gat));
  AND3_X1   g729(.A1(new_n870_), .A2(new_n854_), .A3(new_n882_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n437_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n933_), .B1(new_n931_), .B2(new_n321_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(KEYINPUT125), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT125), .ZN(new_n936_));
  OAI211_X1 g735(.A(new_n933_), .B(new_n936_), .C1(new_n321_), .C2(new_n931_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n937_), .ZN(G1353gat));
  AOI21_X1  g737(.A(new_n650_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n939_));
  OR2_X1    g738(.A1(new_n939_), .A2(KEYINPUT126), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(KEYINPUT126), .ZN(new_n941_));
  NAND3_X1  g740(.A1(new_n928_), .A2(new_n940_), .A3(new_n941_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n943_));
  XOR2_X1   g742(.A(new_n942_), .B(new_n943_), .Z(G1354gat));
  AOI21_X1  g743(.A(G218gat), .B1(new_n928_), .B2(new_n632_), .ZN(new_n945_));
  NAND2_X1  g744(.A1(new_n636_), .A2(G218gat), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(KEYINPUT127), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n945_), .B1(new_n928_), .B2(new_n947_), .ZN(G1355gat));
endmodule


