//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n738_, new_n739_, new_n740_, new_n742_, new_n743_,
    new_n744_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n835_, new_n836_, new_n838_, new_n839_,
    new_n840_, new_n842_, new_n844_, new_n845_, new_n847_, new_n848_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n857_, new_n858_, new_n859_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n888_, new_n889_;
  INV_X1    g000(.A(G106gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G211gat), .B(G218gat), .Z(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G197gat), .ZN(new_n205_));
  AND3_X1   g004(.A1(new_n205_), .A2(KEYINPUT90), .A3(G204gat), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT90), .B1(new_n205_), .B2(G204gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT89), .ZN(new_n210_));
  INV_X1    g009(.A(G204gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT88), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT88), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(G204gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n210_), .B1(new_n215_), .B2(G197gat), .ZN(new_n216_));
  AOI211_X1 g015(.A(KEYINPUT89), .B(new_n205_), .C1(new_n212_), .C2(new_n214_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n209_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n204_), .B1(new_n218_), .B2(KEYINPUT91), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT21), .ZN(new_n220_));
  XNOR2_X1  g019(.A(KEYINPUT88), .B(G204gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT89), .B1(new_n221_), .B2(new_n205_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(new_n213_), .A2(G204gat), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n211_), .A2(KEYINPUT88), .ZN(new_n224_));
  OAI211_X1 g023(.A(new_n210_), .B(G197gat), .C1(new_n223_), .C2(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n208_), .B1(new_n222_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT91), .ZN(new_n227_));
  AOI21_X1  g026(.A(new_n220_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n203_), .B1(new_n226_), .B2(new_n220_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G197gat), .A2(G204gat), .ZN(new_n230_));
  OAI211_X1 g029(.A(KEYINPUT21), .B(new_n230_), .C1(new_n221_), .C2(G197gat), .ZN(new_n231_));
  AOI22_X1  g030(.A1(new_n219_), .A2(new_n228_), .B1(new_n229_), .B2(new_n231_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(KEYINPUT84), .A2(KEYINPUT3), .ZN(new_n233_));
  INV_X1    g032(.A(G141gat), .ZN(new_n234_));
  INV_X1    g033(.A(G148gat), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n233_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G141gat), .A2(G148gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT2), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n240_));
  OAI22_X1  g039(.A1(KEYINPUT84), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n236_), .A2(new_n239_), .A3(new_n240_), .A4(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G155gat), .B(G162gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n246_));
  AND2_X1   g045(.A1(new_n246_), .A2(new_n237_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n234_), .A2(new_n235_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n247_), .B(new_n248_), .C1(new_n243_), .C2(KEYINPUT1), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n245_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(KEYINPUT93), .B(KEYINPUT29), .Z(new_n252_));
  NOR2_X1   g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  OAI211_X1 g052(.A(G228gat), .B(G233gat), .C1(new_n232_), .C2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G78gat), .ZN(new_n255_));
  OAI211_X1 g054(.A(new_n220_), .B(new_n209_), .C1(new_n216_), .C2(new_n217_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n256_), .A2(new_n231_), .A3(new_n204_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n227_), .B(new_n209_), .C1(new_n216_), .C2(new_n217_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT21), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n203_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n257_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT92), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n250_), .A2(KEYINPUT29), .B1(G228gat), .B2(G233gat), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n261_), .A2(new_n262_), .A3(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n262_), .B1(new_n261_), .B2(new_n263_), .ZN(new_n266_));
  OAI211_X1 g065(.A(new_n254_), .B(new_n255_), .C1(new_n265_), .C2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n263_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT92), .B1(new_n232_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n264_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n255_), .B1(new_n271_), .B2(new_n254_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n202_), .B1(new_n268_), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n254_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(G78gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n275_), .A2(G106gat), .A3(new_n267_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n273_), .A2(KEYINPUT87), .A3(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n250_), .A2(KEYINPUT29), .ZN(new_n278_));
  INV_X1    g077(.A(G50gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n278_), .B(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT85), .B(G22gat), .ZN(new_n281_));
  XNOR2_X1  g080(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n281_), .B(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n280_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n277_), .A2(new_n285_), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n273_), .A2(new_n276_), .A3(KEYINPUT87), .A4(new_n284_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G127gat), .B(G134gat), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G113gat), .B(G120gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n292_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n290_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n296_), .B(KEYINPUT31), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G71gat), .B(G99gat), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G227gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G15gat), .B(G43gat), .Z(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  INV_X1    g101(.A(KEYINPUT23), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n303_), .A2(G183gat), .A3(G190gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305_));
  AND3_X1   g104(.A1(new_n305_), .A2(KEYINPUT77), .A3(KEYINPUT23), .ZN(new_n306_));
  AOI21_X1  g105(.A(KEYINPUT77), .B1(new_n305_), .B2(KEYINPUT23), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n304_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(G169gat), .A2(G176gat), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n310_), .A2(G169gat), .A3(G176gat), .ZN(new_n311_));
  INV_X1    g110(.A(G169gat), .ZN(new_n312_));
  INV_X1    g111(.A(G176gat), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT76), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  OAI211_X1 g113(.A(KEYINPUT24), .B(new_n309_), .C1(new_n311_), .C2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT25), .B(G183gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G190gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n312_), .A2(new_n313_), .A3(KEYINPUT76), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n310_), .B1(G169gat), .B2(G176gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n319_), .A2(new_n320_), .A3(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n308_), .A2(new_n315_), .A3(new_n318_), .A4(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n324_));
  NOR2_X1   g123(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n313_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT78), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n305_), .A2(KEYINPUT23), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(new_n304_), .ZN(new_n330_));
  OR2_X1    g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT22), .B(G169gat), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n333_), .A2(KEYINPUT78), .A3(new_n313_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n328_), .A2(new_n332_), .A3(new_n334_), .A4(new_n309_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n323_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT30), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n336_), .B(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n336_), .B(KEYINPUT30), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(new_n339_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n302_), .B1(new_n341_), .B2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n341_), .A2(new_n343_), .A3(new_n302_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(KEYINPUT81), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n348_));
  AOI21_X1  g147(.A(new_n297_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n346_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(new_n344_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT81), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(new_n297_), .B2(new_n348_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n349_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n289_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n250_), .A2(new_n296_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT98), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n245_), .A2(new_n249_), .A3(new_n293_), .A4(new_n295_), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n357_), .A2(new_n358_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(G225gat), .A2(G233gat), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n250_), .A2(KEYINPUT98), .A3(new_n296_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT99), .B(KEYINPUT4), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n357_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n360_), .A2(new_n362_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n365_), .B1(new_n366_), .B2(KEYINPUT4), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n363_), .B1(new_n367_), .B2(new_n361_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G1gat), .B(G29gat), .ZN(new_n369_));
  INV_X1    g168(.A(G85gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT0), .B(G57gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n368_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n373_), .ZN(new_n375_));
  OAI211_X1 g174(.A(new_n363_), .B(new_n375_), .C1(new_n367_), .C2(new_n361_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n374_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT27), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n261_), .A2(new_n336_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n380_), .B(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n316_), .A2(KEYINPUT96), .ZN(new_n384_));
  NOR2_X1   g183(.A1(new_n316_), .A2(KEYINPUT96), .ZN(new_n385_));
  OAI21_X1  g184(.A(new_n317_), .B1(new_n384_), .B2(new_n385_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n321_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n386_), .A2(new_n315_), .A3(new_n330_), .A4(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n308_), .A2(new_n331_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n389_), .A2(new_n309_), .A3(new_n326_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT20), .B1(new_n261_), .B2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n383_), .A2(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n323_), .A2(new_n335_), .ZN(new_n395_));
  OAI211_X1 g194(.A(new_n395_), .B(new_n257_), .C1(new_n259_), .C2(new_n260_), .ZN(new_n396_));
  AND3_X1   g195(.A1(new_n396_), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n397_));
  AOI21_X1  g196(.A(KEYINPUT95), .B1(new_n396_), .B2(KEYINPUT20), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n261_), .A2(new_n391_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR3_X1   g199(.A1(new_n397_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n394_), .B1(new_n401_), .B2(new_n382_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(KEYINPUT97), .B(KEYINPUT18), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G64gat), .B(G92gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406_));
  XOR2_X1   g205(.A(new_n405_), .B(new_n406_), .Z(new_n407_));
  NAND2_X1  g206(.A1(new_n402_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n396_), .A2(KEYINPUT20), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT95), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n396_), .A2(KEYINPUT95), .A3(KEYINPUT20), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n411_), .A2(new_n399_), .A3(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n382_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n393_), .B1(new_n413_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n407_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n408_), .A2(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(new_n397_), .A2(new_n398_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT102), .ZN(new_n420_));
  NAND4_X1  g219(.A1(new_n419_), .A2(new_n420_), .A3(new_n382_), .A4(new_n399_), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n411_), .A2(new_n382_), .A3(new_n399_), .A4(new_n412_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(KEYINPUT102), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT101), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n392_), .A2(new_n424_), .ZN(new_n425_));
  OAI211_X1 g224(.A(KEYINPUT101), .B(KEYINPUT20), .C1(new_n261_), .C2(new_n391_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n425_), .A2(new_n426_), .A3(new_n379_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n414_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n421_), .A2(new_n423_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(new_n407_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n378_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n431_));
  AOI22_X1  g230(.A1(new_n378_), .A2(new_n418_), .B1(new_n430_), .B2(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NOR3_X1   g232(.A1(new_n356_), .A2(new_n377_), .A3(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT103), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT100), .B(KEYINPUT33), .Z(new_n436_));
  NAND3_X1  g235(.A1(new_n366_), .A2(G225gat), .A3(G233gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n373_), .B1(new_n367_), .B2(new_n361_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n374_), .A2(new_n436_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT100), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n368_), .B(new_n373_), .C1(new_n440_), .C2(KEYINPUT33), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n408_), .A2(new_n417_), .A3(new_n439_), .A4(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n416_), .A2(KEYINPUT32), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n429_), .A2(new_n444_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n394_), .B(new_n443_), .C1(new_n401_), .C2(new_n382_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(new_n377_), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n442_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n377_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n289_), .A2(new_n448_), .B1(new_n449_), .B2(new_n432_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n347_), .A2(new_n348_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n297_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(new_n354_), .ZN(new_n454_));
  AOI21_X1  g253(.A(KEYINPUT83), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n349_), .A2(new_n354_), .A3(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n455_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n435_), .B1(new_n450_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n377_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n288_), .A2(new_n432_), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n442_), .ZN(new_n462_));
  AOI21_X1  g261(.A(new_n447_), .B1(new_n444_), .B2(new_n429_), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n287_), .B(new_n286_), .C1(new_n462_), .C2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n458_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n465_), .A2(KEYINPUT103), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n434_), .B1(new_n459_), .B2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G57gat), .B(G64gat), .ZN(new_n469_));
  AND2_X1   g268(.A1(new_n469_), .A2(KEYINPUT11), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(KEYINPUT11), .ZN(new_n471_));
  XNOR2_X1  g270(.A(G71gat), .B(G78gat), .ZN(new_n472_));
  OR3_X1    g271(.A1(new_n470_), .A2(new_n471_), .A3(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n469_), .A2(new_n472_), .A3(KEYINPUT11), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G15gat), .B(G22gat), .ZN(new_n476_));
  INV_X1    g275(.A(G1gat), .ZN(new_n477_));
  INV_X1    g276(.A(G8gat), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT14), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n476_), .A2(new_n479_), .ZN(new_n480_));
  XNOR2_X1  g279(.A(G1gat), .B(G8gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XOR2_X1   g281(.A(new_n475_), .B(new_n482_), .Z(new_n483_));
  NAND2_X1  g282(.A1(G231gat), .A2(G233gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G183gat), .B(G211gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(KEYINPUT75), .B(KEYINPUT16), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G127gat), .B(G155gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  XOR2_X1   g289(.A(new_n490_), .B(KEYINPUT17), .Z(new_n491_));
  OR2_X1    g290(.A1(new_n485_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n490_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n485_), .A2(KEYINPUT17), .A3(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n492_), .A2(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G190gat), .B(G218gat), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G134gat), .B(G162gat), .ZN(new_n498_));
  XOR2_X1   g297(.A(new_n497_), .B(new_n498_), .Z(new_n499_));
  XNOR2_X1  g298(.A(KEYINPUT10), .B(G99gat), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT65), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n500_), .B(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(new_n202_), .ZN(new_n503_));
  INV_X1    g302(.A(G92gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n370_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(KEYINPUT66), .A3(KEYINPUT9), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n507_));
  INV_X1    g306(.A(G99gat), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n507_), .B1(new_n508_), .B2(new_n202_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G85gat), .B(G92gat), .ZN(new_n513_));
  AOI21_X1  g312(.A(KEYINPUT66), .B1(new_n513_), .B2(KEYINPUT9), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n514_), .B1(KEYINPUT9), .B2(new_n505_), .ZN(new_n515_));
  NAND4_X1  g314(.A1(new_n503_), .A2(new_n506_), .A3(new_n512_), .A4(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT67), .ZN(new_n517_));
  AND2_X1   g316(.A1(new_n515_), .A2(new_n512_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT67), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n518_), .A2(new_n503_), .A3(new_n519_), .A4(new_n506_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n513_), .B(KEYINPUT69), .Z(new_n522_));
  INV_X1    g321(.A(KEYINPUT70), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n511_), .B(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n508_), .A2(new_n202_), .ZN(new_n525_));
  AND2_X1   g324(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n526_));
  NOR2_X1   g325(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n528_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n522_), .B1(new_n524_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n530_), .A2(KEYINPUT8), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT8), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n522_), .B(new_n532_), .C1(new_n511_), .C2(new_n529_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n531_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n521_), .A2(new_n534_), .ZN(new_n535_));
  XOR2_X1   g334(.A(G43gat), .B(G50gat), .Z(new_n536_));
  XNOR2_X1  g335(.A(G29gat), .B(G36gat), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n537_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  OAI21_X1  g339(.A(KEYINPUT74), .B1(new_n535_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT73), .ZN(new_n542_));
  AOI22_X1  g341(.A1(new_n517_), .A2(new_n520_), .B1(new_n531_), .B2(new_n533_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(new_n538_), .A4(new_n539_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n541_), .A2(new_n542_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(G232gat), .A2(G233gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(KEYINPUT34), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n546_), .A2(KEYINPUT35), .A3(new_n548_), .ZN(new_n549_));
  XOR2_X1   g348(.A(new_n540_), .B(KEYINPUT15), .Z(new_n550_));
  NAND2_X1  g349(.A1(new_n535_), .A2(new_n550_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n541_), .A2(new_n545_), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n549_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  OR2_X1    g353(.A1(new_n548_), .A2(KEYINPUT35), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n552_), .B1(new_n549_), .B2(new_n555_), .ZN(new_n556_));
  OAI211_X1 g355(.A(new_n496_), .B(new_n499_), .C1(new_n554_), .C2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n549_), .A2(new_n555_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n552_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n499_), .A2(new_n496_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n499_), .A2(new_n496_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .A4(new_n553_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n557_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT37), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  NAND3_X1  g365(.A1(new_n557_), .A2(new_n563_), .A3(KEYINPUT37), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NOR3_X1   g367(.A1(new_n468_), .A2(new_n495_), .A3(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n475_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n535_), .A2(new_n570_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n543_), .A2(new_n475_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(KEYINPUT12), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n475_), .B1(new_n521_), .B2(new_n534_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT12), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G230gat), .A2(G233gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n578_), .B(KEYINPUT64), .Z(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n577_), .A2(new_n580_), .ZN(new_n581_));
  AND3_X1   g380(.A1(new_n521_), .A2(new_n534_), .A3(new_n475_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n579_), .B1(new_n582_), .B2(new_n574_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G120gat), .B(G148gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(G204gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT5), .B(G176gat), .ZN(new_n587_));
  XOR2_X1   g386(.A(new_n586_), .B(new_n587_), .Z(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n589_), .A2(KEYINPUT71), .ZN(new_n590_));
  XOR2_X1   g389(.A(new_n590_), .B(KEYINPUT72), .Z(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n584_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n581_), .A2(new_n583_), .A3(new_n591_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT13), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n593_), .A2(KEYINPUT13), .A3(new_n594_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n482_), .B(new_n540_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n482_), .A2(new_n540_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n601_), .B1(new_n550_), .B2(new_n482_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(G229gat), .A2(G233gat), .ZN(new_n603_));
  MUX2_X1   g402(.A(new_n600_), .B(new_n602_), .S(new_n603_), .Z(new_n604_));
  XNOR2_X1  g403(.A(G113gat), .B(G141gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G169gat), .B(G197gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n604_), .B(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n599_), .A2(new_n609_), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n569_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n377_), .B(KEYINPUT104), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n611_), .A2(new_n477_), .A3(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT38), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n616_), .A2(KEYINPUT105), .ZN(new_n617_));
  INV_X1    g416(.A(new_n564_), .ZN(new_n618_));
  NOR3_X1   g417(.A1(new_n468_), .A2(new_n495_), .A3(new_n618_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n619_), .A2(new_n610_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n477_), .B1(new_n620_), .B2(new_n377_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n614_), .B1(new_n621_), .B2(new_n615_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n616_), .A2(KEYINPUT105), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n617_), .A2(new_n622_), .A3(new_n623_), .ZN(G1324gat));
  NAND3_X1  g423(.A1(new_n611_), .A2(new_n478_), .A3(new_n433_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n478_), .B1(new_n620_), .B2(new_n433_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT39), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n626_), .A2(new_n627_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n625_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT40), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(G1325gat));
  INV_X1    g432(.A(G15gat), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n634_), .B1(new_n620_), .B2(new_n458_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT41), .ZN(new_n636_));
  NAND3_X1  g435(.A1(new_n611_), .A2(new_n634_), .A3(new_n458_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(G1326gat));
  INV_X1    g437(.A(G22gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n611_), .A2(new_n639_), .A3(new_n288_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n620_), .B2(new_n288_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT106), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT42), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n642_), .ZN(new_n645_));
  AND3_X1   g444(.A1(new_n643_), .A2(new_n644_), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n640_), .B1(new_n646_), .B2(new_n647_), .ZN(G1327gat));
  NOR2_X1   g447(.A1(new_n468_), .A2(new_n564_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n495_), .ZN(new_n650_));
  NOR3_X1   g449(.A1(new_n599_), .A2(new_n609_), .A3(new_n650_), .ZN(new_n651_));
  AND2_X1   g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  OR3_X1    g452(.A1(new_n653_), .A2(G29gat), .A3(new_n460_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n568_), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n468_), .A2(KEYINPUT43), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT43), .ZN(new_n657_));
  INV_X1    g456(.A(new_n356_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n658_), .A2(new_n460_), .A3(new_n432_), .ZN(new_n659_));
  AOI21_X1  g458(.A(KEYINPUT103), .B1(new_n465_), .B2(new_n466_), .ZN(new_n660_));
  AOI211_X1 g459(.A(new_n435_), .B(new_n458_), .C1(new_n461_), .C2(new_n464_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n659_), .B1(new_n660_), .B2(new_n661_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n657_), .B1(new_n662_), .B2(new_n568_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n651_), .B1(new_n656_), .B2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT107), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n665_), .A2(KEYINPUT44), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n666_), .ZN(new_n668_));
  OAI211_X1 g467(.A(new_n651_), .B(new_n668_), .C1(new_n656_), .C2(new_n663_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n667_), .A2(new_n613_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT108), .ZN(new_n671_));
  AND3_X1   g470(.A1(new_n670_), .A2(new_n671_), .A3(G29gat), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n670_), .B2(G29gat), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n654_), .B1(new_n672_), .B2(new_n673_), .ZN(G1328gat));
  INV_X1    g473(.A(KEYINPUT110), .ZN(new_n675_));
  INV_X1    g474(.A(G36gat), .ZN(new_n676_));
  NAND4_X1  g475(.A1(new_n652_), .A2(new_n675_), .A3(new_n676_), .A4(new_n433_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n649_), .A2(new_n676_), .A3(new_n651_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT110), .B1(new_n678_), .B2(new_n432_), .ZN(new_n679_));
  XOR2_X1   g478(.A(KEYINPUT111), .B(KEYINPUT45), .Z(new_n680_));
  AND3_X1   g479(.A1(new_n677_), .A2(new_n679_), .A3(new_n680_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n667_), .A2(new_n433_), .A3(new_n669_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT109), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n684_), .A2(new_n685_), .A3(G36gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n684_), .B2(G36gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n683_), .B1(new_n686_), .B2(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT46), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(new_n690_));
  OAI211_X1 g489(.A(new_n683_), .B(KEYINPUT46), .C1(new_n686_), .C2(new_n687_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(G1329gat));
  INV_X1    g491(.A(G43gat), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n693_), .B1(new_n653_), .B2(new_n466_), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n667_), .A2(G43gat), .A3(new_n355_), .A4(new_n669_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n695_), .A2(KEYINPUT112), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n695_), .A2(KEYINPUT112), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n694_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  XNOR2_X1  g497(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n699_));
  INV_X1    g498(.A(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n700_), .ZN(new_n701_));
  OAI211_X1 g500(.A(new_n699_), .B(new_n694_), .C1(new_n696_), .C2(new_n697_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(G1330gat));
  NAND3_X1  g502(.A1(new_n652_), .A2(new_n279_), .A3(new_n288_), .ZN(new_n704_));
  AND3_X1   g503(.A1(new_n667_), .A2(new_n288_), .A3(new_n669_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n704_), .B1(new_n705_), .B2(new_n279_), .ZN(G1331gat));
  INV_X1    g505(.A(new_n599_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n707_), .A2(new_n608_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n619_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(G57gat), .ZN(new_n710_));
  NOR3_X1   g509(.A1(new_n709_), .A2(new_n710_), .A3(new_n460_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n569_), .A2(new_n708_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(new_n613_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n711_), .B1(new_n710_), .B2(new_n714_), .ZN(G1332gat));
  OAI21_X1  g514(.A(G64gat), .B1(new_n709_), .B2(new_n432_), .ZN(new_n716_));
  XOR2_X1   g515(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n717_));
  XNOR2_X1  g516(.A(new_n716_), .B(new_n717_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n432_), .A2(G64gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n718_), .B1(new_n712_), .B2(new_n719_), .ZN(G1333gat));
  OAI21_X1  g519(.A(G71gat), .B1(new_n709_), .B2(new_n466_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT49), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n466_), .A2(G71gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n712_), .B2(new_n723_), .ZN(G1334gat));
  OAI21_X1  g523(.A(G78gat), .B1(new_n709_), .B2(new_n289_), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n725_), .B(KEYINPUT50), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n713_), .A2(new_n255_), .A3(new_n288_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT115), .ZN(G1335gat));
  NOR3_X1   g528(.A1(new_n707_), .A2(new_n608_), .A3(new_n650_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n649_), .A2(new_n730_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT116), .Z(new_n732_));
  NOR2_X1   g531(.A1(new_n612_), .A2(G85gat), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n656_), .A2(new_n663_), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n734_), .A2(new_n377_), .A3(new_n730_), .ZN(new_n735_));
  AOI22_X1  g534(.A1(new_n732_), .A2(new_n733_), .B1(G85gat), .B2(new_n735_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT117), .Z(G1336gat));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n730_), .ZN(new_n738_));
  NOR3_X1   g537(.A1(new_n738_), .A2(new_n504_), .A3(new_n432_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n732_), .A2(new_n433_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n740_), .B2(new_n504_), .ZN(G1337gat));
  NAND3_X1  g540(.A1(new_n732_), .A2(new_n502_), .A3(new_n355_), .ZN(new_n742_));
  OAI21_X1  g541(.A(G99gat), .B1(new_n738_), .B2(new_n466_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n744_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g544(.A1(new_n732_), .A2(new_n202_), .A3(new_n288_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n734_), .A2(new_n288_), .A3(new_n730_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT52), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n747_), .A2(new_n748_), .A3(G106gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n747_), .B2(G106gat), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT53), .ZN(G1339gat));
  OR2_X1    g551(.A1(new_n604_), .A2(new_n607_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n600_), .A2(new_n603_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n602_), .ZN(new_n755_));
  OAI211_X1 g554(.A(new_n607_), .B(new_n754_), .C1(new_n755_), .C2(new_n603_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n753_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n581_), .A2(new_n583_), .A3(new_n589_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n577_), .A2(new_n580_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n543_), .A2(KEYINPUT12), .A3(new_n475_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n582_), .A2(new_n574_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(KEYINPUT12), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT55), .B1(new_n763_), .B2(new_n579_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT55), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n577_), .A2(new_n765_), .A3(new_n580_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n760_), .B1(new_n764_), .B2(new_n766_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT56), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n589_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n765_), .B1(new_n577_), .B2(new_n580_), .ZN(new_n770_));
  AOI211_X1 g569(.A(KEYINPUT55), .B(new_n579_), .C1(new_n573_), .C2(new_n576_), .ZN(new_n771_));
  OAI22_X1  g570(.A1(new_n770_), .A2(new_n771_), .B1(new_n580_), .B2(new_n577_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT56), .B1(new_n772_), .B2(new_n588_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n758_), .B(new_n759_), .C1(new_n769_), .C2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT58), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n768_), .B1(new_n767_), .B2(new_n589_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n772_), .A2(KEYINPUT56), .A3(new_n588_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n779_), .A2(KEYINPUT58), .A3(new_n758_), .A4(new_n759_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n776_), .A2(new_n568_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n759_), .A2(new_n608_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n782_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n757_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n564_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT57), .B(new_n564_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n781_), .A2(new_n787_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT119), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT119), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n781_), .A2(new_n787_), .A3(new_n791_), .A4(new_n788_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n790_), .A2(new_n495_), .A3(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n597_), .A2(new_n609_), .A3(new_n598_), .A4(new_n650_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n794_), .A2(new_n795_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n655_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  XNOR2_X1  g597(.A(new_n798_), .B(KEYINPUT54), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n793_), .A2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n433_), .A2(new_n612_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n658_), .A2(new_n801_), .ZN(new_n802_));
  XOR2_X1   g601(.A(new_n802_), .B(KEYINPUT120), .Z(new_n803_));
  NAND2_X1  g602(.A1(new_n800_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT121), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n800_), .A2(KEYINPUT121), .A3(new_n803_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(G113gat), .B1(new_n808_), .B2(new_n608_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n804_), .A2(KEYINPUT59), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n789_), .A2(new_n495_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT123), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT123), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n789_), .A2(new_n813_), .A3(new_n495_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n812_), .A2(new_n799_), .A3(new_n814_), .ZN(new_n815_));
  XOR2_X1   g614(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n803_), .A3(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n810_), .A2(new_n817_), .ZN(new_n818_));
  AND2_X1   g617(.A1(new_n608_), .A2(G113gat), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n809_), .B1(new_n818_), .B2(new_n819_), .ZN(G1340gat));
  INV_X1    g619(.A(G120gat), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT60), .B1(new_n599_), .B2(new_n821_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n822_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n810_), .A2(new_n599_), .A3(new_n817_), .ZN(new_n824_));
  OAI21_X1  g623(.A(G120gat), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n823_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n825_), .B1(KEYINPUT60), .B2(new_n826_), .ZN(G1341gat));
  NAND4_X1  g626(.A1(new_n810_), .A2(G127gat), .A3(new_n650_), .A4(new_n817_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n495_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n828_), .B1(new_n829_), .B2(G127gat), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(KEYINPUT124), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT124), .ZN(new_n832_));
  OAI211_X1 g631(.A(new_n832_), .B(new_n828_), .C1(new_n829_), .C2(G127gat), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n831_), .A2(new_n833_), .ZN(G1342gat));
  AOI21_X1  g633(.A(G134gat), .B1(new_n808_), .B2(new_n618_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n568_), .A2(G134gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n835_), .B1(new_n818_), .B2(new_n836_), .ZN(G1343gat));
  AND4_X1   g636(.A1(new_n466_), .A2(new_n800_), .A3(new_n288_), .A4(new_n801_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n608_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT125), .B(G141gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(G1344gat));
  NAND2_X1  g640(.A1(new_n838_), .A2(new_n599_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g642(.A1(new_n838_), .A2(new_n650_), .ZN(new_n844_));
  XNOR2_X1  g643(.A(KEYINPUT61), .B(G155gat), .ZN(new_n845_));
  XNOR2_X1  g644(.A(new_n844_), .B(new_n845_), .ZN(G1346gat));
  AOI21_X1  g645(.A(G162gat), .B1(new_n838_), .B2(new_n618_), .ZN(new_n847_));
  AND2_X1   g646(.A1(new_n568_), .A2(G162gat), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n847_), .B1(new_n838_), .B2(new_n848_), .ZN(G1347gat));
  NOR4_X1   g648(.A1(new_n466_), .A2(new_n288_), .A3(new_n432_), .A4(new_n613_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n815_), .A2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(G169gat), .B1(new_n851_), .B2(new_n609_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n851_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n608_), .A3(new_n333_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n852_), .ZN(new_n855_));
  MUX2_X1   g654(.A(new_n852_), .B(new_n855_), .S(KEYINPUT62), .Z(G1348gat));
  AOI21_X1  g655(.A(G176gat), .B1(new_n853_), .B2(new_n599_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n800_), .A2(new_n850_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n707_), .A2(new_n313_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n858_), .B2(new_n859_), .ZN(G1349gat));
  AOI21_X1  g659(.A(G183gat), .B1(new_n858_), .B2(new_n650_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n495_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n861_), .B1(new_n853_), .B2(new_n862_), .ZN(G1350gat));
  OAI21_X1  g662(.A(G190gat), .B1(new_n851_), .B2(new_n655_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n618_), .A2(new_n317_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n864_), .B1(new_n851_), .B2(new_n865_), .ZN(G1351gat));
  NOR3_X1   g665(.A1(new_n289_), .A2(new_n458_), .A3(new_n432_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n800_), .A2(new_n460_), .A3(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n868_), .A2(new_n609_), .ZN(new_n869_));
  XNOR2_X1  g668(.A(new_n869_), .B(new_n205_), .ZN(G1352gat));
  INV_X1    g669(.A(new_n868_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(new_n599_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(G204gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n221_), .B2(new_n872_), .ZN(G1353gat));
  INV_X1    g673(.A(KEYINPUT63), .ZN(new_n875_));
  INV_X1    g674(.A(G211gat), .ZN(new_n876_));
  OAI21_X1  g675(.A(new_n650_), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(KEYINPUT126), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n871_), .A2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(KEYINPUT127), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT127), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n871_), .A2(new_n881_), .A3(new_n878_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n875_), .A2(new_n876_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND4_X1  g684(.A1(new_n880_), .A2(new_n875_), .A3(new_n876_), .A4(new_n882_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1354gat));
  AND3_X1   g686(.A1(new_n871_), .A2(G218gat), .A3(new_n568_), .ZN(new_n888_));
  AOI21_X1  g687(.A(G218gat), .B1(new_n871_), .B2(new_n618_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1355gat));
endmodule


