//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 0 1 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n856_,
    new_n857_, new_n859_, new_n860_, new_n861_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n898_, new_n899_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_;
  AND2_X1   g000(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n202_));
  NOR2_X1   g001(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(G176gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(KEYINPUT80), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n208_));
  INV_X1    g007(.A(G183gat), .ZN(new_n209_));
  INV_X1    g008(.A(G190gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n208_), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND3_X1  g010(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n212_));
  OAI211_X1 g011(.A(new_n211_), .B(new_n212_), .C1(G183gat), .C2(G190gat), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n205_), .B1(new_n202_), .B2(new_n203_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT80), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND4_X1  g015(.A1(new_n206_), .A2(new_n207_), .A3(new_n213_), .A4(new_n216_), .ZN(new_n217_));
  NOR3_X1   g016(.A1(KEYINPUT79), .A2(G169gat), .A3(G176gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(KEYINPUT79), .B1(G169gat), .B2(G176gat), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT24), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n220_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n207_), .B1(new_n222_), .B2(new_n218_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n221_), .B1(new_n223_), .B2(KEYINPUT24), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT25), .B(G183gat), .ZN(new_n225_));
  XNOR2_X1  g024(.A(KEYINPUT26), .B(G190gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n217_), .B1(new_n224_), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G227gat), .A2(G233gat), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n230_), .B(KEYINPUT81), .Z(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT30), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n229_), .B(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(G15gat), .B(G43gat), .Z(new_n234_));
  XNOR2_X1  g033(.A(new_n233_), .B(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G71gat), .B(G99gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n237_), .A2(KEYINPUT83), .ZN(new_n238_));
  OR2_X1    g037(.A1(new_n235_), .A2(new_n236_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT83), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n235_), .A2(new_n236_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n239_), .A2(new_n240_), .A3(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G127gat), .B(G134gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(G113gat), .ZN(new_n244_));
  INV_X1    g043(.A(G120gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G113gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n243_), .B(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(G120gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  XOR2_X1   g049(.A(KEYINPUT82), .B(KEYINPUT31), .Z(new_n251_));
  XNOR2_X1  g050(.A(new_n250_), .B(new_n251_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n238_), .A2(new_n242_), .A3(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n242_), .A2(new_n252_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(KEYINPUT84), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT84), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n253_), .A2(new_n254_), .A3(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n256_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G197gat), .B(G204gat), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(G211gat), .A2(G218gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT21), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G211gat), .A2(G218gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n263_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n265_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT87), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n267_), .A2(new_n262_), .A3(new_n268_), .ZN(new_n269_));
  OAI211_X1 g068(.A(new_n261_), .B(new_n266_), .C1(new_n269_), .C2(new_n264_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n263_), .A2(KEYINPUT87), .A3(new_n265_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n271_), .A2(KEYINPUT21), .A3(new_n260_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT88), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n270_), .A2(KEYINPUT88), .A3(new_n272_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n229_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(G226gat), .A2(G233gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n279_), .B(KEYINPUT19), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  AND3_X1   g080(.A1(new_n227_), .A2(new_n211_), .A3(new_n212_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n223_), .A2(KEYINPUT24), .ZN(new_n283_));
  INV_X1    g082(.A(G169gat), .ZN(new_n284_));
  AOI21_X1  g083(.A(KEYINPUT24), .B1(new_n284_), .B2(new_n205_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n282_), .B1(new_n283_), .B2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n273_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n213_), .A2(new_n207_), .A3(new_n214_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  AND4_X1   g088(.A1(KEYINPUT20), .A2(new_n278_), .A3(new_n281_), .A4(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n282_), .B1(new_n283_), .B2(new_n221_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n275_), .A2(new_n292_), .A3(new_n217_), .A4(new_n276_), .ZN(new_n293_));
  AND3_X1   g092(.A1(new_n293_), .A2(KEYINPUT93), .A3(KEYINPUT20), .ZN(new_n294_));
  AOI21_X1  g093(.A(KEYINPUT93), .B1(new_n293_), .B2(KEYINPUT20), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n286_), .A2(new_n288_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n273_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NOR3_X1   g097(.A1(new_n294_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n291_), .B1(new_n299_), .B2(new_n281_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT18), .B(G64gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(G92gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G8gat), .B(G36gat), .ZN(new_n303_));
  XOR2_X1   g102(.A(new_n302_), .B(new_n303_), .Z(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n300_), .A2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n293_), .A2(KEYINPUT20), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT93), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n307_), .A2(new_n308_), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n293_), .A2(KEYINPUT93), .A3(KEYINPUT20), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(new_n297_), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n290_), .B1(new_n311_), .B2(new_n280_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n304_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n306_), .A2(KEYINPUT94), .A3(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT27), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT94), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n316_), .A3(new_n304_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n314_), .A2(new_n315_), .A3(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319_));
  NOR2_X1   g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n322_), .B(KEYINPUT3), .Z(new_n323_));
  NAND2_X1  g122(.A1(G141gat), .A2(G148gat), .ZN(new_n324_));
  XOR2_X1   g123(.A(new_n324_), .B(KEYINPUT2), .Z(new_n325_));
  OAI21_X1  g124(.A(new_n321_), .B1(new_n323_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n322_), .B1(new_n321_), .B2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n319_), .A2(KEYINPUT1), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n328_), .A2(new_n329_), .A3(new_n324_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n250_), .A2(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n246_), .A2(new_n249_), .A3(new_n330_), .A4(new_n326_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(KEYINPUT4), .A3(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G225gat), .A2(G233gat), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT4), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n250_), .A2(new_n337_), .A3(new_n331_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n334_), .A2(new_n336_), .A3(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n339_), .A2(KEYINPUT95), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n332_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT95), .ZN(new_n342_));
  NAND4_X1  g141(.A1(new_n334_), .A2(new_n342_), .A3(new_n336_), .A4(new_n338_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n340_), .A2(new_n341_), .A3(new_n343_), .ZN(new_n344_));
  XOR2_X1   g143(.A(G1gat), .B(G29gat), .Z(new_n345_));
  XNOR2_X1  g144(.A(G57gat), .B(G85gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT96), .B(KEYINPUT0), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n344_), .A2(new_n349_), .ZN(new_n350_));
  INV_X1    g149(.A(new_n349_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n340_), .A2(new_n341_), .A3(new_n351_), .A4(new_n343_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n331_), .A2(KEYINPUT29), .ZN(new_n354_));
  XNOR2_X1  g153(.A(KEYINPUT85), .B(KEYINPUT28), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n354_), .A2(new_n355_), .ZN(new_n357_));
  XNOR2_X1  g156(.A(G22gat), .B(G50gat), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  OR3_X1    g158(.A1(new_n356_), .A2(new_n357_), .A3(new_n359_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n359_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n331_), .A2(KEYINPUT29), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G228gat), .A2(G233gat), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n363_), .B(KEYINPUT86), .Z(new_n364_));
  NAND3_X1  g163(.A1(new_n277_), .A2(new_n362_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n287_), .A2(KEYINPUT89), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT89), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n273_), .A2(new_n367_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n366_), .A2(new_n368_), .B1(KEYINPUT29), .B2(new_n331_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n365_), .B1(new_n369_), .B2(new_n363_), .ZN(new_n370_));
  XNOR2_X1  g169(.A(G78gat), .B(G106gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(KEYINPUT90), .ZN(new_n372_));
  AOI21_X1  g171(.A(KEYINPUT91), .B1(new_n370_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n372_), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n365_), .B(new_n374_), .C1(new_n369_), .C2(new_n363_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  NOR3_X1   g176(.A1(new_n370_), .A2(KEYINPUT91), .A3(new_n372_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n360_), .B(new_n361_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n360_), .A2(new_n361_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n370_), .A2(new_n371_), .ZN(new_n381_));
  INV_X1    g180(.A(KEYINPUT92), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n375_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n376_), .A2(KEYINPUT92), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n380_), .A2(new_n381_), .A3(new_n383_), .A4(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n353_), .B1(new_n379_), .B2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n366_), .A2(new_n368_), .ZN(new_n387_));
  OAI211_X1 g186(.A(new_n278_), .B(KEYINPUT20), .C1(new_n296_), .C2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n280_), .ZN(new_n389_));
  OAI21_X1  g188(.A(new_n389_), .B1(new_n311_), .B2(new_n280_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(new_n305_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n391_), .A2(new_n313_), .A3(KEYINPUT27), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n318_), .A2(new_n386_), .A3(new_n392_), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT100), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  NAND4_X1  g194(.A1(new_n318_), .A2(new_n386_), .A3(new_n392_), .A4(KEYINPUT100), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n379_), .A2(new_n385_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n314_), .A2(new_n317_), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n334_), .A2(new_n335_), .A3(new_n338_), .ZN(new_n400_));
  XOR2_X1   g199(.A(new_n400_), .B(KEYINPUT98), .Z(new_n401_));
  NAND3_X1  g200(.A1(new_n332_), .A2(new_n333_), .A3(new_n336_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(new_n349_), .ZN(new_n403_));
  XOR2_X1   g202(.A(new_n403_), .B(KEYINPUT97), .Z(new_n404_));
  NAND2_X1  g203(.A1(new_n401_), .A2(new_n404_), .ZN(new_n405_));
  OR2_X1    g204(.A1(new_n405_), .A2(KEYINPUT99), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n352_), .B(KEYINPUT33), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(KEYINPUT99), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n399_), .A2(new_n406_), .A3(new_n407_), .A4(new_n408_), .ZN(new_n409_));
  AND2_X1   g208(.A1(new_n304_), .A2(KEYINPUT32), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n390_), .A2(new_n410_), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n353_), .B(new_n411_), .C1(new_n300_), .C2(new_n410_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n398_), .B1(new_n409_), .B2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n259_), .B1(new_n397_), .B2(new_n413_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT101), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  AND2_X1   g215(.A1(new_n318_), .A2(new_n392_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n418_), .A2(new_n255_), .A3(new_n398_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n353_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  OAI211_X1 g220(.A(new_n259_), .B(KEYINPUT101), .C1(new_n397_), .C2(new_n413_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n416_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  AND2_X1   g222(.A1(G57gat), .A2(G64gat), .ZN(new_n424_));
  NOR2_X1   g223(.A1(G57gat), .A2(G64gat), .ZN(new_n425_));
  NOR2_X1   g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT11), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT65), .ZN(new_n430_));
  NOR2_X1   g229(.A1(G71gat), .A2(G78gat), .ZN(new_n431_));
  AOI21_X1  g230(.A(new_n431_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G71gat), .A2(G78gat), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n430_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(G57gat), .ZN(new_n435_));
  INV_X1    g234(.A(G64gat), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G57gat), .A2(G64gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n427_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n431_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n433_), .A3(new_n440_), .ZN(new_n441_));
  NOR2_X1   g240(.A1(new_n441_), .A2(KEYINPUT65), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n429_), .B1(new_n434_), .B2(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n432_), .A2(new_n430_), .A3(new_n433_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(KEYINPUT65), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n444_), .A2(new_n428_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT64), .ZN(new_n448_));
  OAI21_X1  g247(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NOR3_X1   g249(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n448_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G99gat), .A2(G106gat), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND3_X1  g254(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n456_));
  AND2_X1   g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT7), .ZN(new_n458_));
  INV_X1    g257(.A(G99gat), .ZN(new_n459_));
  INV_X1    g258(.A(G106gat), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n459_), .A3(new_n460_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(KEYINPUT64), .A3(new_n449_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n452_), .A2(new_n457_), .A3(new_n462_), .ZN(new_n463_));
  XOR2_X1   g262(.A(G85gat), .B(G92gat), .Z(new_n464_));
  NAND3_X1  g263(.A1(new_n463_), .A2(KEYINPUT8), .A3(new_n464_), .ZN(new_n465_));
  XOR2_X1   g264(.A(KEYINPUT10), .B(G99gat), .Z(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(new_n460_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n464_), .A2(KEYINPUT9), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT9), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(G85gat), .A3(G92gat), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n467_), .A2(new_n468_), .A3(new_n470_), .A4(new_n457_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n461_), .A2(new_n455_), .A3(new_n456_), .A4(new_n449_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(new_n464_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT8), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(new_n465_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n447_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n465_), .A2(new_n471_), .A3(new_n475_), .ZN(new_n478_));
  NAND4_X1  g277(.A1(new_n478_), .A2(KEYINPUT12), .A3(new_n446_), .A4(new_n443_), .ZN(new_n479_));
  AND2_X1   g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G230gat), .A2(G233gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n446_), .A3(new_n443_), .ZN(new_n482_));
  XOR2_X1   g281(.A(KEYINPUT66), .B(KEYINPUT12), .Z(new_n483_));
  NAND2_X1  g282(.A1(new_n482_), .A2(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n480_), .A2(new_n481_), .A3(new_n484_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n477_), .A2(new_n482_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n485_), .B1(new_n481_), .B2(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G120gat), .B(G148gat), .ZN(new_n488_));
  INV_X1    g287(.A(G204gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n488_), .B(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n490_), .B(KEYINPUT5), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(new_n205_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n487_), .B(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT67), .B(KEYINPUT13), .Z(new_n495_));
  OR2_X1    g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n494_), .B1(KEYINPUT67), .B2(KEYINPUT13), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(new_n498_), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G113gat), .B(G141gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(new_n284_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(G197gat), .ZN(new_n502_));
  XOR2_X1   g301(.A(new_n502_), .B(KEYINPUT78), .Z(new_n503_));
  XNOR2_X1  g302(.A(G15gat), .B(G22gat), .ZN(new_n504_));
  INV_X1    g303(.A(G1gat), .ZN(new_n505_));
  INV_X1    g304(.A(G8gat), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT14), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n504_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G1gat), .B(G8gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  XOR2_X1   g309(.A(G29gat), .B(G36gat), .Z(new_n511_));
  INV_X1    g310(.A(G43gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G29gat), .B(G36gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n514_), .A2(G43gat), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n513_), .A2(G50gat), .A3(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(G50gat), .B1(new_n513_), .B2(new_n515_), .ZN(new_n517_));
  OAI21_X1  g316(.A(KEYINPUT69), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(G50gat), .ZN(new_n519_));
  INV_X1    g318(.A(new_n515_), .ZN(new_n520_));
  NOR2_X1   g319(.A1(new_n514_), .A2(G43gat), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n519_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT69), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n513_), .A2(G50gat), .A3(new_n515_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n518_), .A2(KEYINPUT15), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(KEYINPUT15), .B1(new_n518_), .B2(new_n525_), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n510_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(G229gat), .A2(G233gat), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n522_), .A2(new_n524_), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(new_n510_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n529_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n531_), .A2(new_n510_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT76), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n530_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n533_), .A2(KEYINPUT76), .A3(new_n535_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n538_), .A2(new_n539_), .A3(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n534_), .A2(new_n541_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n503_), .B1(new_n542_), .B2(KEYINPUT77), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT77), .ZN(new_n544_));
  INV_X1    g343(.A(new_n503_), .ZN(new_n545_));
  AOI211_X1 g344(.A(new_n544_), .B(new_n545_), .C1(new_n534_), .C2(new_n541_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n543_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n499_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G190gat), .B(G218gat), .ZN(new_n550_));
  XNOR2_X1  g349(.A(new_n550_), .B(G134gat), .ZN(new_n551_));
  XOR2_X1   g350(.A(new_n551_), .B(G162gat), .Z(new_n552_));
  INV_X1    g351(.A(KEYINPUT36), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n478_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n531_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n476_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT34), .ZN(new_n559_));
  OR2_X1    g358(.A1(new_n559_), .A2(KEYINPUT35), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT70), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n559_), .A2(KEYINPUT35), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT68), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n555_), .A2(new_n562_), .A3(new_n563_), .A4(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n563_), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n565_), .A2(new_n563_), .ZN(new_n568_));
  INV_X1    g367(.A(KEYINPUT15), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n516_), .A2(new_n517_), .A3(KEYINPUT69), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n523_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n569_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  AOI21_X1  g371(.A(new_n476_), .B1(new_n572_), .B2(new_n526_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n567_), .B(new_n568_), .C1(new_n573_), .C2(new_n561_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n554_), .B1(new_n566_), .B2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(KEYINPUT37), .B1(new_n575_), .B2(KEYINPUT71), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n576_), .A2(KEYINPUT72), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT72), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n578_), .B(KEYINPUT37), .C1(new_n575_), .C2(KEYINPUT71), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n575_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n566_), .A2(new_n574_), .A3(new_n554_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n552_), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n581_), .A2(new_n582_), .B1(KEYINPUT36), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n580_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G183gat), .B(G211gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(G155gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XOR2_X1   g389(.A(KEYINPUT74), .B(G127gat), .Z(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n592_), .B(KEYINPUT17), .ZN(new_n593_));
  NAND2_X1  g392(.A1(G231gat), .A2(G233gat), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n510_), .B(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(new_n595_), .B(new_n447_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT17), .ZN(new_n598_));
  OR3_X1    g397(.A1(new_n596_), .A2(new_n598_), .A3(new_n592_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT75), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n577_), .A2(new_n584_), .A3(new_n579_), .ZN(new_n602_));
  AND3_X1   g401(.A1(new_n586_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  AND3_X1   g402(.A1(new_n423_), .A2(new_n549_), .A3(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n353_), .B(KEYINPUT102), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n505_), .A3(new_n606_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT38), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n423_), .A2(new_n584_), .A3(new_n549_), .A4(new_n600_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n609_), .B2(new_n420_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(G1324gat));
  NAND3_X1  g410(.A1(new_n604_), .A2(new_n506_), .A3(new_n418_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT103), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(G8gat), .B1(new_n609_), .B2(new_n417_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT39), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  OR2_X1    g416(.A1(new_n615_), .A2(new_n616_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n614_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT40), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n614_), .A2(new_n617_), .A3(KEYINPUT40), .A4(new_n618_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(G1325gat));
  INV_X1    g422(.A(G15gat), .ZN(new_n624_));
  INV_X1    g423(.A(new_n259_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n604_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G15gat), .B1(new_n609_), .B2(new_n259_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n627_), .A2(KEYINPUT104), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(KEYINPUT104), .ZN(new_n629_));
  AND3_X1   g428(.A1(new_n628_), .A2(KEYINPUT41), .A3(new_n629_), .ZN(new_n630_));
  AOI21_X1  g429(.A(KEYINPUT41), .B1(new_n628_), .B2(new_n629_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n626_), .B1(new_n630_), .B2(new_n631_), .ZN(G1326gat));
  XOR2_X1   g431(.A(new_n398_), .B(KEYINPUT105), .Z(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  OAI21_X1  g433(.A(G22gat), .B1(new_n609_), .B2(new_n634_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n635_), .B(KEYINPUT42), .ZN(new_n636_));
  INV_X1    g435(.A(G22gat), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n604_), .A2(new_n637_), .A3(new_n633_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n636_), .A2(new_n638_), .ZN(G1327gat));
  INV_X1    g438(.A(new_n601_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n549_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n423_), .A2(new_n585_), .A3(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(G29gat), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n353_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n586_), .A2(new_n602_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n423_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n647_), .A2(KEYINPUT43), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n423_), .A2(new_n649_), .A3(new_n646_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n641_), .B1(new_n648_), .B2(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n651_), .A2(KEYINPUT44), .ZN(new_n652_));
  AND3_X1   g451(.A1(new_n423_), .A2(new_n649_), .A3(new_n646_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n649_), .B1(new_n423_), .B2(new_n646_), .ZN(new_n654_));
  OAI211_X1 g453(.A(KEYINPUT44), .B(new_n642_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n606_), .ZN(new_n656_));
  OAI211_X1 g455(.A(KEYINPUT106), .B(G29gat), .C1(new_n652_), .C2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n642_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT44), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n661_), .A2(new_n606_), .A3(new_n655_), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT106), .B1(new_n662_), .B2(G29gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n645_), .B1(new_n658_), .B2(new_n663_), .ZN(G1328gat));
  INV_X1    g463(.A(KEYINPUT46), .ZN(new_n665_));
  INV_X1    g464(.A(G36gat), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n417_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n667_), .B2(new_n655_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n643_), .A2(new_n666_), .A3(new_n418_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT45), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n669_), .B(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n665_), .B1(new_n668_), .B2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n418_), .B1(new_n651_), .B2(KEYINPUT44), .ZN(new_n673_));
  INV_X1    g472(.A(new_n655_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G36gat), .B1(new_n673_), .B2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n669_), .B(KEYINPUT45), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n675_), .A2(KEYINPUT46), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n672_), .A2(new_n677_), .ZN(G1329gat));
  NAND2_X1  g477(.A1(new_n643_), .A2(new_n625_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n679_), .A2(new_n512_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n254_), .B(new_n253_), .C1(new_n651_), .C2(KEYINPUT44), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n655_), .A2(G43gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n680_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT47), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT47), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n685_), .B(new_n680_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(G1330gat));
  NAND2_X1  g486(.A1(new_n633_), .A2(new_n519_), .ZN(new_n688_));
  XOR2_X1   g487(.A(new_n688_), .B(KEYINPUT107), .Z(new_n689_));
  NAND2_X1  g488(.A1(new_n643_), .A2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n398_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n652_), .A2(new_n674_), .A3(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(new_n690_), .B1(new_n692_), .B2(new_n519_), .ZN(G1331gat));
  NAND2_X1  g492(.A1(new_n499_), .A2(new_n548_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n694_), .A2(new_n640_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n423_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n584_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n697_), .A2(new_n435_), .A3(new_n420_), .ZN(new_n698_));
  AND3_X1   g497(.A1(new_n696_), .A2(new_n602_), .A3(new_n586_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(new_n606_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n698_), .B1(new_n700_), .B2(new_n435_), .ZN(G1332gat));
  INV_X1    g500(.A(new_n697_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n702_), .A2(new_n418_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n703_), .A2(G64gat), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT108), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n703_), .A2(new_n706_), .A3(G64gat), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n705_), .A2(KEYINPUT48), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n706_), .B1(new_n703_), .B2(G64gat), .ZN(new_n710_));
  AOI211_X1 g509(.A(KEYINPUT108), .B(new_n436_), .C1(new_n702_), .C2(new_n418_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n709_), .B1(new_n710_), .B2(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n699_), .A2(new_n436_), .A3(new_n418_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n708_), .A2(new_n712_), .A3(new_n713_), .ZN(G1333gat));
  OAI21_X1  g513(.A(G71gat), .B1(new_n697_), .B2(new_n259_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT49), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n259_), .A2(G71gat), .ZN(new_n717_));
  XNOR2_X1  g516(.A(new_n717_), .B(KEYINPUT109), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n699_), .A2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n716_), .A2(new_n719_), .ZN(G1334gat));
  INV_X1    g519(.A(G78gat), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n699_), .A2(new_n721_), .A3(new_n633_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n696_), .A2(new_n584_), .A3(new_n633_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT50), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(G78gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G78gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT110), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n727_), .B(new_n728_), .ZN(G1335gat));
  AND2_X1   g528(.A1(new_n423_), .A2(new_n585_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n694_), .A2(new_n601_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n732_), .ZN(new_n733_));
  AOI21_X1  g532(.A(G85gat), .B1(new_n733_), .B2(new_n606_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT111), .ZN(new_n735_));
  AOI211_X1 g534(.A(new_n601_), .B(new_n694_), .C1(new_n648_), .C2(new_n650_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n736_), .A2(G85gat), .A3(new_n353_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n735_), .A2(new_n737_), .ZN(G1336gat));
  NAND3_X1  g537(.A1(new_n736_), .A2(G92gat), .A3(new_n418_), .ZN(new_n739_));
  INV_X1    g538(.A(G92gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n740_), .B1(new_n732_), .B2(new_n417_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n739_), .A2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT112), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n739_), .A2(new_n744_), .A3(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1337gat));
  AOI21_X1  g545(.A(new_n459_), .B1(new_n736_), .B2(new_n625_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(KEYINPUT51), .ZN(new_n749_));
  INV_X1    g548(.A(new_n466_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n732_), .A2(new_n750_), .A3(new_n255_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n748_), .A2(new_n749_), .A3(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(KEYINPUT51), .B1(new_n747_), .B2(new_n751_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n753_), .A2(new_n754_), .ZN(G1338gat));
  NAND3_X1  g554(.A1(new_n733_), .A2(new_n460_), .A3(new_n398_), .ZN(new_n756_));
  OAI211_X1 g555(.A(new_n398_), .B(new_n731_), .C1(new_n653_), .C2(new_n654_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758_));
  AND3_X1   g557(.A1(new_n757_), .A2(new_n758_), .A3(G106gat), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n758_), .B1(new_n757_), .B2(G106gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n756_), .B1(new_n759_), .B2(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n761_), .A2(KEYINPUT53), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT53), .ZN(new_n763_));
  OAI211_X1 g562(.A(new_n763_), .B(new_n756_), .C1(new_n759_), .C2(new_n760_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n762_), .A2(new_n764_), .ZN(G1339gat));
  INV_X1    g564(.A(KEYINPUT113), .ZN(new_n766_));
  NAND4_X1  g565(.A1(new_n603_), .A2(new_n766_), .A3(new_n498_), .A4(new_n548_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n586_), .A2(new_n548_), .A3(new_n601_), .A4(new_n602_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT113), .B1(new_n768_), .B2(new_n499_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT54), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n767_), .A2(new_n769_), .A3(KEYINPUT54), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT115), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT55), .ZN(new_n776_));
  INV_X1    g575(.A(new_n481_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n776_), .B1(new_n777_), .B2(KEYINPUT114), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n484_), .A2(new_n477_), .A3(new_n479_), .A4(new_n779_), .ZN(new_n780_));
  NOR2_X1   g579(.A1(new_n481_), .A2(KEYINPUT55), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n779_), .B1(new_n480_), .B2(new_n484_), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n775_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n484_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n477_), .A2(new_n479_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n778_), .B1(new_n785_), .B2(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n787_), .B(KEYINPUT115), .C1(new_n781_), .C2(new_n780_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n784_), .A2(new_n493_), .A3(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n789_), .A2(KEYINPUT56), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT56), .ZN(new_n791_));
  NAND4_X1  g590(.A1(new_n784_), .A2(new_n791_), .A3(new_n788_), .A4(new_n493_), .ZN(new_n792_));
  AND2_X1   g591(.A1(new_n790_), .A2(new_n792_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n487_), .A2(new_n493_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n793_), .A2(KEYINPUT116), .A3(new_n794_), .A4(new_n547_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n529_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n539_), .B1(new_n796_), .B2(new_n532_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n538_), .A2(new_n540_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n530_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n502_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n534_), .A2(new_n541_), .A3(new_n502_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n494_), .A2(new_n802_), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n790_), .A2(new_n547_), .A3(new_n794_), .A4(new_n792_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT116), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n795_), .A2(new_n803_), .A3(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(KEYINPUT57), .A3(new_n584_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT119), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n807_), .A2(KEYINPUT119), .A3(KEYINPUT57), .A4(new_n584_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT57), .B1(new_n807_), .B2(new_n584_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n790_), .A2(new_n794_), .A3(new_n802_), .A4(new_n792_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(KEYINPUT58), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n814_), .A2(new_n815_), .A3(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n646_), .A3(new_n819_), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n813_), .B1(KEYINPUT118), .B2(new_n820_), .ZN(new_n821_));
  OR2_X1    g620(.A1(new_n820_), .A2(KEYINPUT118), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n812_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(new_n600_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n774_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n419_), .A2(new_n606_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n547_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT59), .B1(new_n825_), .B2(new_n826_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT59), .ZN(new_n830_));
  XOR2_X1   g629(.A(new_n826_), .B(KEYINPUT120), .Z(new_n831_));
  XNOR2_X1  g630(.A(new_n804_), .B(KEYINPUT116), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n585_), .B1(new_n832_), .B2(new_n803_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n820_), .B1(new_n833_), .B2(KEYINPUT57), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT121), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n834_), .A2(new_n835_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n836_));
  OAI211_X1 g635(.A(KEYINPUT121), .B(new_n820_), .C1(new_n833_), .C2(KEYINPUT57), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n601_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  OAI211_X1 g637(.A(new_n830_), .B(new_n831_), .C1(new_n838_), .C2(new_n774_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT122), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n829_), .A2(new_n839_), .A3(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n840_), .B1(new_n829_), .B2(new_n839_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n548_), .A2(new_n247_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n828_), .B1(new_n843_), .B2(new_n844_), .ZN(G1340gat));
  XNOR2_X1  g644(.A(KEYINPUT123), .B(G120gat), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n498_), .A2(new_n846_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n827_), .B1(KEYINPUT60), .B2(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n849_), .B2(KEYINPUT60), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n849_), .A2(new_n499_), .A3(new_n829_), .A4(new_n839_), .ZN(new_n851_));
  AND2_X1   g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1341gat));
  AOI21_X1  g651(.A(G127gat), .B1(new_n827_), .B2(new_n601_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n600_), .A2(G127gat), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n853_), .B1(new_n843_), .B2(new_n854_), .ZN(G1342gat));
  AOI21_X1  g654(.A(G134gat), .B1(new_n827_), .B2(new_n585_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n646_), .A2(G134gat), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n856_), .B1(new_n843_), .B2(new_n857_), .ZN(G1343gat));
  NOR3_X1   g657(.A1(new_n825_), .A2(new_n691_), .A3(new_n625_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n418_), .A2(new_n605_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n547_), .A3(new_n860_), .ZN(new_n861_));
  XNOR2_X1  g660(.A(new_n861_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g661(.A1(new_n859_), .A2(new_n499_), .A3(new_n860_), .ZN(new_n863_));
  XNOR2_X1  g662(.A(new_n863_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g663(.A1(new_n859_), .A2(new_n601_), .A3(new_n860_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT61), .B(G155gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1346gat));
  AND3_X1   g666(.A1(new_n859_), .A2(new_n585_), .A3(new_n860_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n859_), .A2(new_n646_), .A3(new_n860_), .ZN(new_n869_));
  MUX2_X1   g668(.A(new_n868_), .B(new_n869_), .S(G162gat), .Z(G1347gat));
  INV_X1    g669(.A(KEYINPUT62), .ZN(new_n871_));
  INV_X1    g670(.A(new_n820_), .ZN(new_n872_));
  OAI21_X1  g671(.A(new_n835_), .B1(new_n813_), .B2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n812_), .A2(new_n837_), .A3(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n774_), .B1(new_n874_), .B2(new_n640_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n259_), .A2(new_n606_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n876_), .A2(new_n418_), .A3(new_n634_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n875_), .A2(new_n548_), .A3(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n871_), .B1(new_n878_), .B2(new_n284_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n878_), .A2(new_n204_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n877_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n881_), .B(new_n547_), .C1(new_n838_), .C2(new_n774_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n882_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n883_));
  NAND3_X1  g682(.A1(new_n879_), .A2(new_n880_), .A3(new_n883_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT124), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  NAND4_X1  g685(.A1(new_n879_), .A2(KEYINPUT124), .A3(new_n883_), .A4(new_n880_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n886_), .A2(new_n887_), .ZN(G1348gat));
  NOR2_X1   g687(.A1(new_n875_), .A2(new_n877_), .ZN(new_n889_));
  AOI21_X1  g688(.A(G176gat), .B1(new_n889_), .B2(new_n499_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n823_), .A2(new_n824_), .ZN(new_n891_));
  INV_X1    g690(.A(new_n774_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n893_), .A2(new_n691_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n876_), .A2(new_n418_), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n894_), .A2(new_n205_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n890_), .B1(new_n896_), .B2(new_n499_), .ZN(G1349gat));
  OR3_X1    g696(.A1(new_n894_), .A2(new_n640_), .A3(new_n895_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n824_), .A2(new_n225_), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n898_), .A2(new_n209_), .B1(new_n889_), .B2(new_n899_), .ZN(G1350gat));
  NAND3_X1  g699(.A1(new_n889_), .A2(new_n585_), .A3(new_n226_), .ZN(new_n901_));
  AND2_X1   g700(.A1(new_n889_), .A2(new_n646_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n902_), .B2(new_n210_), .ZN(G1351gat));
  NOR3_X1   g702(.A1(new_n417_), .A2(new_n353_), .A3(new_n691_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n893_), .A2(new_n259_), .A3(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n547_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n499_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n489_), .A2(KEYINPUT125), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1353gat));
  AOI211_X1 g710(.A(KEYINPUT63), .B(G211gat), .C1(new_n906_), .C2(new_n600_), .ZN(new_n912_));
  XOR2_X1   g711(.A(KEYINPUT63), .B(G211gat), .Z(new_n913_));
  AND3_X1   g712(.A1(new_n906_), .A2(new_n600_), .A3(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n912_), .A2(new_n914_), .ZN(G1354gat));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(new_n905_), .B2(new_n584_), .ZN(new_n917_));
  INV_X1    g716(.A(G218gat), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n825_), .A2(new_n625_), .ZN(new_n919_));
  NAND4_X1  g718(.A1(new_n919_), .A2(KEYINPUT126), .A3(new_n585_), .A4(new_n904_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n917_), .A2(new_n918_), .A3(new_n920_), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n906_), .A2(G218gat), .A3(new_n646_), .ZN(new_n922_));
  AND2_X1   g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1355gat));
endmodule


