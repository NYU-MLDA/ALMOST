//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n863_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n870_,
    new_n871_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n960_, new_n961_, new_n962_, new_n963_, new_n965_,
    new_n966_, new_n968_, new_n970_, new_n971_, new_n972_, new_n973_,
    new_n974_, new_n975_, new_n976_, new_n977_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n999_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1008_,
    new_n1009_, new_n1010_, new_n1011_, new_n1013_, new_n1014_, new_n1015_,
    new_n1017_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1029_, new_n1030_,
    new_n1031_;
  INV_X1    g000(.A(KEYINPUT7), .ZN(new_n202_));
  INV_X1    g001(.A(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G85gat), .A2(G92gat), .ZN(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G85gat), .A2(G92gat), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n213_), .A2(new_n214_), .A3(KEYINPUT8), .ZN(new_n215_));
  AOI21_X1  g014(.A(KEYINPUT66), .B1(new_n211_), .B2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n211_), .A2(KEYINPUT66), .A3(new_n215_), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n213_), .A2(new_n214_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n207_), .A2(KEYINPUT67), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n222_), .A2(KEYINPUT6), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n206_), .B1(new_n221_), .B2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n205_), .A2(new_n210_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  AND3_X1   g025(.A1(new_n221_), .A2(new_n223_), .A3(new_n206_), .ZN(new_n227_));
  INV_X1    g026(.A(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n220_), .B1(new_n226_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT8), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n217_), .B(new_n218_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n231_));
  AND2_X1   g030(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n232_));
  NOR2_X1   g031(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT64), .ZN(new_n234_));
  NOR3_X1   g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT64), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n204_), .B1(new_n235_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT9), .ZN(new_n240_));
  NOR3_X1   g039(.A1(new_n213_), .A2(new_n214_), .A3(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n240_), .A2(G85gat), .A3(G92gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n208_), .A2(new_n242_), .A3(new_n209_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n239_), .A2(KEYINPUT65), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n236_), .A2(KEYINPUT64), .A3(new_n237_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n234_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n248_));
  AOI21_X1  g047(.A(G106gat), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  AND3_X1   g048(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(G85gat), .ZN(new_n253_));
  INV_X1    g052(.A(G92gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n255_), .A2(KEYINPUT9), .A3(new_n212_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n252_), .A2(new_n256_), .A3(new_n242_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n246_), .B1(new_n249_), .B2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n245_), .A2(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G71gat), .B(G78gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G57gat), .B(G64gat), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT11), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n260_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n261_), .A2(KEYINPUT11), .ZN(new_n265_));
  XNOR2_X1  g064(.A(new_n264_), .B(new_n265_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n231_), .A2(new_n259_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G230gat), .A2(G233gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  NOR3_X1   g068(.A1(new_n227_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n270_));
  OAI21_X1  g069(.A(KEYINPUT8), .B1(new_n270_), .B2(new_n220_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n211_), .A2(KEYINPUT66), .A3(new_n215_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n272_), .A2(new_n216_), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n271_), .A2(new_n273_), .B1(new_n258_), .B2(new_n245_), .ZN(new_n274_));
  OAI21_X1  g073(.A(KEYINPUT12), .B1(new_n274_), .B2(new_n266_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n231_), .A2(new_n259_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT12), .ZN(new_n277_));
  INV_X1    g076(.A(new_n266_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n276_), .A2(new_n277_), .A3(new_n278_), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n269_), .B1(new_n275_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n268_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n274_), .A2(new_n266_), .ZN(new_n283_));
  AND3_X1   g082(.A1(new_n231_), .A2(new_n259_), .A3(new_n266_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n282_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  AND2_X1   g084(.A1(new_n285_), .A2(KEYINPUT68), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT68), .ZN(new_n287_));
  OAI211_X1 g086(.A(new_n287_), .B(new_n282_), .C1(new_n283_), .C2(new_n284_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n281_), .B1(new_n286_), .B2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(G120gat), .B(G148gat), .ZN(new_n291_));
  INV_X1    g090(.A(G204gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G176gat), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n293_), .B(new_n294_), .Z(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n290_), .A2(KEYINPUT69), .A3(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n285_), .A2(KEYINPUT68), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n280_), .B1(new_n299_), .B2(new_n288_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n298_), .B1(new_n300_), .B2(new_n295_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  OAI211_X1 g101(.A(new_n281_), .B(new_n295_), .C1(new_n286_), .C2(new_n289_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n300_), .A2(KEYINPUT70), .A3(new_n295_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n302_), .A2(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT13), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT81), .ZN(new_n311_));
  XOR2_X1   g110(.A(G1gat), .B(G8gat), .Z(new_n312_));
  INV_X1    g111(.A(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(G1gat), .A2(G8gat), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT14), .ZN(new_n315_));
  INV_X1    g114(.A(G15gat), .ZN(new_n316_));
  INV_X1    g115(.A(G22gat), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G15gat), .A2(G22gat), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n315_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n320_), .A2(KEYINPUT75), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n320_), .A2(KEYINPUT75), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n313_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n323_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(new_n312_), .A3(new_n321_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(G29gat), .B(G36gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G43gat), .B(G50gat), .Z(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G43gat), .B(G50gat), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n328_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n331_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n327_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT80), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n311_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n334_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n338_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n339_), .A2(KEYINPUT80), .A3(KEYINPUT81), .ZN(new_n340_));
  OAI22_X1  g139(.A1(new_n337_), .A2(new_n340_), .B1(new_n334_), .B2(new_n327_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n335_), .A2(new_n336_), .A3(new_n311_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n327_), .A2(new_n334_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT81), .B1(new_n339_), .B2(KEYINPUT80), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n342_), .A2(new_n343_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G229gat), .A2(G233gat), .ZN(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n341_), .A2(new_n345_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT15), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n334_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n331_), .A2(KEYINPUT15), .A3(new_n333_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n327_), .A2(new_n352_), .ZN(new_n353_));
  NOR3_X1   g152(.A1(new_n353_), .A2(new_n347_), .A3(new_n339_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n348_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G113gat), .B(G141gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G169gat), .ZN(new_n358_));
  INV_X1    g157(.A(G197gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(new_n358_), .B(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n356_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n348_), .A2(new_n355_), .A3(new_n360_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT78), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G231gat), .A2(G233gat), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n366_), .B(KEYINPUT76), .Z(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n324_), .A2(new_n326_), .A3(new_n368_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n278_), .A3(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n266_), .B1(new_n373_), .B2(new_n369_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT17), .ZN(new_n376_));
  XNOR2_X1  g175(.A(G183gat), .B(G211gat), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G127gat), .B(G155gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  XNOR2_X1  g178(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n379_), .B(new_n380_), .ZN(new_n381_));
  OR3_X1    g180(.A1(new_n375_), .A2(new_n376_), .A3(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n381_), .B(KEYINPUT17), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n375_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT79), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n384_), .A2(KEYINPUT79), .ZN(new_n386_));
  AND4_X1   g185(.A1(new_n365_), .A2(new_n382_), .A3(new_n385_), .A4(new_n386_), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n386_), .A2(new_n385_), .B1(new_n382_), .B2(new_n365_), .ZN(new_n388_));
  OR2_X1    g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n302_), .A2(new_n307_), .A3(KEYINPUT13), .ZN(new_n390_));
  NAND4_X1  g189(.A1(new_n310_), .A2(new_n364_), .A3(new_n389_), .A4(new_n390_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n391_), .A2(KEYINPUT100), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n391_), .A2(KEYINPUT100), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(G57gat), .B(G85gat), .Z(new_n395_));
  XNOR2_X1  g194(.A(G1gat), .B(G29gat), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n395_), .B(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G127gat), .B(G134gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(G113gat), .B(G120gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(new_n400_), .B(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G155gat), .B(G162gat), .ZN(new_n404_));
  INV_X1    g203(.A(G141gat), .ZN(new_n405_));
  INV_X1    g204(.A(G148gat), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  OAI21_X1  g206(.A(KEYINPUT89), .B1(new_n407_), .B2(KEYINPUT3), .ZN(new_n408_));
  NOR2_X1   g207(.A1(G141gat), .A2(G148gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT89), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n409_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G141gat), .A2(G148gat), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT2), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n417_));
  OAI21_X1  g216(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n416_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n404_), .B1(new_n413_), .B2(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n407_), .A2(new_n414_), .A3(new_n421_), .ZN(new_n422_));
  XOR2_X1   g221(.A(G155gat), .B(G162gat), .Z(new_n423_));
  INV_X1    g222(.A(KEYINPUT1), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n403_), .B1(new_n420_), .B2(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n418_), .A2(new_n417_), .ZN(new_n427_));
  NOR4_X1   g226(.A1(KEYINPUT89), .A2(KEYINPUT3), .A3(G141gat), .A4(G148gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n410_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n427_), .B(new_n416_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n425_), .B1(new_n423_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n402_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n426_), .A2(new_n432_), .A3(KEYINPUT4), .ZN(new_n433_));
  OR3_X1    g232(.A1(new_n431_), .A2(KEYINPUT4), .A3(new_n402_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(G225gat), .A2(G233gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(new_n437_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n437_), .B1(new_n426_), .B2(new_n432_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n399_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n436_), .B1(new_n433_), .B2(new_n434_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n399_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n442_), .A2(new_n443_), .A3(new_n439_), .ZN(new_n444_));
  NOR2_X1   g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT86), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G227gat), .A2(G233gat), .ZN(new_n448_));
  XOR2_X1   g247(.A(new_n448_), .B(KEYINPUT85), .Z(new_n449_));
  XNOR2_X1  g248(.A(G71gat), .B(G99gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(KEYINPUT82), .A2(G190gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(KEYINPUT26), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT26), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(KEYINPUT82), .A3(G190gat), .ZN(new_n455_));
  INV_X1    g254(.A(G183gat), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n456_), .A2(KEYINPUT25), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT25), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n458_), .A2(G183gat), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n453_), .A2(new_n455_), .A3(new_n457_), .A4(new_n459_), .ZN(new_n460_));
  NOR2_X1   g259(.A1(G169gat), .A2(G176gat), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(G169gat), .A2(G176gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(KEYINPUT24), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT24), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  AND3_X1   g265(.A1(new_n460_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(G183gat), .A2(G190gat), .ZN(new_n468_));
  AND2_X1   g267(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n469_));
  NOR2_X1   g268(.A1(KEYINPUT83), .A2(KEYINPUT23), .ZN(new_n470_));
  OAI21_X1  g269(.A(new_n468_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT84), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT84), .ZN(new_n473_));
  OAI211_X1 g272(.A(new_n473_), .B(new_n468_), .C1(new_n469_), .C2(new_n470_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n468_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT23), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n472_), .A2(new_n474_), .A3(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n467_), .A2(new_n478_), .ZN(new_n479_));
  XNOR2_X1  g278(.A(KEYINPUT22), .B(G169gat), .ZN(new_n480_));
  INV_X1    g279(.A(G176gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n468_), .A2(KEYINPUT23), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n469_), .A2(new_n470_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(new_n485_), .B2(new_n475_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(G183gat), .A2(G190gat), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n463_), .B(new_n482_), .C1(new_n486_), .C2(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n479_), .A2(new_n488_), .A3(KEYINPUT30), .ZN(new_n489_));
  AOI21_X1  g288(.A(KEYINPUT30), .B1(new_n479_), .B2(new_n488_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n451_), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G15gat), .B(G43gat), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT30), .ZN(new_n493_));
  NAND3_X1  g292(.A1(new_n460_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n494_));
  AOI22_X1  g293(.A1(new_n471_), .A2(KEYINPUT84), .B1(new_n476_), .B2(new_n475_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n494_), .B1(new_n474_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n482_), .A2(new_n463_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n487_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n485_), .A2(new_n475_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n483_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n497_), .B1(new_n498_), .B2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(new_n493_), .B1(new_n496_), .B2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n479_), .A2(new_n488_), .A3(KEYINPUT30), .ZN(new_n503_));
  INV_X1    g302(.A(new_n451_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n502_), .A2(new_n503_), .A3(new_n504_), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n491_), .A2(new_n492_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n492_), .B1(new_n491_), .B2(new_n505_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n447_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n492_), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n489_), .A2(new_n490_), .A3(new_n451_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n504_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n509_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n491_), .A2(new_n492_), .A3(new_n505_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(KEYINPUT86), .A3(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n402_), .B(KEYINPUT31), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n515_), .B(KEYINPUT87), .Z(new_n516_));
  NAND3_X1  g315(.A1(new_n508_), .A2(new_n514_), .A3(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n515_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n518_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n517_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT88), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n517_), .A2(new_n522_), .A3(new_n519_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT93), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G78gat), .B(G106gat), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n526_));
  AND2_X1   g325(.A1(G197gat), .A2(G204gat), .ZN(new_n527_));
  NOR2_X1   g326(.A1(G197gat), .A2(G204gat), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT21), .ZN(new_n529_));
  NOR3_X1   g328(.A1(new_n527_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G211gat), .B(G218gat), .Z(new_n531_));
  NAND3_X1  g330(.A1(new_n530_), .A2(new_n531_), .A3(KEYINPUT90), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT90), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n359_), .A2(new_n292_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G197gat), .A2(G204gat), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(KEYINPUT21), .A3(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G211gat), .B(G218gat), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n533_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n532_), .A2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n529_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n540_), .A2(new_n536_), .A3(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(G228gat), .A2(G233gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT29), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n430_), .A2(new_n423_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n425_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n526_), .B1(new_n544_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT29), .B1(new_n420_), .B2(new_n425_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n550_), .A2(KEYINPUT91), .A3(new_n543_), .A4(new_n542_), .ZN(new_n551_));
  AND2_X1   g350(.A1(new_n549_), .A2(new_n551_), .ZN(new_n552_));
  AND2_X1   g351(.A1(new_n539_), .A2(new_n541_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n553_), .B1(new_n550_), .B2(KEYINPUT92), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT92), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n555_), .B(KEYINPUT29), .C1(new_n420_), .C2(new_n425_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n543_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n525_), .B1(new_n552_), .B2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT92), .B1(new_n431_), .B2(new_n545_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(new_n556_), .A3(new_n542_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n543_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n549_), .A2(new_n551_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n525_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n562_), .A2(new_n563_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n431_), .A2(new_n545_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT28), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(G22gat), .B(G50gat), .Z(new_n569_));
  NAND3_X1  g368(.A1(new_n431_), .A2(KEYINPUT28), .A3(new_n545_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n568_), .A2(new_n569_), .A3(new_n570_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n569_), .B1(new_n568_), .B2(new_n570_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  AND4_X1   g372(.A1(new_n524_), .A2(new_n558_), .A3(new_n565_), .A4(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n565_), .A2(KEYINPUT93), .ZN(new_n575_));
  AOI22_X1  g374(.A1(new_n575_), .A2(new_n573_), .B1(new_n558_), .B2(new_n565_), .ZN(new_n576_));
  NOR2_X1   g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G8gat), .B(G36gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT18), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(G64gat), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n580_), .A2(G92gat), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(G92gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  AND2_X1   g382(.A1(new_n457_), .A2(new_n459_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT26), .B(G190gat), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND4_X1  g385(.A1(new_n500_), .A2(new_n464_), .A3(new_n466_), .A4(new_n586_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n487_), .B1(new_n495_), .B2(new_n474_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n587_), .B1(new_n588_), .B2(new_n497_), .ZN(new_n589_));
  OR2_X1    g388(.A1(new_n589_), .A2(new_n542_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(G226gat), .A2(G233gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT19), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT20), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n479_), .A2(new_n488_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n594_), .B1(new_n595_), .B2(new_n542_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n590_), .A2(new_n593_), .A3(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n496_), .A2(new_n501_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n594_), .B1(new_n598_), .B2(new_n553_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n589_), .A2(new_n542_), .ZN(new_n600_));
  AOI21_X1  g399(.A(new_n593_), .B1(new_n599_), .B2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n583_), .B1(new_n597_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n599_), .A2(new_n600_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n592_), .ZN(new_n604_));
  AND2_X1   g403(.A1(new_n581_), .A2(new_n582_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n590_), .A2(new_n593_), .A3(new_n596_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n604_), .A2(new_n605_), .A3(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n433_), .A2(new_n434_), .A3(new_n436_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n426_), .A2(new_n432_), .A3(new_n437_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n608_), .A2(new_n399_), .A3(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT95), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT95), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n608_), .A2(new_n612_), .A3(new_n399_), .A4(new_n609_), .ZN(new_n613_));
  NAND4_X1  g412(.A1(new_n602_), .A2(new_n607_), .A3(new_n611_), .A4(new_n613_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n443_), .B1(new_n442_), .B2(new_n439_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  OAI211_X1 g416(.A(KEYINPUT33), .B(new_n443_), .C1(new_n442_), .C2(new_n439_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n581_), .A2(KEYINPUT32), .A3(new_n582_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n604_), .A2(new_n606_), .A3(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n621_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n589_), .A2(KEYINPUT96), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(new_n553_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n589_), .A2(KEYINPUT96), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n596_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(new_n592_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n599_), .A2(new_n593_), .A3(new_n600_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n620_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  OAI22_X1  g428(.A1(new_n614_), .A2(new_n619_), .B1(new_n622_), .B2(new_n629_), .ZN(new_n630_));
  AND4_X1   g429(.A1(new_n521_), .A2(new_n523_), .A3(new_n577_), .A4(new_n630_), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n574_), .A2(new_n576_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n521_), .A2(new_n632_), .A3(new_n523_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n577_), .A2(new_n520_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n627_), .A2(new_n628_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n583_), .B(KEYINPUT97), .ZN(new_n637_));
  OAI211_X1 g436(.A(KEYINPUT27), .B(new_n607_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(KEYINPUT27), .B1(new_n602_), .B2(new_n607_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT98), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(new_n640_), .ZN(new_n641_));
  AOI211_X1 g440(.A(KEYINPUT98), .B(KEYINPUT27), .C1(new_n602_), .C2(new_n607_), .ZN(new_n642_));
  OAI211_X1 g441(.A(new_n445_), .B(new_n638_), .C1(new_n641_), .C2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n643_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n631_), .B1(new_n635_), .B2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n352_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n276_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n226_), .A2(new_n228_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n230_), .B1(new_n648_), .B2(new_n219_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n217_), .A2(new_n218_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n259_), .B(new_n334_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(G232gat), .A2(G233gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT34), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n653_), .A2(KEYINPUT35), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND4_X1  g454(.A1(new_n647_), .A2(KEYINPUT71), .A3(new_n651_), .A4(new_n655_), .ZN(new_n656_));
  AND3_X1   g455(.A1(new_n231_), .A2(new_n334_), .A3(new_n259_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n352_), .B1(new_n231_), .B2(new_n259_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n653_), .A2(KEYINPUT35), .ZN(new_n659_));
  NOR3_X1   g458(.A1(new_n657_), .A2(new_n658_), .A3(new_n659_), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT71), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n654_), .B1(new_n651_), .B2(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n656_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(G218gat), .ZN(new_n664_));
  XNOR2_X1  g463(.A(G134gat), .B(G162gat), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT72), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(G190gat), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n665_), .B(KEYINPUT72), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n670_), .A2(G190gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n664_), .B1(new_n669_), .B2(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(G190gat), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n667_), .A2(new_n668_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n673_), .A2(new_n674_), .A3(G218gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT36), .B1(new_n672_), .B2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n663_), .A2(new_n676_), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n651_), .B1(new_n274_), .B2(new_n352_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT71), .B1(new_n274_), .B2(new_n334_), .ZN(new_n679_));
  OAI22_X1  g478(.A1(new_n678_), .A2(new_n659_), .B1(new_n679_), .B2(new_n654_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n672_), .A2(new_n675_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT36), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(new_n676_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n680_), .A2(new_n656_), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(KEYINPUT73), .B1(new_n677_), .B2(new_n685_), .ZN(new_n686_));
  AND2_X1   g485(.A1(new_n685_), .A2(KEYINPUT73), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT101), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n645_), .A2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n394_), .A2(new_n446_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G1gat), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT73), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n680_), .A2(new_n656_), .A3(new_n684_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n676_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n695_), .B1(new_n680_), .B2(new_n656_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n693_), .B1(new_n694_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT37), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n685_), .A2(KEYINPUT73), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n697_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT74), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n698_), .B1(new_n677_), .B2(new_n685_), .ZN(new_n702_));
  INV_X1    g501(.A(new_n702_), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n700_), .A2(new_n701_), .A3(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n701_), .B1(new_n700_), .B2(new_n703_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(new_n645_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n391_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n445_), .A2(G1gat), .ZN(new_n712_));
  AND3_X1   g511(.A1(new_n710_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n711_), .B1(new_n710_), .B2(new_n712_), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n692_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT102), .ZN(G1324gat));
  OR2_X1    g515(.A1(new_n641_), .A2(new_n642_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n638_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n392_), .A2(new_n718_), .A3(new_n690_), .A4(new_n393_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT39), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(new_n720_), .A3(G8gat), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n720_), .B1(new_n719_), .B2(G8gat), .ZN(new_n722_));
  INV_X1    g521(.A(new_n718_), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n723_), .A2(G8gat), .ZN(new_n724_));
  OAI22_X1  g523(.A1(new_n721_), .A2(new_n722_), .B1(new_n709_), .B2(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(KEYINPUT103), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT103), .ZN(new_n727_));
  OAI221_X1 g526(.A(new_n727_), .B1(new_n709_), .B2(new_n724_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n728_));
  AND3_X1   g527(.A1(new_n726_), .A2(KEYINPUT40), .A3(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(KEYINPUT40), .B1(new_n726_), .B2(new_n728_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n729_), .A2(new_n730_), .ZN(G1325gat));
  AND3_X1   g530(.A1(new_n517_), .A2(new_n522_), .A3(new_n519_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n522_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n710_), .A2(new_n316_), .A3(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n394_), .A2(new_n735_), .A3(new_n690_), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n737_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT41), .B1(new_n737_), .B2(G15gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n736_), .B1(new_n738_), .B2(new_n739_), .ZN(G1326gat));
  NAND3_X1  g539(.A1(new_n710_), .A2(new_n317_), .A3(new_n632_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n394_), .A2(new_n632_), .A3(new_n690_), .ZN(new_n742_));
  XOR2_X1   g541(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n743_));
  AND3_X1   g542(.A1(new_n742_), .A2(G22gat), .A3(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n742_), .B2(G22gat), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n741_), .B1(new_n744_), .B2(new_n745_), .ZN(G1327gat));
  INV_X1    g545(.A(new_n688_), .ZN(new_n747_));
  NOR3_X1   g546(.A1(new_n645_), .A2(new_n747_), .A3(new_n389_), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n302_), .A2(new_n307_), .A3(KEYINPUT13), .ZN(new_n749_));
  AOI21_X1  g548(.A(KEYINPUT13), .B1(new_n302_), .B2(new_n307_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n364_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n748_), .A2(new_n754_), .ZN(new_n755_));
  OR3_X1    g554(.A1(new_n755_), .A2(G29gat), .A3(new_n445_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT44), .ZN(new_n757_));
  NOR3_X1   g556(.A1(new_n686_), .A2(KEYINPUT37), .A3(new_n687_), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT74), .B1(new_n758_), .B2(new_n702_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n700_), .A2(new_n701_), .A3(new_n703_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n759_), .A2(new_n760_), .A3(new_n761_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n645_), .A2(new_n762_), .ZN(new_n763_));
  NOR3_X1   g562(.A1(new_n732_), .A2(new_n733_), .A3(new_n577_), .ZN(new_n764_));
  INV_X1    g563(.A(new_n634_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n644_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n631_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT106), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n704_), .A2(new_n705_), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT106), .B1(new_n759_), .B2(new_n761_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n768_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n763_), .B1(new_n772_), .B2(KEYINPUT43), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n387_), .A2(new_n388_), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n751_), .A2(new_n774_), .A3(new_n364_), .A4(new_n775_), .ZN(new_n776_));
  NAND4_X1  g575(.A1(new_n310_), .A2(new_n775_), .A3(new_n364_), .A4(new_n390_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT105), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n757_), .B1(new_n773_), .B2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n776_), .A2(new_n778_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n769_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n759_), .A2(KEYINPUT106), .A3(new_n761_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n760_), .B1(new_n784_), .B2(new_n768_), .ZN(new_n785_));
  OAI211_X1 g584(.A(KEYINPUT44), .B(new_n781_), .C1(new_n785_), .C2(new_n763_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n780_), .A2(new_n446_), .A3(new_n786_), .ZN(new_n787_));
  AND3_X1   g586(.A1(new_n787_), .A2(KEYINPUT107), .A3(G29gat), .ZN(new_n788_));
  AOI21_X1  g587(.A(KEYINPUT107), .B1(new_n787_), .B2(G29gat), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n756_), .B1(new_n788_), .B2(new_n789_), .ZN(G1328gat));
  NOR3_X1   g589(.A1(new_n755_), .A2(G36gat), .A3(new_n723_), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT45), .Z(new_n792_));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n793_));
  INV_X1    g592(.A(G36gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n781_), .B1(new_n785_), .B2(new_n763_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n723_), .B1(new_n795_), .B2(new_n757_), .ZN(new_n796_));
  AOI211_X1 g595(.A(new_n793_), .B(new_n794_), .C1(new_n796_), .C2(new_n786_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n780_), .A2(new_n718_), .A3(new_n786_), .ZN(new_n798_));
  AOI21_X1  g597(.A(KEYINPUT108), .B1(new_n798_), .B2(G36gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n792_), .B1(new_n797_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT46), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n800_), .A2(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n792_), .B(KEYINPUT46), .C1(new_n797_), .C2(new_n799_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(G1329gat));
  NAND4_X1  g603(.A1(new_n780_), .A2(G43gat), .A3(new_n520_), .A4(new_n786_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n755_), .A2(new_n734_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n805_), .B1(G43gat), .B2(new_n806_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(new_n807_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g607(.A1(new_n780_), .A2(new_n632_), .A3(new_n786_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n809_), .A2(KEYINPUT109), .A3(G50gat), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT109), .B1(new_n809_), .B2(G50gat), .ZN(new_n811_));
  NOR2_X1   g610(.A1(new_n577_), .A2(G50gat), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT110), .ZN(new_n813_));
  OAI22_X1  g612(.A1(new_n810_), .A2(new_n811_), .B1(new_n755_), .B2(new_n813_), .ZN(G1331gat));
  NOR2_X1   g613(.A1(new_n775_), .A2(new_n364_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n752_), .A2(new_n815_), .ZN(new_n816_));
  NOR3_X1   g615(.A1(new_n816_), .A2(new_n645_), .A3(new_n706_), .ZN(new_n817_));
  INV_X1    g616(.A(G57gat), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n817_), .A2(new_n818_), .A3(new_n446_), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n816_), .A2(new_n689_), .A3(new_n645_), .ZN(new_n820_));
  AND2_X1   g619(.A1(new_n820_), .A2(new_n446_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n821_), .B2(new_n818_), .ZN(G1332gat));
  INV_X1    g621(.A(G64gat), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n823_), .B1(new_n820_), .B2(new_n718_), .ZN(new_n824_));
  XOR2_X1   g623(.A(new_n824_), .B(KEYINPUT48), .Z(new_n825_));
  NAND2_X1  g624(.A1(new_n718_), .A2(new_n823_), .ZN(new_n826_));
  XOR2_X1   g625(.A(new_n826_), .B(KEYINPUT111), .Z(new_n827_));
  NAND2_X1  g626(.A1(new_n817_), .A2(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n825_), .A2(new_n828_), .ZN(G1333gat));
  INV_X1    g628(.A(G71gat), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n830_), .B1(new_n820_), .B2(new_n735_), .ZN(new_n831_));
  XOR2_X1   g630(.A(new_n831_), .B(KEYINPUT49), .Z(new_n832_));
  NAND3_X1  g631(.A1(new_n817_), .A2(new_n830_), .A3(new_n735_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(G1334gat));
  INV_X1    g633(.A(G78gat), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n835_), .B1(new_n820_), .B2(new_n632_), .ZN(new_n836_));
  XOR2_X1   g635(.A(new_n836_), .B(KEYINPUT50), .Z(new_n837_));
  NAND3_X1  g636(.A1(new_n817_), .A2(new_n835_), .A3(new_n632_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(new_n838_), .ZN(G1335gat));
  INV_X1    g638(.A(new_n773_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n751_), .A2(new_n364_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n775_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n840_), .A2(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(G85gat), .B1(new_n844_), .B2(new_n445_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n748_), .A2(new_n841_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(new_n253_), .A3(new_n446_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n845_), .A2(new_n848_), .ZN(G1336gat));
  OAI21_X1  g648(.A(G92gat), .B1(new_n844_), .B2(new_n723_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n847_), .A2(new_n254_), .A3(new_n718_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(G1337gat));
  NAND3_X1  g651(.A1(new_n840_), .A2(new_n735_), .A3(new_n843_), .ZN(new_n853_));
  AOI22_X1  g652(.A1(new_n517_), .A2(new_n519_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n854_));
  AOI22_X1  g653(.A1(new_n853_), .A2(G99gat), .B1(new_n847_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n856_), .A2(KEYINPUT113), .A3(KEYINPUT51), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT113), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT51), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n858_), .B1(new_n855_), .B2(new_n859_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT112), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n856_), .B2(KEYINPUT51), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n855_), .A2(KEYINPUT112), .A3(new_n859_), .ZN(new_n863_));
  OAI22_X1  g662(.A1(new_n857_), .A2(new_n860_), .B1(new_n862_), .B2(new_n863_), .ZN(G1338gat));
  INV_X1    g663(.A(KEYINPUT114), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n843_), .B(new_n632_), .C1(new_n785_), .C2(new_n763_), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(G106gat), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n866_), .A2(G106gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(KEYINPUT114), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n847_), .A2(new_n204_), .A3(new_n632_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n867_), .A2(new_n868_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n871_), .A2(new_n872_), .A3(new_n873_), .A4(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n870_), .A2(KEYINPUT114), .ZN(new_n876_));
  NOR3_X1   g675(.A1(new_n876_), .A2(new_n868_), .A3(new_n867_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n874_), .A2(new_n873_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT53), .B1(new_n877_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n875_), .A2(new_n879_), .ZN(G1339gat));
  NAND2_X1  g679(.A1(new_n723_), .A2(new_n446_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  AOI22_X1  g681(.A1(new_n305_), .A2(new_n306_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n284_), .B1(new_n279_), .B2(new_n275_), .ZN(new_n884_));
  OAI22_X1  g683(.A1(new_n280_), .A2(KEYINPUT55), .B1(new_n884_), .B2(new_n268_), .ZN(new_n885_));
  AND2_X1   g684(.A1(new_n280_), .A2(KEYINPUT55), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n296_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT115), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n887_), .A2(new_n888_), .A3(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n295_), .A2(new_n889_), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n891_), .B1(new_n885_), .B2(new_n886_), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(new_n893_), .ZN(new_n894_));
  OAI211_X1 g693(.A(KEYINPUT116), .B(new_n891_), .C1(new_n885_), .C2(new_n886_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n890_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n888_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n883_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(KEYINPUT117), .ZN(new_n899_));
  INV_X1    g698(.A(KEYINPUT117), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n900_), .B(new_n883_), .C1(new_n896_), .C2(new_n897_), .ZN(new_n901_));
  NAND3_X1  g700(.A1(new_n341_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n335_), .A2(new_n347_), .ZN(new_n903_));
  OAI211_X1 g702(.A(new_n902_), .B(new_n361_), .C1(new_n353_), .C2(new_n903_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n904_), .A2(new_n363_), .ZN(new_n905_));
  INV_X1    g704(.A(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n308_), .A2(new_n906_), .ZN(new_n907_));
  NAND3_X1  g706(.A1(new_n899_), .A2(new_n901_), .A3(new_n907_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n908_), .A2(new_n747_), .ZN(new_n909_));
  XOR2_X1   g708(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(new_n911_));
  AND2_X1   g710(.A1(new_n747_), .A2(KEYINPUT57), .ZN(new_n912_));
  AOI21_X1  g711(.A(new_n905_), .B1(new_n305_), .B2(new_n306_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n887_), .A2(new_n889_), .ZN(new_n914_));
  INV_X1    g713(.A(new_n892_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n913_), .B(KEYINPUT58), .C1(new_n914_), .C2(new_n915_), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT58), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n906_), .A2(new_n307_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n915_), .B1(new_n889_), .B2(new_n887_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n917_), .B1(new_n918_), .B2(new_n919_), .ZN(new_n920_));
  AND2_X1   g719(.A1(new_n916_), .A2(new_n920_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n908_), .A2(new_n912_), .B1(new_n921_), .B2(new_n706_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n389_), .B1(new_n911_), .B2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n751_), .A2(new_n815_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n706_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(KEYINPUT54), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n765_), .B(new_n882_), .C1(new_n923_), .C2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(KEYINPUT59), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n908_), .A2(new_n912_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n921_), .A2(new_n706_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n929_), .A2(new_n930_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n910_), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n932_), .B1(new_n908_), .B2(new_n747_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n775_), .B1(new_n931_), .B2(new_n933_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n925_), .B(new_n935_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n881_), .B1(new_n934_), .B2(new_n936_), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT59), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n937_), .A2(new_n938_), .A3(new_n765_), .ZN(new_n939_));
  NAND3_X1  g738(.A1(new_n928_), .A2(new_n939_), .A3(new_n364_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(G113gat), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT119), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n927_), .A2(new_n942_), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n937_), .A2(KEYINPUT119), .A3(new_n765_), .ZN(new_n944_));
  NOR2_X1   g743(.A1(new_n753_), .A2(G113gat), .ZN(new_n945_));
  NAND3_X1  g744(.A1(new_n943_), .A2(new_n944_), .A3(new_n945_), .ZN(new_n946_));
  NAND2_X1  g745(.A1(new_n941_), .A2(new_n946_), .ZN(G1340gat));
  NAND3_X1  g746(.A1(new_n928_), .A2(new_n939_), .A3(new_n752_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n948_), .A2(G120gat), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n751_), .A2(G120gat), .ZN(new_n950_));
  MUX2_X1   g749(.A(new_n950_), .B(G120gat), .S(KEYINPUT60), .Z(new_n951_));
  NAND3_X1  g750(.A1(new_n943_), .A2(new_n944_), .A3(new_n951_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n949_), .A2(new_n952_), .ZN(G1341gat));
  AND2_X1   g752(.A1(new_n928_), .A2(new_n939_), .ZN(new_n954_));
  INV_X1    g753(.A(G127gat), .ZN(new_n955_));
  NOR2_X1   g754(.A1(new_n775_), .A2(new_n955_), .ZN(new_n956_));
  XNOR2_X1  g755(.A(new_n956_), .B(KEYINPUT120), .ZN(new_n957_));
  NAND3_X1  g756(.A1(new_n943_), .A2(new_n944_), .A3(new_n389_), .ZN(new_n958_));
  AOI22_X1  g757(.A1(new_n954_), .A2(new_n957_), .B1(new_n958_), .B2(new_n955_), .ZN(G1342gat));
  NAND2_X1  g758(.A1(new_n706_), .A2(G134gat), .ZN(new_n960_));
  XOR2_X1   g759(.A(new_n960_), .B(KEYINPUT121), .Z(new_n961_));
  NAND3_X1  g760(.A1(new_n943_), .A2(new_n944_), .A3(new_n689_), .ZN(new_n962_));
  INV_X1    g761(.A(G134gat), .ZN(new_n963_));
  AOI22_X1  g762(.A1(new_n954_), .A2(new_n961_), .B1(new_n962_), .B2(new_n963_), .ZN(G1343gat));
  OAI211_X1 g763(.A(new_n764_), .B(new_n882_), .C1(new_n923_), .C2(new_n926_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n965_), .A2(new_n753_), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(new_n405_), .ZN(G1344gat));
  NOR2_X1   g766(.A1(new_n965_), .A2(new_n751_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n968_), .B(new_n406_), .ZN(G1345gat));
  OAI21_X1  g768(.A(KEYINPUT122), .B1(new_n965_), .B2(new_n775_), .ZN(new_n970_));
  INV_X1    g769(.A(KEYINPUT122), .ZN(new_n971_));
  NAND4_X1  g770(.A1(new_n937_), .A2(new_n971_), .A3(new_n764_), .A4(new_n389_), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n970_), .A2(new_n972_), .ZN(new_n973_));
  XNOR2_X1  g772(.A(KEYINPUT61), .B(G155gat), .ZN(new_n974_));
  INV_X1    g773(.A(new_n974_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n973_), .A2(new_n975_), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n970_), .A2(new_n972_), .A3(new_n974_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n976_), .A2(new_n977_), .ZN(G1346gat));
  INV_X1    g777(.A(new_n965_), .ZN(new_n979_));
  AOI21_X1  g778(.A(G162gat), .B1(new_n979_), .B2(new_n689_), .ZN(new_n980_));
  INV_X1    g779(.A(G162gat), .ZN(new_n981_));
  AOI21_X1  g780(.A(new_n981_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n982_));
  AOI21_X1  g781(.A(new_n980_), .B1(new_n979_), .B2(new_n982_), .ZN(G1347gat));
  NAND2_X1  g782(.A1(new_n934_), .A2(new_n936_), .ZN(new_n984_));
  NOR4_X1   g783(.A1(new_n723_), .A2(new_n446_), .A3(new_n734_), .A4(new_n632_), .ZN(new_n985_));
  NAND2_X1  g784(.A1(new_n984_), .A2(new_n985_), .ZN(new_n986_));
  INV_X1    g785(.A(new_n986_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n364_), .A2(new_n480_), .ZN(new_n988_));
  XOR2_X1   g787(.A(new_n988_), .B(KEYINPUT124), .Z(new_n989_));
  NAND2_X1  g788(.A1(new_n987_), .A2(new_n989_), .ZN(new_n990_));
  OAI211_X1 g789(.A(new_n364_), .B(new_n985_), .C1(new_n923_), .C2(new_n926_), .ZN(new_n991_));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n992_));
  NAND3_X1  g791(.A1(new_n991_), .A2(new_n992_), .A3(G169gat), .ZN(new_n993_));
  AOI21_X1  g792(.A(new_n992_), .B1(new_n991_), .B2(G169gat), .ZN(new_n994_));
  OAI21_X1  g793(.A(new_n993_), .B1(new_n994_), .B2(KEYINPUT123), .ZN(new_n995_));
  INV_X1    g794(.A(KEYINPUT123), .ZN(new_n996_));
  AOI211_X1 g795(.A(new_n996_), .B(new_n992_), .C1(new_n991_), .C2(G169gat), .ZN(new_n997_));
  OAI21_X1  g796(.A(new_n990_), .B1(new_n995_), .B2(new_n997_), .ZN(G1348gat));
  NOR2_X1   g797(.A1(new_n986_), .A2(new_n751_), .ZN(new_n999_));
  XNOR2_X1  g798(.A(new_n999_), .B(new_n481_), .ZN(G1349gat));
  INV_X1    g799(.A(KEYINPUT125), .ZN(new_n1001_));
  NAND3_X1  g800(.A1(new_n984_), .A2(new_n389_), .A3(new_n985_), .ZN(new_n1002_));
  OAI21_X1  g801(.A(new_n1001_), .B1(new_n1002_), .B2(new_n584_), .ZN(new_n1003_));
  NAND2_X1  g802(.A1(new_n1002_), .A2(new_n456_), .ZN(new_n1004_));
  NAND2_X1  g803(.A1(new_n1003_), .A2(new_n1004_), .ZN(new_n1005_));
  NOR3_X1   g804(.A1(new_n1002_), .A2(new_n1001_), .A3(new_n584_), .ZN(new_n1006_));
  NOR2_X1   g805(.A1(new_n1005_), .A2(new_n1006_), .ZN(G1350gat));
  NAND3_X1  g806(.A1(new_n987_), .A2(new_n689_), .A3(new_n585_), .ZN(new_n1008_));
  NAND3_X1  g807(.A1(new_n984_), .A2(new_n706_), .A3(new_n985_), .ZN(new_n1009_));
  AND3_X1   g808(.A1(new_n1009_), .A2(KEYINPUT126), .A3(G190gat), .ZN(new_n1010_));
  AOI21_X1  g809(.A(KEYINPUT126), .B1(new_n1009_), .B2(G190gat), .ZN(new_n1011_));
  OAI21_X1  g810(.A(new_n1008_), .B1(new_n1010_), .B2(new_n1011_), .ZN(G1351gat));
  NOR3_X1   g811(.A1(new_n723_), .A2(new_n446_), .A3(new_n633_), .ZN(new_n1013_));
  NAND2_X1  g812(.A1(new_n984_), .A2(new_n1013_), .ZN(new_n1014_));
  NOR2_X1   g813(.A1(new_n1014_), .A2(new_n753_), .ZN(new_n1015_));
  XNOR2_X1  g814(.A(new_n1015_), .B(new_n359_), .ZN(G1352gat));
  NOR2_X1   g815(.A1(new_n1014_), .A2(new_n751_), .ZN(new_n1017_));
  XNOR2_X1  g816(.A(new_n1017_), .B(new_n292_), .ZN(G1353gat));
  INV_X1    g817(.A(KEYINPUT63), .ZN(new_n1019_));
  AOI21_X1  g818(.A(new_n775_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1020_));
  OAI211_X1 g819(.A(new_n1013_), .B(new_n1020_), .C1(new_n923_), .C2(new_n926_), .ZN(new_n1021_));
  NAND2_X1  g820(.A1(new_n1021_), .A2(KEYINPUT127), .ZN(new_n1022_));
  INV_X1    g821(.A(G211gat), .ZN(new_n1023_));
  INV_X1    g822(.A(KEYINPUT127), .ZN(new_n1024_));
  NAND4_X1  g823(.A1(new_n984_), .A2(new_n1024_), .A3(new_n1013_), .A4(new_n1020_), .ZN(new_n1025_));
  AND4_X1   g824(.A1(new_n1019_), .A2(new_n1022_), .A3(new_n1023_), .A4(new_n1025_), .ZN(new_n1026_));
  AOI22_X1  g825(.A1(new_n1022_), .A2(new_n1025_), .B1(new_n1019_), .B2(new_n1023_), .ZN(new_n1027_));
  NOR2_X1   g826(.A1(new_n1026_), .A2(new_n1027_), .ZN(G1354gat));
  INV_X1    g827(.A(new_n706_), .ZN(new_n1029_));
  OAI21_X1  g828(.A(G218gat), .B1(new_n1014_), .B2(new_n1029_), .ZN(new_n1030_));
  NAND2_X1  g829(.A1(new_n689_), .A2(new_n664_), .ZN(new_n1031_));
  OAI21_X1  g830(.A(new_n1030_), .B1(new_n1014_), .B2(new_n1031_), .ZN(G1355gat));
endmodule


