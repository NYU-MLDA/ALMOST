//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n901_, new_n903_, new_n904_, new_n905_, new_n906_, new_n908_,
    new_n909_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n925_, new_n926_, new_n928_, new_n929_,
    new_n930_, new_n932_, new_n933_, new_n935_, new_n936_, new_n937_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_, new_n951_;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G169gat), .B(G197gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  XNOR2_X1  g004(.A(G29gat), .B(G36gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n206_), .B(G50gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT75), .B(G43gat), .ZN(new_n208_));
  XOR2_X1   g007(.A(new_n207_), .B(new_n208_), .Z(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT78), .B(G1gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G8gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT14), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G15gat), .B(G22gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(G1gat), .B(G8gat), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n212_), .A2(new_n213_), .A3(new_n215_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n209_), .A2(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n207_), .A2(new_n208_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n207_), .A2(new_n208_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n223_), .A2(new_n218_), .A3(new_n217_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n220_), .A2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G229gat), .A2(G233gat), .ZN(new_n226_));
  INV_X1    g025(.A(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n225_), .A2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT81), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT81), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n225_), .A2(new_n230_), .A3(new_n227_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT15), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n223_), .A2(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(KEYINPUT15), .B1(new_n221_), .B2(new_n222_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n226_), .B(new_n220_), .C1(new_n236_), .C2(new_n219_), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n205_), .B1(new_n232_), .B2(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n229_), .A2(new_n237_), .A3(new_n231_), .A4(new_n205_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n238_), .A2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(G85gat), .ZN(new_n242_));
  INV_X1    g041(.A(G92gat), .ZN(new_n243_));
  NOR3_X1   g042(.A1(new_n242_), .A2(new_n243_), .A3(KEYINPUT9), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT9), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n245_), .B1(G85gat), .B2(G92gat), .ZN(new_n246_));
  OAI22_X1  g045(.A1(new_n244_), .A2(new_n246_), .B1(G85gat), .B2(G92gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G99gat), .A2(G106gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n248_), .A2(KEYINPUT66), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n250_), .A2(G99gat), .A3(G106gat), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT6), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT67), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT6), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n249_), .A2(new_n251_), .A3(new_n253_), .A4(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n249_), .A2(new_n251_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(new_n255_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n247_), .A2(new_n256_), .A3(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT65), .B(G106gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT10), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(G99gat), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(G99gat), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n265_), .A2(KEYINPUT10), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n264_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(KEYINPUT64), .B1(new_n263_), .B2(new_n266_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n261_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n260_), .A2(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G71gat), .B(G78gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G57gat), .B(G64gat), .ZN(new_n275_));
  OR2_X1    g074(.A1(new_n275_), .A2(KEYINPUT11), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(KEYINPUT11), .ZN(new_n277_));
  AOI21_X1  g076(.A(new_n274_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n277_), .A2(new_n274_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  OR2_X1    g079(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n281_));
  NAND2_X1  g080(.A1(KEYINPUT68), .A2(KEYINPUT7), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(G106gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n265_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n283_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n282_), .A2(new_n265_), .A3(new_n284_), .ZN(new_n287_));
  NAND4_X1  g086(.A1(new_n259_), .A2(new_n286_), .A3(new_n287_), .A4(new_n256_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT69), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n287_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n285_), .B2(new_n283_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n292_), .A2(KEYINPUT69), .A3(new_n256_), .A4(new_n259_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT8), .ZN(new_n294_));
  XOR2_X1   g093(.A(G85gat), .B(G92gat), .Z(new_n295_));
  NAND4_X1  g094(.A1(new_n290_), .A2(new_n293_), .A3(new_n294_), .A4(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  AND3_X1   g096(.A1(new_n249_), .A2(new_n251_), .A3(KEYINPUT70), .ZN(new_n298_));
  AOI21_X1  g097(.A(KEYINPUT70), .B1(new_n249_), .B2(new_n251_), .ZN(new_n299_));
  OAI21_X1  g098(.A(KEYINPUT6), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n250_), .B1(G99gat), .B2(G106gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n248_), .A2(KEYINPUT66), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n301_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND3_X1  g103(.A1(new_n249_), .A2(new_n251_), .A3(KEYINPUT70), .ZN(new_n305_));
  NAND3_X1  g104(.A1(new_n304_), .A2(new_n252_), .A3(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(new_n300_), .A2(new_n306_), .A3(new_n292_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n294_), .B1(new_n307_), .B2(new_n295_), .ZN(new_n308_));
  OAI211_X1 g107(.A(new_n273_), .B(new_n280_), .C1(new_n297_), .C2(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n307_), .A2(new_n295_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n310_), .A2(KEYINPUT8), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n272_), .B1(new_n311_), .B2(new_n296_), .ZN(new_n312_));
  NOR3_X1   g111(.A1(new_n312_), .A2(KEYINPUT71), .A3(new_n280_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT71), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n273_), .B1(new_n297_), .B2(new_n308_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n280_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n314_), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n309_), .B1(new_n313_), .B2(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(G230gat), .A2(G233gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT12), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(new_n312_), .B2(new_n280_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n269_), .A2(new_n270_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n261_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n259_), .A2(new_n256_), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n325_), .A2(KEYINPUT73), .A3(new_n326_), .A4(new_n247_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n328_), .B1(new_n260_), .B2(new_n271_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n330_), .B1(new_n297_), .B2(new_n308_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n280_), .A2(new_n321_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n322_), .A2(new_n319_), .A3(new_n309_), .A4(new_n333_), .ZN(new_n334_));
  AOI22_X1  g133(.A1(new_n318_), .A2(new_n320_), .B1(new_n334_), .B2(KEYINPUT72), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT71), .B1(new_n312_), .B2(new_n280_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n315_), .A2(new_n314_), .A3(new_n316_), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n336_), .A2(new_n337_), .B1(new_n312_), .B2(new_n280_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT72), .ZN(new_n339_));
  NOR3_X1   g138(.A1(new_n338_), .A2(new_n339_), .A3(new_n319_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n335_), .A2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT5), .B(G176gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n342_), .B(G204gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(G120gat), .B(G148gat), .ZN(new_n344_));
  XOR2_X1   g143(.A(new_n343_), .B(new_n344_), .Z(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n341_), .A2(new_n346_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n335_), .B2(new_n340_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n347_), .A2(KEYINPUT13), .A3(new_n348_), .ZN(new_n349_));
  AOI21_X1  g148(.A(KEYINPUT13), .B1(new_n347_), .B2(new_n348_), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n351_), .A2(KEYINPUT74), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(KEYINPUT74), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n241_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT22), .B1(KEYINPUT87), .B2(G169gat), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT22), .ZN(new_n356_));
  OAI21_X1  g155(.A(G169gat), .B1(new_n356_), .B2(KEYINPUT86), .ZN(new_n357_));
  NAND2_X1  g156(.A1(KEYINPUT87), .A2(G169gat), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT86), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n355_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n361_));
  OR3_X1    g160(.A1(new_n361_), .A2(KEYINPUT88), .A3(G176gat), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G169gat), .A2(G176gat), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT88), .B1(new_n361_), .B2(G176gat), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(KEYINPUT89), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT23), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n367_), .B1(G183gat), .B2(G190gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n368_), .B(KEYINPUT90), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(G183gat), .A3(G190gat), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n371_), .B1(G183gat), .B2(G190gat), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT89), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n362_), .A2(new_n373_), .A3(new_n363_), .A4(new_n364_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n366_), .A2(new_n372_), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT30), .ZN(new_n376_));
  INV_X1    g175(.A(new_n370_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n377_), .A2(new_n368_), .ZN(new_n378_));
  INV_X1    g177(.A(G169gat), .ZN(new_n379_));
  INV_X1    g178(.A(G176gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n381_), .A2(KEYINPUT24), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n383_), .B(KEYINPUT85), .ZN(new_n384_));
  INV_X1    g183(.A(G190gat), .ZN(new_n385_));
  OR3_X1    g184(.A1(new_n385_), .A2(KEYINPUT82), .A3(KEYINPUT26), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT25), .B(G183gat), .ZN(new_n387_));
  OAI21_X1  g186(.A(KEYINPUT26), .B1(new_n385_), .B2(KEYINPUT82), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n386_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(KEYINPUT83), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n381_), .A2(KEYINPUT24), .A3(new_n363_), .ZN(new_n391_));
  XNOR2_X1  g190(.A(new_n391_), .B(KEYINPUT84), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n384_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n375_), .A2(new_n376_), .A3(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n376_), .B1(new_n375_), .B2(new_n393_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT92), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT92), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G227gat), .A2(G233gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(KEYINPUT91), .ZN(new_n401_));
  XOR2_X1   g200(.A(G15gat), .B(G43gat), .Z(new_n402_));
  XNOR2_X1  g201(.A(new_n401_), .B(new_n402_), .ZN(new_n403_));
  XOR2_X1   g202(.A(G71gat), .B(G99gat), .Z(new_n404_));
  XNOR2_X1  g203(.A(new_n403_), .B(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n397_), .A2(new_n399_), .A3(new_n406_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n396_), .A2(KEYINPUT92), .A3(new_n405_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT93), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G127gat), .B(G134gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G113gat), .B(G120gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n412_), .B(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT31), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n407_), .A2(KEYINPUT93), .A3(new_n408_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n411_), .A2(new_n416_), .A3(new_n417_), .ZN(new_n418_));
  XOR2_X1   g217(.A(G155gat), .B(G162gat), .Z(new_n419_));
  INV_X1    g218(.A(KEYINPUT1), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G141gat), .A2(G148gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT94), .ZN(new_n424_));
  INV_X1    g223(.A(G141gat), .ZN(new_n425_));
  INV_X1    g224(.A(G148gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NAND4_X1  g226(.A1(new_n421_), .A2(new_n422_), .A3(new_n424_), .A4(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT2), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(new_n430_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(KEYINPUT95), .A2(KEYINPUT3), .ZN(new_n432_));
  XNOR2_X1  g231(.A(new_n427_), .B(new_n432_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n431_), .B(new_n433_), .C1(new_n430_), .C2(new_n423_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n419_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT96), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n434_), .A2(KEYINPUT96), .A3(new_n419_), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n429_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n414_), .ZN(new_n440_));
  AND3_X1   g239(.A1(new_n434_), .A2(KEYINPUT96), .A3(new_n419_), .ZN(new_n441_));
  AOI21_X1  g240(.A(KEYINPUT96), .B1(new_n434_), .B2(new_n419_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n428_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n414_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n440_), .A2(new_n445_), .A3(KEYINPUT4), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT4), .ZN(new_n447_));
  NAND3_X1  g246(.A1(new_n443_), .A2(new_n447_), .A3(new_n444_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(KEYINPUT104), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G225gat), .A2(G233gat), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT104), .ZN(new_n452_));
  NAND4_X1  g251(.A1(new_n443_), .A2(new_n452_), .A3(new_n447_), .A4(new_n444_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n446_), .A2(new_n449_), .A3(new_n451_), .A4(new_n453_), .ZN(new_n454_));
  AND2_X1   g253(.A1(new_n440_), .A2(new_n445_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n450_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G1gat), .B(G29gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(G85gat), .ZN(new_n458_));
  XOR2_X1   g257(.A(KEYINPUT0), .B(G57gat), .Z(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n454_), .A2(new_n456_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n460_), .B1(new_n454_), .B2(new_n456_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n409_), .A2(new_n410_), .A3(new_n415_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n418_), .A2(new_n463_), .A3(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT107), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT29), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n439_), .A2(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(G22gat), .B(G50gat), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT28), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n469_), .B(new_n471_), .ZN(new_n472_));
  XOR2_X1   g271(.A(G78gat), .B(G106gat), .Z(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT97), .B1(new_n439_), .B2(new_n468_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G228gat), .A2(G233gat), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G197gat), .A2(G204gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT98), .B(G204gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  OAI211_X1 g277(.A(KEYINPUT21), .B(new_n476_), .C1(new_n478_), .C2(G197gat), .ZN(new_n479_));
  XOR2_X1   g278(.A(G211gat), .B(G218gat), .Z(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(G197gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(G204gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(new_n483_), .B1(new_n478_), .B2(new_n482_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n479_), .B(new_n481_), .C1(new_n484_), .C2(KEYINPUT21), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n484_), .A2(KEYINPUT21), .A3(new_n480_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT97), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n443_), .A2(new_n488_), .A3(KEYINPUT29), .ZN(new_n489_));
  NAND4_X1  g288(.A1(new_n474_), .A2(new_n475_), .A3(new_n487_), .A4(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n439_), .A2(new_n468_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT99), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n487_), .B(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(G228gat), .B(G233gat), .C1(new_n491_), .C2(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n473_), .B1(new_n490_), .B2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n472_), .B1(new_n495_), .B2(KEYINPUT100), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n490_), .A2(new_n494_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n473_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n490_), .A2(new_n494_), .A3(new_n473_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n496_), .A2(new_n501_), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n499_), .A2(KEYINPUT100), .A3(new_n500_), .A4(new_n472_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(G226gat), .A2(G233gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT19), .ZN(new_n507_));
  INV_X1    g306(.A(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n487_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n375_), .A2(new_n509_), .A3(new_n393_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT20), .ZN(new_n511_));
  XNOR2_X1  g310(.A(KEYINPUT22), .B(G169gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(new_n380_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n363_), .B(KEYINPUT101), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT102), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n513_), .A2(new_n514_), .A3(KEYINPUT102), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  OAI22_X1  g318(.A1(new_n377_), .A2(new_n368_), .B1(G183gat), .B2(G190gat), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT26), .B(G190gat), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n382_), .B1(new_n387_), .B2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n523_), .A2(new_n391_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n524_), .A2(new_n371_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n511_), .B1(new_n526_), .B2(new_n487_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n508_), .B1(new_n510_), .B2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G8gat), .B(G36gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(new_n243_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT18), .B(G64gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n509_), .B1(new_n375_), .B2(new_n393_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT103), .B1(new_n526_), .B2(new_n487_), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n519_), .A2(new_n520_), .B1(new_n524_), .B2(new_n371_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT103), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n509_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n536_), .A2(new_n539_), .A3(KEYINPUT20), .A4(new_n508_), .ZN(new_n540_));
  OAI211_X1 g339(.A(new_n529_), .B(new_n534_), .C1(new_n535_), .C2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n540_), .A2(new_n535_), .ZN(new_n542_));
  OAI21_X1  g341(.A(new_n533_), .B1(new_n542_), .B2(new_n528_), .ZN(new_n543_));
  AOI21_X1  g342(.A(KEYINPUT27), .B1(new_n541_), .B2(new_n543_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n542_), .A2(new_n533_), .A3(new_n528_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT106), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  NOR4_X1   g346(.A1(new_n542_), .A2(new_n528_), .A3(KEYINPUT106), .A4(new_n533_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n547_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT27), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n510_), .A2(new_n527_), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n551_), .A2(new_n507_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  AOI211_X1 g352(.A(new_n511_), .B(new_n535_), .C1(new_n493_), .C2(new_n537_), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n553_), .B1(new_n554_), .B2(new_n508_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n550_), .B1(new_n555_), .B2(new_n533_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n544_), .B1(new_n549_), .B2(new_n556_), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n467_), .B1(new_n505_), .B2(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n535_), .B1(new_n493_), .B2(new_n537_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n508_), .B1(new_n559_), .B2(KEYINPUT20), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n533_), .B1(new_n560_), .B2(new_n552_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n545_), .A2(new_n546_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n541_), .A2(KEYINPUT106), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n561_), .A2(new_n562_), .A3(new_n563_), .A4(KEYINPUT27), .ZN(new_n564_));
  INV_X1    g363(.A(new_n544_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n564_), .A2(new_n502_), .A3(new_n503_), .A4(new_n565_), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n566_), .A2(KEYINPUT107), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n466_), .B1(new_n558_), .B2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n418_), .A2(new_n464_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n504_), .A2(new_n463_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n564_), .A2(new_n565_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  NAND4_X1  g371(.A1(new_n446_), .A2(new_n449_), .A3(new_n450_), .A4(new_n453_), .ZN(new_n573_));
  OR2_X1    g372(.A1(new_n573_), .A2(KEYINPUT105), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(KEYINPUT105), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n460_), .B1(new_n455_), .B2(new_n451_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n543_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n578_), .A2(new_n545_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n461_), .A2(KEYINPUT33), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n454_), .A2(new_n456_), .A3(new_n460_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT33), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  NAND4_X1  g382(.A1(new_n577_), .A2(new_n579_), .A3(new_n580_), .A4(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(KEYINPUT32), .B(new_n534_), .C1(new_n560_), .C2(new_n552_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n542_), .A2(new_n528_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT32), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n586_), .B1(new_n587_), .B2(new_n533_), .ZN(new_n588_));
  OAI211_X1 g387(.A(new_n585_), .B(new_n588_), .C1(new_n461_), .C2(new_n462_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n504_), .B1(new_n584_), .B2(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n569_), .B1(new_n572_), .B2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n568_), .A2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n331_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n312_), .A2(new_n209_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT34), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n595_), .A2(KEYINPUT35), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(KEYINPUT35), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n597_), .A2(KEYINPUT35), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n593_), .A2(new_n599_), .A3(new_n600_), .A4(new_n594_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n598_), .A2(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G134gat), .B(G162gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(G218gat), .ZN(new_n604_));
  XOR2_X1   g403(.A(KEYINPUT76), .B(G190gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT36), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(KEYINPUT36), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n602_), .A2(new_n608_), .A3(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n598_), .A2(new_n601_), .A3(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n610_), .A2(KEYINPUT77), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n613_), .A3(KEYINPUT37), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT37), .ZN(new_n615_));
  OAI211_X1 g414(.A(new_n610_), .B(new_n611_), .C1(KEYINPUT77), .C2(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G231gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n219_), .B(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(new_n316_), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT79), .Z(new_n621_));
  XOR2_X1   g420(.A(G127gat), .B(G155gat), .Z(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(G211gat), .ZN(new_n623_));
  XOR2_X1   g422(.A(KEYINPUT16), .B(G183gat), .Z(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(KEYINPUT17), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n621_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n625_), .A2(KEYINPUT17), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n626_), .A2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n620_), .A2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT80), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n620_), .A2(KEYINPUT80), .A3(new_n629_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n627_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n617_), .A2(new_n634_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n354_), .A2(new_n592_), .A3(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT108), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n636_), .B(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n463_), .A2(new_n210_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n638_), .A2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT109), .B(KEYINPUT38), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  AND2_X1   g441(.A1(new_n354_), .A2(new_n592_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n612_), .B(KEYINPUT110), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n644_), .A2(new_n634_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n463_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G1gat), .ZN(new_n649_));
  INV_X1    g448(.A(new_n641_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n638_), .A2(new_n650_), .A3(new_n639_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n642_), .A2(new_n649_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT111), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  NAND4_X1  g453(.A1(new_n642_), .A2(KEYINPUT111), .A3(new_n649_), .A4(new_n651_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1324gat));
  INV_X1    g455(.A(G8gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n638_), .A2(new_n657_), .A3(new_n571_), .ZN(new_n658_));
  NAND4_X1  g457(.A1(new_n354_), .A2(new_n571_), .A3(new_n592_), .A4(new_n645_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(G8gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n660_), .B(KEYINPUT39), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(KEYINPUT112), .B(KEYINPUT40), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n662_), .B(new_n663_), .ZN(G1325gat));
  INV_X1    g463(.A(KEYINPUT41), .ZN(new_n665_));
  INV_X1    g464(.A(new_n569_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n646_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT113), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n667_), .A2(new_n668_), .A3(G15gat), .ZN(new_n669_));
  INV_X1    g468(.A(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n668_), .B1(new_n667_), .B2(G15gat), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n665_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n671_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n673_), .A2(KEYINPUT41), .A3(new_n669_), .ZN(new_n674_));
  OR3_X1    g473(.A1(new_n636_), .A2(G15gat), .A3(new_n569_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n672_), .A2(new_n674_), .A3(new_n675_), .ZN(G1326gat));
  INV_X1    g475(.A(G22gat), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n677_), .B1(new_n646_), .B2(new_n504_), .ZN(new_n678_));
  XOR2_X1   g477(.A(new_n678_), .B(KEYINPUT42), .Z(new_n679_));
  NAND2_X1  g478(.A1(new_n504_), .A2(new_n677_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n636_), .B2(new_n680_), .ZN(G1327gat));
  INV_X1    g480(.A(new_n634_), .ZN(new_n682_));
  NOR2_X1   g481(.A1(new_n682_), .A2(new_n612_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n643_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n647_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n584_), .A2(new_n589_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n505_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n557_), .A2(new_n463_), .A3(new_n504_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n666_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n505_), .A2(new_n557_), .A3(new_n467_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n566_), .A2(KEYINPUT107), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n465_), .B1(new_n691_), .B2(new_n692_), .ZN(new_n693_));
  OAI211_X1 g492(.A(new_n686_), .B(new_n617_), .C1(new_n690_), .C2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT114), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND4_X1  g495(.A1(new_n592_), .A2(KEYINPUT114), .A3(new_n686_), .A4(new_n617_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n617_), .B1(new_n690_), .B2(new_n693_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT43), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n696_), .A2(new_n697_), .A3(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n354_), .A2(new_n634_), .ZN(new_n701_));
  AND3_X1   g500(.A1(new_n700_), .A2(KEYINPUT44), .A3(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT44), .B1(new_n700_), .B2(new_n701_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n702_), .A2(new_n703_), .A3(new_n463_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n685_), .B1(new_n704_), .B2(G29gat), .ZN(G1328gat));
  INV_X1    g504(.A(G36gat), .ZN(new_n706_));
  NAND4_X1  g505(.A1(new_n643_), .A2(new_n706_), .A3(new_n571_), .A4(new_n683_), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n707_), .B(KEYINPUT45), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n702_), .A2(new_n703_), .A3(new_n557_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n708_), .B1(new_n709_), .B2(new_n706_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT46), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n708_), .B(KEYINPUT46), .C1(new_n709_), .C2(new_n706_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1329gat));
  NOR2_X1   g513(.A1(new_n702_), .A2(new_n703_), .ZN(new_n715_));
  INV_X1    g514(.A(G43gat), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n569_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n684_), .A2(new_n666_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(new_n716_), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n718_), .A2(KEYINPUT47), .A3(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT47), .B1(new_n718_), .B2(new_n720_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n721_), .A2(new_n722_), .ZN(G1330gat));
  AOI21_X1  g522(.A(G50gat), .B1(new_n684_), .B2(new_n504_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n504_), .A2(G50gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n715_), .B2(new_n725_), .ZN(G1331gat));
  NAND2_X1  g525(.A1(new_n352_), .A2(new_n353_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n241_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n729_), .A2(new_n592_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n730_), .A2(new_n645_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n731_), .A2(G57gat), .A3(new_n647_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n730_), .A2(new_n635_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n463_), .B1(new_n733_), .B2(KEYINPUT115), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(KEYINPUT115), .B2(new_n733_), .ZN(new_n735_));
  INV_X1    g534(.A(G57gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n732_), .B1(new_n735_), .B2(new_n736_), .ZN(G1332gat));
  INV_X1    g536(.A(G64gat), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n733_), .A2(new_n738_), .A3(new_n571_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n731_), .A2(new_n571_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(G64gat), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n741_), .A2(KEYINPUT48), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n741_), .A2(KEYINPUT48), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n739_), .B1(new_n742_), .B2(new_n743_), .ZN(G1333gat));
  INV_X1    g543(.A(G71gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n733_), .A2(new_n745_), .A3(new_n666_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n731_), .A2(new_n666_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G71gat), .ZN(new_n748_));
  AND2_X1   g547(.A1(new_n748_), .A2(KEYINPUT49), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n748_), .A2(KEYINPUT49), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(G1334gat));
  INV_X1    g550(.A(G78gat), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n733_), .A2(new_n752_), .A3(new_n504_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n731_), .A2(new_n504_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n754_), .A2(G78gat), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n755_), .A2(KEYINPUT50), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(KEYINPUT50), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(G1335gat));
  AND3_X1   g557(.A1(new_n700_), .A2(new_n634_), .A3(new_n729_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(new_n647_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(G85gat), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n730_), .A2(new_n683_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n762_), .A2(new_n242_), .A3(new_n647_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n761_), .A2(new_n763_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(KEYINPUT116), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT116), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n761_), .A2(new_n766_), .A3(new_n763_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1336gat));
  AOI21_X1  g567(.A(G92gat), .B1(new_n762_), .B2(new_n571_), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n557_), .A2(new_n243_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT117), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n759_), .B2(new_n771_), .ZN(G1337gat));
  NAND2_X1  g571(.A1(new_n759_), .A2(new_n666_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n569_), .B1(new_n270_), .B2(new_n269_), .ZN(new_n774_));
  AOI22_X1  g573(.A1(new_n773_), .A2(G99gat), .B1(new_n762_), .B2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT118), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(KEYINPUT51), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n775_), .B(new_n777_), .ZN(G1338gat));
  NAND3_X1  g577(.A1(new_n762_), .A2(new_n324_), .A3(new_n504_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n700_), .A2(new_n504_), .A3(new_n634_), .A4(new_n729_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(G106gat), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n781_), .B1(new_n780_), .B2(G106gat), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n779_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT53), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786_));
  OAI211_X1 g585(.A(new_n779_), .B(new_n786_), .C1(new_n782_), .C2(new_n783_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n785_), .A2(new_n787_), .ZN(G1339gat));
  NAND2_X1  g587(.A1(new_n209_), .A2(KEYINPUT15), .ZN(new_n789_));
  INV_X1    g588(.A(new_n235_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n219_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n220_), .ZN(new_n792_));
  OAI21_X1  g591(.A(KEYINPUT121), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT121), .ZN(new_n794_));
  OAI211_X1 g593(.A(new_n794_), .B(new_n220_), .C1(new_n236_), .C2(new_n219_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n793_), .A2(new_n795_), .A3(new_n227_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n225_), .A2(new_n226_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n796_), .A2(new_n204_), .A3(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(new_n239_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n799_), .B1(new_n341_), .B2(new_n346_), .ZN(new_n800_));
  AOI22_X1  g599(.A1(new_n332_), .A2(new_n331_), .B1(new_n312_), .B2(new_n280_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n319_), .B1(new_n801_), .B2(new_n322_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT55), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n334_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n801_), .A2(KEYINPUT55), .A3(new_n319_), .A4(new_n322_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT56), .B1(new_n806_), .B2(new_n345_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT56), .ZN(new_n808_));
  AOI211_X1 g607(.A(new_n808_), .B(new_n346_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n800_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT58), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n800_), .B(KEYINPUT58), .C1(new_n807_), .C2(new_n809_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n617_), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT122), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n812_), .A2(new_n617_), .A3(KEYINPUT122), .A4(new_n813_), .ZN(new_n817_));
  INV_X1    g616(.A(new_n612_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n311_), .A2(new_n296_), .B1(new_n329_), .B2(new_n327_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n332_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n309_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT12), .B1(new_n315_), .B2(new_n316_), .ZN(new_n822_));
  NOR3_X1   g621(.A1(new_n821_), .A2(new_n822_), .A3(new_n320_), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n320_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(KEYINPUT55), .B2(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(new_n805_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n345_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(KEYINPUT120), .A3(new_n808_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n346_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(KEYINPUT56), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(KEYINPUT56), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n828_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n241_), .B1(new_n341_), .B2(new_n346_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n347_), .A2(new_n348_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n799_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n818_), .B1(new_n835_), .B2(new_n838_), .ZN(new_n839_));
  AOI22_X1  g638(.A1(new_n816_), .A2(new_n817_), .B1(new_n839_), .B2(KEYINPUT57), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841_));
  AOI22_X1  g640(.A1(new_n833_), .A2(new_n834_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n841_), .B1(new_n842_), .B2(new_n818_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n682_), .B1(new_n840_), .B2(new_n843_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n635_), .A2(new_n351_), .A3(new_n241_), .ZN(new_n845_));
  AND2_X1   g644(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n846_));
  NOR2_X1   g645(.A1(KEYINPUT119), .A2(KEYINPUT54), .ZN(new_n847_));
  NOR2_X1   g646(.A1(new_n846_), .A2(new_n847_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n845_), .A2(new_n848_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n635_), .A2(new_n351_), .A3(new_n241_), .A4(new_n846_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n844_), .A2(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n691_), .A2(new_n692_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(new_n647_), .A3(new_n666_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n852_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(G113gat), .B1(new_n855_), .B2(new_n728_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n851_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n839_), .A2(KEYINPUT57), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n858_), .A2(new_n843_), .A3(new_n814_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(new_n634_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n857_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(KEYINPUT59), .ZN(new_n862_));
  INV_X1    g661(.A(new_n854_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(KEYINPUT123), .ZN(new_n865_));
  OAI21_X1  g664(.A(KEYINPUT59), .B1(new_n852_), .B2(new_n854_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT123), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n861_), .A2(new_n867_), .A3(new_n862_), .A4(new_n863_), .ZN(new_n868_));
  AND4_X1   g667(.A1(new_n728_), .A2(new_n865_), .A3(new_n866_), .A4(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n856_), .B1(new_n869_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g669(.A(new_n727_), .ZN(new_n871_));
  XOR2_X1   g670(.A(KEYINPUT124), .B(G120gat), .Z(new_n872_));
  AND2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  OAI221_X1 g672(.A(new_n863_), .B1(new_n873_), .B2(KEYINPUT60), .C1(new_n844_), .C2(new_n851_), .ZN(new_n874_));
  AND4_X1   g673(.A1(new_n866_), .A2(new_n865_), .A3(new_n868_), .A4(new_n874_), .ZN(new_n875_));
  OR2_X1    g674(.A1(new_n874_), .A2(KEYINPUT60), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n875_), .A2(new_n871_), .B1(new_n872_), .B2(new_n876_), .ZN(G1341gat));
  AOI21_X1  g676(.A(G127gat), .B1(new_n855_), .B2(new_n682_), .ZN(new_n878_));
  AND4_X1   g677(.A1(G127gat), .A2(new_n865_), .A3(new_n866_), .A4(new_n868_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n878_), .B1(new_n879_), .B2(new_n682_), .ZN(G1342gat));
  AOI21_X1  g679(.A(G134gat), .B1(new_n855_), .B2(new_n644_), .ZN(new_n881_));
  AND4_X1   g680(.A1(G134gat), .A2(new_n865_), .A3(new_n866_), .A4(new_n868_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n882_), .B2(new_n617_), .ZN(G1343gat));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n647_), .B(new_n569_), .C1(new_n844_), .C2(new_n851_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n505_), .A2(new_n571_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n884_), .B1(new_n885_), .B2(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n816_), .A2(new_n817_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n889_), .A2(new_n843_), .A3(new_n858_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(new_n634_), .ZN(new_n891_));
  AOI21_X1  g690(.A(new_n666_), .B1(new_n891_), .B2(new_n857_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n892_), .A2(KEYINPUT125), .A3(new_n647_), .A4(new_n886_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n888_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n894_), .A2(new_n728_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n895_), .A2(G141gat), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n894_), .A2(new_n425_), .A3(new_n728_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(G1344gat));
  NAND2_X1  g697(.A1(new_n894_), .A2(new_n871_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(G148gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n894_), .A2(new_n426_), .A3(new_n871_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n900_), .A2(new_n901_), .ZN(G1345gat));
  XNOR2_X1  g701(.A(KEYINPUT61), .B(G155gat), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n903_), .B1(new_n894_), .B2(new_n682_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n903_), .ZN(new_n905_));
  AOI211_X1 g704(.A(new_n634_), .B(new_n905_), .C1(new_n888_), .C2(new_n893_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n904_), .A2(new_n906_), .ZN(G1346gat));
  NAND2_X1  g706(.A1(new_n894_), .A2(new_n644_), .ZN(new_n908_));
  INV_X1    g707(.A(G162gat), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n909_), .B1(new_n888_), .B2(new_n893_), .ZN(new_n910_));
  AOI22_X1  g709(.A1(new_n908_), .A2(new_n909_), .B1(new_n910_), .B2(new_n617_), .ZN(G1347gat));
  NOR3_X1   g710(.A1(new_n465_), .A2(new_n504_), .A3(new_n557_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n913_), .B1(new_n857_), .B2(new_n860_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n379_), .B1(new_n914_), .B2(new_n728_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n914_), .A2(new_n728_), .A3(new_n512_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(KEYINPUT62), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n917_), .B1(new_n919_), .B2(new_n915_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(KEYINPUT126), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n922_));
  OAI211_X1 g721(.A(new_n917_), .B(new_n922_), .C1(new_n919_), .C2(new_n915_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n921_), .A2(new_n923_), .ZN(G1348gat));
  AOI21_X1  g723(.A(G176gat), .B1(new_n914_), .B2(new_n871_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n852_), .A2(new_n380_), .A3(new_n913_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n925_), .B1(new_n926_), .B2(new_n871_), .ZN(G1349gat));
  NOR2_X1   g726(.A1(new_n857_), .A2(new_n913_), .ZN(new_n928_));
  AOI21_X1  g727(.A(G183gat), .B1(new_n928_), .B2(new_n682_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n634_), .A2(new_n387_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n929_), .B1(new_n914_), .B2(new_n930_), .ZN(G1350gat));
  NAND3_X1  g730(.A1(new_n914_), .A2(new_n522_), .A3(new_n644_), .ZN(new_n932_));
  AND2_X1   g731(.A1(new_n914_), .A2(new_n617_), .ZN(new_n933_));
  OAI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(new_n385_), .ZN(G1351gat));
  NOR2_X1   g733(.A1(new_n570_), .A2(new_n557_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n892_), .A2(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n241_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(new_n482_), .ZN(G1352gat));
  NOR2_X1   g737(.A1(new_n936_), .A2(new_n727_), .ZN(new_n939_));
  MUX2_X1   g738(.A(G204gat), .B(new_n477_), .S(new_n939_), .Z(G1353gat));
  OAI22_X1  g739(.A1(new_n936_), .A2(new_n634_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n941_));
  XNOR2_X1  g740(.A(KEYINPUT63), .B(G211gat), .ZN(new_n942_));
  NAND4_X1  g741(.A1(new_n892_), .A2(new_n682_), .A3(new_n935_), .A4(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n944_), .A2(KEYINPUT127), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n946_));
  NAND3_X1  g745(.A1(new_n941_), .A2(new_n946_), .A3(new_n943_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n945_), .A2(new_n947_), .ZN(G1354gat));
  INV_X1    g747(.A(G218gat), .ZN(new_n949_));
  NOR2_X1   g748(.A1(new_n936_), .A2(new_n949_), .ZN(new_n950_));
  NAND3_X1  g749(.A1(new_n892_), .A2(new_n644_), .A3(new_n935_), .ZN(new_n951_));
  AOI22_X1  g750(.A1(new_n950_), .A2(new_n617_), .B1(new_n949_), .B2(new_n951_), .ZN(G1355gat));
endmodule


