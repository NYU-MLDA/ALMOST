//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:40 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n797_, new_n798_, new_n799_, new_n801_, new_n802_, new_n803_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_;
  INV_X1    g000(.A(KEYINPUT17), .ZN(new_n202_));
  XOR2_X1   g001(.A(G127gat), .B(G155gat), .Z(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT16), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G183gat), .B(G211gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G15gat), .B(G22gat), .ZN(new_n207_));
  INV_X1    g006(.A(G1gat), .ZN(new_n208_));
  INV_X1    g007(.A(G8gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(new_n208_), .B2(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n207_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G1gat), .B(G8gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n211_), .B(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G231gat), .A2(G233gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n213_), .B(new_n214_), .ZN(new_n215_));
  XNOR2_X1  g014(.A(G57gat), .B(G64gat), .ZN(new_n216_));
  OR2_X1    g015(.A1(new_n216_), .A2(KEYINPUT11), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(KEYINPUT11), .ZN(new_n218_));
  XOR2_X1   g017(.A(G71gat), .B(G78gat), .Z(new_n219_));
  NAND3_X1  g018(.A1(new_n217_), .A2(new_n218_), .A3(new_n219_), .ZN(new_n220_));
  OR2_X1    g019(.A1(new_n218_), .A2(new_n219_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n215_), .B(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT70), .ZN(new_n225_));
  AOI211_X1 g024(.A(new_n202_), .B(new_n206_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n226_), .B1(new_n225_), .B2(new_n224_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n206_), .B(new_n202_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT83), .ZN(new_n229_));
  AOI21_X1  g028(.A(new_n228_), .B1(new_n224_), .B2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n230_), .B1(new_n229_), .B2(new_n224_), .ZN(new_n231_));
  AND2_X1   g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(new_n232_), .B(KEYINPUT84), .ZN(new_n233_));
  INV_X1    g032(.A(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT7), .ZN(new_n235_));
  INV_X1    g034(.A(G99gat), .ZN(new_n236_));
  INV_X1    g035(.A(G106gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G99gat), .A2(G106gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n242_), .B(KEYINPUT6), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n241_), .A2(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT8), .ZN(new_n245_));
  XOR2_X1   g044(.A(G85gat), .B(G92gat), .Z(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n245_), .A3(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n248_));
  XNOR2_X1  g047(.A(KEYINPUT67), .B(KEYINPUT6), .ZN(new_n249_));
  OAI211_X1 g048(.A(new_n238_), .B(new_n239_), .C1(new_n249_), .C2(new_n242_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT6), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT67), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT6), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n252_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n242_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n248_), .B(new_n246_), .C1(new_n250_), .C2(new_n257_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n258_), .A2(KEYINPUT8), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n242_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n249_), .A2(new_n242_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n261_), .A2(new_n241_), .A3(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n248_), .B1(new_n263_), .B2(new_n246_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n247_), .B1(new_n259_), .B2(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(KEYINPUT10), .B(G99gat), .Z(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n237_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n267_), .B(KEYINPUT65), .ZN(new_n268_));
  XNOR2_X1  g067(.A(KEYINPUT66), .B(G85gat), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT9), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n269_), .A2(new_n270_), .A3(G92gat), .ZN(new_n271_));
  INV_X1    g070(.A(new_n246_), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n271_), .B(new_n243_), .C1(new_n270_), .C2(new_n272_), .ZN(new_n273_));
  OR2_X1    g072(.A1(new_n268_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n265_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n275_), .A2(new_n223_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n275_), .A2(new_n223_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT12), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(G230gat), .A2(G233gat), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT64), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n247_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n260_), .A2(new_n240_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n272_), .B1(new_n284_), .B2(new_n262_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n245_), .B1(new_n285_), .B2(new_n248_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n250_), .A2(new_n257_), .ZN(new_n287_));
  OAI21_X1  g086(.A(KEYINPUT68), .B1(new_n287_), .B2(new_n272_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n283_), .B1(new_n286_), .B2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(new_n268_), .A2(new_n273_), .ZN(new_n290_));
  OAI21_X1  g089(.A(KEYINPUT69), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n265_), .A2(new_n274_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n223_), .A2(new_n225_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n222_), .A2(KEYINPUT70), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n295_), .A2(KEYINPUT12), .A3(new_n296_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n279_), .B(new_n282_), .C1(new_n294_), .C2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n288_), .A2(KEYINPUT8), .A3(new_n258_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n290_), .B1(new_n299_), .B2(new_n247_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n222_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(new_n276_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n281_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n303_), .ZN(new_n304_));
  XOR2_X1   g103(.A(G120gat), .B(G148gat), .Z(new_n305_));
  XNOR2_X1  g104(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G176gat), .B(G204gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT72), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n304_), .A2(new_n310_), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n298_), .A2(new_n303_), .A3(new_n309_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(KEYINPUT73), .A2(KEYINPUT13), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n313_), .B1(new_n316_), .B2(new_n314_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(KEYINPUT81), .B(KEYINPUT37), .Z(new_n319_));
  XNOR2_X1  g118(.A(G29gat), .B(G36gat), .ZN(new_n320_));
  OR2_X1    g119(.A1(new_n320_), .A2(KEYINPUT76), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(KEYINPUT76), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  XNOR2_X1  g122(.A(G43gat), .B(G50gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n323_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n321_), .A2(new_n322_), .A3(new_n324_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n328_), .B(KEYINPUT15), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n291_), .A2(new_n293_), .A3(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G232gat), .A2(G233gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(new_n331_), .B(new_n332_), .ZN(new_n333_));
  XOR2_X1   g132(.A(KEYINPUT75), .B(KEYINPUT35), .Z(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n335_), .ZN(new_n336_));
  AOI22_X1  g135(.A1(new_n300_), .A2(new_n328_), .B1(new_n334_), .B2(new_n333_), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n330_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n336_), .B1(new_n330_), .B2(new_n337_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n341_));
  XOR2_X1   g140(.A(G190gat), .B(G218gat), .Z(new_n342_));
  XNOR2_X1  g141(.A(G134gat), .B(G162gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT36), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(new_n346_), .B(KEYINPUT77), .Z(new_n347_));
  NAND3_X1  g146(.A1(new_n340_), .A2(new_n341_), .A3(new_n347_), .ZN(new_n348_));
  AND3_X1   g147(.A1(new_n265_), .A2(new_n274_), .A3(new_n292_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n292_), .B1(new_n265_), .B2(new_n274_), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT15), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n328_), .B(new_n351_), .ZN(new_n352_));
  NOR3_X1   g151(.A1(new_n349_), .A2(new_n350_), .A3(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n300_), .A2(new_n328_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n333_), .A2(new_n334_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n335_), .B1(new_n353_), .B2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n330_), .A2(new_n336_), .A3(new_n337_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(new_n358_), .A3(new_n347_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT78), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n319_), .B1(new_n348_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n357_), .A2(KEYINPUT79), .A3(new_n358_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n344_), .B(KEYINPUT36), .ZN(new_n366_));
  AOI21_X1  g165(.A(KEYINPUT80), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT80), .ZN(new_n368_));
  INV_X1    g167(.A(new_n366_), .ZN(new_n369_));
  AOI211_X1 g168(.A(new_n368_), .B(new_n369_), .C1(new_n363_), .C2(new_n364_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n361_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n348_), .A2(new_n360_), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n366_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT37), .ZN(new_n376_));
  AND3_X1   g175(.A1(new_n371_), .A2(new_n372_), .A3(new_n376_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n372_), .B1(new_n371_), .B2(new_n376_), .ZN(new_n378_));
  OAI211_X1 g177(.A(new_n234_), .B(new_n318_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT85), .ZN(new_n380_));
  OR2_X1    g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n379_), .A2(new_n380_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(G227gat), .A2(G233gat), .ZN(new_n383_));
  XOR2_X1   g182(.A(new_n383_), .B(KEYINPUT90), .Z(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT30), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(KEYINPUT31), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G15gat), .B(G43gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n388_), .B(KEYINPUT89), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n389_), .B(G71gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(G99gat), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n392_), .B1(G183gat), .B2(G190gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G183gat), .A2(G190gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(KEYINPUT88), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT88), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n396_), .A2(G183gat), .A3(G190gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n395_), .A2(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n393_), .B1(new_n398_), .B2(new_n392_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(KEYINPUT25), .B(G183gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT26), .B(G190gat), .ZN(new_n401_));
  AND2_X1   g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  NOR3_X1   g201(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n399_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(G169gat), .ZN(new_n405_));
  INV_X1    g204(.A(G176gat), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT24), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(G169gat), .A2(G176gat), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT87), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT24), .ZN(new_n410_));
  AOI21_X1  g209(.A(new_n410_), .B1(G169gat), .B2(G176gat), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT87), .ZN(new_n412_));
  INV_X1    g211(.A(new_n408_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n411_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n394_), .A2(new_n392_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n398_), .B2(KEYINPUT23), .ZN(new_n418_));
  NOR2_X1   g217(.A1(G183gat), .A2(G190gat), .ZN(new_n419_));
  INV_X1    g218(.A(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n418_), .A2(new_n420_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(G169gat), .ZN(new_n423_));
  AOI22_X1  g222(.A1(new_n404_), .A2(new_n415_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n391_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n390_), .B(new_n236_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n399_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n403_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n415_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n421_), .A2(new_n423_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(G127gat), .B(G134gat), .Z(new_n433_));
  XOR2_X1   g232(.A(G113gat), .B(G120gat), .Z(new_n434_));
  XOR2_X1   g233(.A(new_n433_), .B(new_n434_), .Z(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  AND3_X1   g235(.A1(new_n425_), .A2(new_n432_), .A3(new_n436_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n436_), .B1(new_n425_), .B2(new_n432_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n387_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n425_), .A2(new_n432_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n440_), .A2(new_n435_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n425_), .A2(new_n432_), .A3(new_n436_), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n441_), .A2(new_n386_), .A3(new_n442_), .ZN(new_n443_));
  AND2_X1   g242(.A1(new_n439_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  XOR2_X1   g244(.A(G22gat), .B(G50gat), .Z(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G141gat), .A2(G148gat), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT92), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n450_), .A2(KEYINPUT2), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT2), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n448_), .A2(new_n449_), .A3(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT91), .ZN(new_n454_));
  OAI22_X1  g253(.A1(new_n454_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n455_));
  NOR2_X1   g254(.A1(G141gat), .A2(G148gat), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT3), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n456_), .A2(KEYINPUT91), .A3(new_n457_), .ZN(new_n458_));
  NAND4_X1  g257(.A1(new_n451_), .A2(new_n453_), .A3(new_n455_), .A4(new_n458_), .ZN(new_n459_));
  OR2_X1    g258(.A1(G155gat), .A2(G162gat), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G155gat), .A2(G162gat), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n459_), .A2(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT29), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT1), .ZN(new_n465_));
  NOR2_X1   g264(.A1(new_n461_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n448_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n466_), .A2(new_n467_), .A3(new_n456_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n460_), .A2(new_n465_), .A3(new_n461_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n463_), .A2(new_n464_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT28), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT93), .ZN(new_n473_));
  AOI22_X1  g272(.A1(new_n459_), .A2(new_n462_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT28), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n474_), .A2(new_n475_), .A3(new_n464_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n472_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n473_), .B1(new_n472_), .B2(new_n476_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n447_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n476_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n475_), .B1(new_n474_), .B2(new_n464_), .ZN(new_n481_));
  OAI21_X1  g280(.A(KEYINPUT93), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n472_), .A2(new_n473_), .A3(new_n476_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n482_), .A2(new_n446_), .A3(new_n483_), .ZN(new_n484_));
  AND2_X1   g283(.A1(new_n479_), .A2(new_n484_), .ZN(new_n485_));
  OR2_X1    g284(.A1(new_n485_), .A2(KEYINPUT98), .ZN(new_n486_));
  XOR2_X1   g285(.A(G211gat), .B(G218gat), .Z(new_n487_));
  INV_X1    g286(.A(KEYINPUT21), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G197gat), .B(G204gat), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n487_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(G204gat), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n491_), .A2(KEYINPUT96), .A3(G197gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(G197gat), .ZN(new_n493_));
  INV_X1    g292(.A(G197gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n494_), .A2(G204gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  OAI211_X1 g295(.A(KEYINPUT21), .B(new_n492_), .C1(new_n496_), .C2(KEYINPUT96), .ZN(new_n497_));
  NOR2_X1   g296(.A1(new_n489_), .A2(new_n488_), .ZN(new_n498_));
  AOI22_X1  g297(.A1(new_n490_), .A2(new_n497_), .B1(new_n487_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n463_), .A2(new_n470_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n499_), .B1(KEYINPUT29), .B2(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(KEYINPUT94), .A2(G228gat), .ZN(new_n502_));
  NOR2_X1   g301(.A1(KEYINPUT94), .A2(G228gat), .ZN(new_n503_));
  OAI21_X1  g302(.A(G233gat), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT95), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n501_), .A2(new_n505_), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n506_), .B(KEYINPUT97), .C1(new_n501_), .C2(new_n504_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(KEYINPUT97), .B2(new_n506_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n479_), .A2(new_n484_), .A3(KEYINPUT98), .ZN(new_n509_));
  XOR2_X1   g308(.A(G78gat), .B(G106gat), .Z(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  AND3_X1   g310(.A1(new_n508_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n511_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n486_), .B1(new_n512_), .B2(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n508_), .A2(new_n509_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(new_n510_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n485_), .A2(KEYINPUT98), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n508_), .A2(new_n509_), .A3(new_n511_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n516_), .A2(new_n517_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n514_), .A2(new_n519_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(G8gat), .B(G36gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n521_), .B(KEYINPUT18), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G64gat), .B(G92gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n522_), .B(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G226gat), .A2(G233gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(KEYINPUT19), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n499_), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT20), .B1(new_n431_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n403_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT101), .B1(new_n418_), .B2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT26), .ZN(new_n532_));
  NOR2_X1   g331(.A1(new_n532_), .A2(G190gat), .ZN(new_n533_));
  INV_X1    g332(.A(G190gat), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n534_), .A2(KEYINPUT26), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT99), .B1(new_n533_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(KEYINPUT26), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n532_), .A2(G190gat), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT99), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n537_), .A2(new_n538_), .A3(new_n539_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n536_), .A2(new_n400_), .A3(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT100), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n407_), .A2(new_n542_), .ZN(new_n543_));
  OAI211_X1 g342(.A(KEYINPUT100), .B(KEYINPUT24), .C1(new_n405_), .C2(new_n406_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n413_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n541_), .A2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n392_), .B1(new_n395_), .B2(new_n397_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT101), .ZN(new_n548_));
  NOR4_X1   g347(.A1(new_n547_), .A2(new_n417_), .A3(new_n548_), .A4(new_n403_), .ZN(new_n549_));
  NOR3_X1   g348(.A1(new_n531_), .A2(new_n546_), .A3(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n423_), .B1(new_n399_), .B2(new_n419_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n528_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n553_));
  AOI21_X1  g352(.A(new_n529_), .B1(new_n553_), .B2(KEYINPUT102), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT102), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n555_), .B(new_n528_), .C1(new_n550_), .C2(new_n552_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n527_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT20), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n558_), .B1(new_n431_), .B2(new_n528_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n398_), .A2(KEYINPUT23), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n560_), .A2(new_n416_), .A3(new_n530_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(new_n548_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n418_), .A2(KEYINPUT101), .A3(new_n530_), .ZN(new_n563_));
  NAND4_X1  g362(.A1(new_n562_), .A2(new_n563_), .A3(new_n541_), .A4(new_n545_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n564_), .A2(new_n499_), .A3(new_n551_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n559_), .A2(new_n565_), .A3(new_n527_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n524_), .B1(new_n557_), .B2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n558_), .B1(new_n424_), .B2(new_n499_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n499_), .B1(new_n564_), .B2(new_n551_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n569_), .B1(new_n570_), .B2(new_n555_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n556_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n526_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n524_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n573_), .A2(new_n574_), .A3(new_n566_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n568_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT27), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n531_), .A2(new_n546_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n552_), .B1(new_n578_), .B2(new_n563_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT102), .B1(new_n579_), .B2(new_n499_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n580_), .A2(new_n556_), .A3(new_n569_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n567_), .B1(new_n581_), .B2(new_n526_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n577_), .B1(new_n582_), .B2(new_n574_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n559_), .A2(new_n565_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n526_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n585_), .B1(new_n581_), .B2(new_n526_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(new_n524_), .ZN(new_n587_));
  AOI22_X1  g386(.A1(new_n576_), .A2(new_n577_), .B1(new_n583_), .B2(new_n587_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n520_), .A2(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n435_), .A2(new_n500_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT4), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n436_), .A2(new_n474_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n593_), .A2(KEYINPUT103), .A3(new_n590_), .ZN(new_n594_));
  OR3_X1    g393(.A1(new_n435_), .A2(new_n500_), .A3(KEYINPUT103), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n592_), .B1(new_n596_), .B2(new_n591_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(G225gat), .A2(G233gat), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n596_), .A2(new_n598_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(G1gat), .B(G29gat), .Z(new_n603_));
  XNOR2_X1  g402(.A(G57gat), .B(G85gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT104), .B(KEYINPUT0), .ZN(new_n606_));
  XOR2_X1   g405(.A(new_n605_), .B(new_n606_), .Z(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n607_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n600_), .A2(new_n609_), .A3(new_n601_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n589_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(KEYINPUT105), .A2(KEYINPUT33), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n576_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n610_), .A2(new_n613_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n609_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n596_), .B(KEYINPUT106), .Z(new_n618_));
  OAI21_X1  g417(.A(new_n617_), .B1(new_n618_), .B2(new_n598_), .ZN(new_n619_));
  NAND4_X1  g418(.A1(new_n614_), .A2(new_n615_), .A3(new_n616_), .A4(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT32), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n582_), .B1(new_n621_), .B2(new_n524_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n586_), .A2(KEYINPUT32), .A3(new_n574_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n611_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  AOI21_X1  g423(.A(new_n520_), .B1(new_n620_), .B2(new_n624_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n445_), .B1(new_n612_), .B2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(KEYINPUT108), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT107), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n557_), .A2(new_n524_), .A3(new_n567_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n574_), .B1(new_n573_), .B2(new_n566_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n577_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n587_), .A2(new_n575_), .A3(KEYINPUT27), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n631_), .A2(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n628_), .B1(new_n520_), .B2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n588_), .A2(KEYINPUT107), .A3(new_n519_), .A4(new_n514_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n608_), .A2(new_n610_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n637_), .A2(new_n444_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n627_), .B1(new_n636_), .B2(new_n639_), .ZN(new_n640_));
  AOI211_X1 g439(.A(KEYINPUT108), .B(new_n638_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n626_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n329_), .A2(new_n213_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n213_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n328_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G229gat), .A2(G233gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n643_), .A2(new_n645_), .A3(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n328_), .B(new_n644_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n646_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n647_), .A2(new_n650_), .ZN(new_n651_));
  XOR2_X1   g450(.A(G113gat), .B(G141gat), .Z(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT86), .ZN(new_n653_));
  XOR2_X1   g452(.A(G169gat), .B(G197gat), .Z(new_n654_));
  XNOR2_X1  g453(.A(new_n653_), .B(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(new_n651_), .B(new_n655_), .Z(new_n656_));
  AND2_X1   g455(.A1(new_n642_), .A2(new_n656_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n381_), .A2(new_n382_), .A3(new_n657_), .ZN(new_n658_));
  INV_X1    g457(.A(KEYINPUT109), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND4_X1  g459(.A1(new_n381_), .A2(KEYINPUT109), .A3(new_n382_), .A4(new_n657_), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n637_), .A2(G1gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT110), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT110), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n660_), .A2(new_n665_), .A3(new_n661_), .A4(new_n662_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT38), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n373_), .B1(new_n367_), .B2(new_n370_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n642_), .A2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT112), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n318_), .A2(new_n656_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n232_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT111), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n672_), .A2(new_n611_), .A3(new_n676_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(G1gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n664_), .A2(KEYINPUT38), .A3(new_n666_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n669_), .A2(new_n678_), .A3(new_n679_), .ZN(G1324gat));
  NAND4_X1  g479(.A1(new_n660_), .A2(new_n209_), .A3(new_n633_), .A4(new_n661_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n672_), .A2(new_n633_), .A3(new_n676_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT39), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n682_), .A2(new_n683_), .A3(G8gat), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n683_), .B1(new_n682_), .B2(G8gat), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT40), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  OAI211_X1 g487(.A(KEYINPUT40), .B(new_n681_), .C1(new_n684_), .C2(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n688_), .A2(new_n689_), .ZN(G1325gat));
  AND2_X1   g489(.A1(new_n660_), .A2(new_n661_), .ZN(new_n691_));
  INV_X1    g490(.A(G15gat), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(new_n692_), .A3(new_n444_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n672_), .A2(new_n444_), .A3(new_n676_), .ZN(new_n694_));
  AND3_X1   g493(.A1(new_n694_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT41), .B1(new_n694_), .B2(G15gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n693_), .B1(new_n695_), .B2(new_n696_), .ZN(G1326gat));
  INV_X1    g496(.A(G22gat), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n691_), .A2(new_n698_), .A3(new_n520_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n672_), .A2(new_n520_), .A3(new_n676_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(G22gat), .ZN(new_n701_));
  AND2_X1   g500(.A1(new_n701_), .A2(KEYINPUT42), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n701_), .A2(KEYINPUT42), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(G1327gat));
  INV_X1    g503(.A(new_n670_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n705_), .A2(new_n233_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n318_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n657_), .A2(new_n708_), .ZN(new_n709_));
  OR3_X1    g508(.A1(new_n709_), .A2(G29gat), .A3(new_n637_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n673_), .A2(new_n234_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n377_), .A2(new_n378_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n642_), .A2(new_n712_), .A3(new_n713_), .ZN(new_n714_));
  AOI21_X1  g513(.A(new_n713_), .B1(new_n642_), .B2(new_n712_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n711_), .B1(new_n714_), .B2(new_n715_), .ZN(new_n716_));
  INV_X1    g515(.A(KEYINPUT44), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n716_), .A2(new_n717_), .ZN(new_n718_));
  OAI211_X1 g517(.A(KEYINPUT44), .B(new_n711_), .C1(new_n714_), .C2(new_n715_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n720_), .A2(KEYINPUT113), .A3(new_n611_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(G29gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(KEYINPUT113), .B1(new_n720_), .B2(new_n611_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n710_), .B1(new_n722_), .B2(new_n723_), .ZN(G1328gat));
  NAND3_X1  g523(.A1(new_n718_), .A2(new_n633_), .A3(new_n719_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(G36gat), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n588_), .A2(G36gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n657_), .A2(new_n708_), .A3(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT45), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(new_n730_));
  INV_X1    g529(.A(new_n730_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n726_), .A2(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT46), .B1(new_n732_), .B2(KEYINPUT114), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n730_), .B1(new_n725_), .B2(G36gat), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT114), .ZN(new_n735_));
  INV_X1    g534(.A(KEYINPUT46), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n734_), .A2(new_n735_), .A3(new_n736_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n733_), .A2(new_n737_), .ZN(G1329gat));
  NOR3_X1   g537(.A1(new_n709_), .A2(G43gat), .A3(new_n445_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n720_), .A2(new_n444_), .ZN(new_n741_));
  INV_X1    g540(.A(G43gat), .ZN(new_n742_));
  OAI211_X1 g541(.A(KEYINPUT47), .B(new_n740_), .C1(new_n741_), .C2(new_n742_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT47), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n742_), .B1(new_n720_), .B2(new_n444_), .ZN(new_n745_));
  OAI21_X1  g544(.A(new_n744_), .B1(new_n745_), .B2(new_n739_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n743_), .A2(new_n746_), .ZN(G1330gat));
  NAND2_X1  g546(.A1(new_n720_), .A2(new_n520_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n748_), .A2(G50gat), .ZN(new_n749_));
  INV_X1    g548(.A(new_n520_), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n750_), .A2(G50gat), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT115), .Z(new_n752_));
  OAI21_X1  g551(.A(new_n749_), .B1(new_n709_), .B2(new_n752_), .ZN(G1331gat));
  NOR2_X1   g552(.A1(new_n233_), .A2(new_n656_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n672_), .A2(new_n707_), .A3(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(G57gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n757_), .B1(new_n611_), .B2(KEYINPUT117), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n758_), .B1(KEYINPUT117), .B2(new_n757_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n712_), .A2(new_n233_), .A3(new_n318_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n656_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n642_), .A2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n637_), .B1(new_n763_), .B2(KEYINPUT116), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n764_), .B1(KEYINPUT116), .B2(new_n763_), .ZN(new_n765_));
  AOI22_X1  g564(.A1(new_n756_), .A2(new_n759_), .B1(new_n765_), .B2(new_n757_), .ZN(G1332gat));
  INV_X1    g565(.A(new_n763_), .ZN(new_n767_));
  INV_X1    g566(.A(G64gat), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n767_), .A2(new_n768_), .A3(new_n633_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT48), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n756_), .A2(new_n633_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n770_), .B1(new_n771_), .B2(G64gat), .ZN(new_n772_));
  AOI211_X1 g571(.A(KEYINPUT48), .B(new_n768_), .C1(new_n756_), .C2(new_n633_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n769_), .B1(new_n772_), .B2(new_n773_), .ZN(G1333gat));
  OR3_X1    g573(.A1(new_n763_), .A2(G71gat), .A3(new_n445_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n756_), .A2(new_n444_), .ZN(new_n776_));
  XOR2_X1   g575(.A(KEYINPUT118), .B(KEYINPUT49), .Z(new_n777_));
  AND3_X1   g576(.A1(new_n776_), .A2(G71gat), .A3(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n777_), .B1(new_n776_), .B2(G71gat), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(G1334gat));
  INV_X1    g579(.A(G78gat), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n767_), .A2(new_n781_), .A3(new_n520_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n756_), .A2(new_n520_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(G78gat), .ZN(new_n785_));
  AOI211_X1 g584(.A(KEYINPUT50), .B(new_n781_), .C1(new_n756_), .C2(new_n520_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n782_), .B1(new_n785_), .B2(new_n786_), .ZN(G1335gat));
  NAND4_X1  g586(.A1(new_n762_), .A2(new_n233_), .A3(new_n707_), .A4(new_n705_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT119), .ZN(new_n789_));
  XNOR2_X1  g588(.A(new_n788_), .B(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(G85gat), .B1(new_n790_), .B2(new_n611_), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n714_), .A2(new_n715_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n234_), .A2(new_n318_), .A3(new_n656_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n611_), .A2(new_n269_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n791_), .B1(new_n794_), .B2(new_n795_), .ZN(G1336gat));
  AOI21_X1  g595(.A(G92gat), .B1(new_n790_), .B2(new_n633_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n633_), .A2(G92gat), .ZN(new_n798_));
  XOR2_X1   g597(.A(new_n798_), .B(KEYINPUT120), .Z(new_n799_));
  AOI21_X1  g598(.A(new_n797_), .B1(new_n794_), .B2(new_n799_), .ZN(G1337gat));
  NAND2_X1  g599(.A1(new_n794_), .A2(new_n444_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(G99gat), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n790_), .A2(new_n266_), .A3(new_n444_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n802_), .A2(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(KEYINPUT51), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT51), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n802_), .A2(new_n806_), .A3(new_n803_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n805_), .A2(new_n807_), .ZN(G1338gat));
  NAND3_X1  g607(.A1(new_n790_), .A2(new_n237_), .A3(new_n520_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n792_), .A2(new_n520_), .A3(new_n793_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n810_), .A2(new_n811_), .A3(G106gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n811_), .B1(new_n810_), .B2(G106gat), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n809_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT53), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n809_), .B(new_n816_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1339gat));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819_));
  OAI21_X1  g618(.A(KEYINPUT122), .B1(new_n298_), .B2(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n301_), .A2(KEYINPUT12), .ZN(new_n821_));
  NOR2_X1   g620(.A1(new_n349_), .A2(new_n350_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n297_), .ZN(new_n823_));
  AOI22_X1  g622(.A1(new_n276_), .A2(new_n821_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT122), .ZN(new_n825_));
  NAND4_X1  g624(.A1(new_n824_), .A2(new_n825_), .A3(KEYINPUT55), .A4(new_n282_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n279_), .B1(new_n294_), .B2(new_n297_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(new_n281_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n298_), .A2(new_n819_), .ZN(new_n829_));
  NAND4_X1  g628(.A1(new_n820_), .A2(new_n826_), .A3(new_n828_), .A4(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n310_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT56), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n830_), .A2(KEYINPUT56), .A3(new_n310_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n651_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n643_), .A2(new_n645_), .A3(new_n649_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n655_), .B1(new_n648_), .B2(new_n646_), .ZN(new_n838_));
  AOI22_X1  g637(.A1(new_n836_), .A2(new_n655_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  AND2_X1   g638(.A1(new_n839_), .A2(new_n312_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n835_), .A2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n835_), .A2(KEYINPUT58), .A3(new_n840_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n712_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846_));
  NAND4_X1  g645(.A1(new_n830_), .A2(KEYINPUT123), .A3(KEYINPUT56), .A4(new_n310_), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n847_), .A2(new_n312_), .A3(new_n656_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n833_), .A2(new_n849_), .A3(new_n834_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n848_), .A2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n313_), .A2(new_n839_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n846_), .B1(new_n853_), .B2(new_n670_), .ZN(new_n854_));
  AOI211_X1 g653(.A(KEYINPUT57), .B(new_n705_), .C1(new_n851_), .C2(new_n852_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n845_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n233_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n318_), .B(new_n754_), .C1(new_n377_), .C2(new_n378_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859_));
  OR3_X1    g658(.A1(new_n858_), .A2(new_n859_), .A3(KEYINPUT54), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n859_), .B1(new_n858_), .B2(KEYINPUT54), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(KEYINPUT54), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n857_), .A2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT59), .ZN(new_n865_));
  NAND3_X1  g664(.A1(new_n636_), .A2(new_n444_), .A3(new_n611_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n864_), .A2(new_n865_), .A3(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n856_), .A2(new_n674_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n866_), .B1(new_n869_), .B2(new_n863_), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n868_), .B1(new_n865_), .B2(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(G113gat), .B1(new_n871_), .B2(new_n761_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n870_), .ZN(new_n873_));
  OR3_X1    g672(.A1(new_n873_), .A2(G113gat), .A3(new_n761_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(G1340gat));
  OAI21_X1  g674(.A(G120gat), .B1(new_n871_), .B2(new_n318_), .ZN(new_n876_));
  INV_X1    g675(.A(G120gat), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n318_), .B2(KEYINPUT60), .ZN(new_n878_));
  OAI211_X1 g677(.A(new_n870_), .B(new_n878_), .C1(KEYINPUT60), .C2(new_n877_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n876_), .A2(new_n879_), .ZN(G1341gat));
  OAI21_X1  g679(.A(G127gat), .B1(new_n871_), .B2(new_n674_), .ZN(new_n881_));
  OR3_X1    g680(.A1(new_n873_), .A2(G127gat), .A3(new_n233_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n881_), .A2(new_n882_), .ZN(G1342gat));
  INV_X1    g682(.A(new_n712_), .ZN(new_n884_));
  OAI21_X1  g683(.A(G134gat), .B1(new_n871_), .B2(new_n884_), .ZN(new_n885_));
  OR3_X1    g684(.A1(new_n873_), .A2(G134gat), .A3(new_n670_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1343gat));
  NAND2_X1  g686(.A1(new_n869_), .A2(new_n863_), .ZN(new_n888_));
  NOR3_X1   g687(.A1(new_n589_), .A2(new_n444_), .A3(new_n637_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n890_), .A2(new_n761_), .ZN(new_n891_));
  XOR2_X1   g690(.A(KEYINPUT124), .B(G141gat), .Z(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1344gat));
  NAND3_X1  g692(.A1(new_n888_), .A2(new_n707_), .A3(new_n889_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g694(.A1(new_n890_), .A2(new_n233_), .ZN(new_n896_));
  XOR2_X1   g695(.A(KEYINPUT61), .B(G155gat), .Z(new_n897_));
  XNOR2_X1  g696(.A(new_n896_), .B(new_n897_), .ZN(G1346gat));
  OAI21_X1  g697(.A(G162gat), .B1(new_n890_), .B2(new_n884_), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n670_), .A2(G162gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n890_), .B2(new_n900_), .ZN(G1347gat));
  INV_X1    g700(.A(KEYINPUT22), .ZN(new_n902_));
  NOR3_X1   g701(.A1(new_n638_), .A2(new_n520_), .A3(new_n588_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n864_), .A2(new_n902_), .A3(new_n656_), .A4(new_n903_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n904_), .A2(KEYINPUT62), .A3(new_n405_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(KEYINPUT62), .ZN(new_n906_));
  AND3_X1   g705(.A1(new_n864_), .A2(new_n656_), .A3(new_n903_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT62), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n405_), .B1(new_n907_), .B2(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n905_), .B1(new_n906_), .B2(new_n909_), .ZN(G1348gat));
  NAND2_X1  g709(.A1(new_n864_), .A2(new_n903_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  AOI21_X1  g711(.A(G176gat), .B1(new_n912_), .B2(new_n707_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n888_), .A2(new_n903_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n318_), .A2(new_n406_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n913_), .B1(new_n914_), .B2(new_n915_), .ZN(G1349gat));
  AOI21_X1  g715(.A(G183gat), .B1(new_n914_), .B2(new_n234_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n911_), .A2(new_n674_), .A3(new_n400_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n911_), .B2(new_n884_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n705_), .A2(new_n536_), .A3(new_n540_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n911_), .B2(new_n921_), .ZN(G1351gat));
  NOR4_X1   g721(.A1(new_n750_), .A2(new_n444_), .A3(new_n611_), .A4(new_n588_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n888_), .A2(new_n923_), .ZN(new_n924_));
  NOR2_X1   g723(.A1(new_n924_), .A2(new_n761_), .ZN(new_n925_));
  XNOR2_X1  g724(.A(new_n925_), .B(new_n494_), .ZN(G1352gat));
  AND2_X1   g725(.A1(new_n888_), .A2(new_n923_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n927_), .A2(new_n707_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n491_), .A2(KEYINPUT125), .ZN(new_n929_));
  XNOR2_X1  g728(.A(new_n928_), .B(new_n929_), .ZN(G1353gat));
  INV_X1    g729(.A(KEYINPUT63), .ZN(new_n931_));
  INV_X1    g730(.A(G211gat), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n232_), .B1(new_n931_), .B2(new_n932_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(KEYINPUT126), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n927_), .A2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n931_), .A2(new_n932_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n935_), .B(new_n936_), .ZN(G1354gat));
  OR3_X1    g736(.A1(new_n924_), .A2(G218gat), .A3(new_n670_), .ZN(new_n938_));
  OAI21_X1  g737(.A(G218gat), .B1(new_n924_), .B2(new_n884_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1355gat));
endmodule


