//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:46 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n586_, new_n587_,
    new_n588_, new_n589_, new_n591_, new_n592_, new_n593_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n630_, new_n631_, new_n632_, new_n634_,
    new_n635_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n755_, new_n756_, new_n757_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n767_, new_n769_,
    new_n770_, new_n772_, new_n773_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n831_, new_n832_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT20), .ZN(new_n203_));
  NOR2_X1   g002(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(G169gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(KEYINPUT86), .B(G190gat), .Z(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(G183gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(G183gat), .A2(G190gat), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT23), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n208_), .B(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n205_), .B1(new_n207_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT24), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G169gat), .A2(G176gat), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n210_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G169gat), .ZN(new_n215_));
  INV_X1    g014(.A(G176gat), .ZN(new_n216_));
  OAI21_X1  g015(.A(KEYINPUT24), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n214_), .B1(new_n213_), .B2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(G183gat), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n219_), .A2(KEYINPUT85), .ZN(new_n220_));
  XOR2_X1   g019(.A(new_n220_), .B(KEYINPUT25), .Z(new_n221_));
  NOR2_X1   g020(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n222_), .B1(new_n206_), .B2(KEYINPUT26), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n221_), .A2(new_n223_), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n211_), .B1(new_n218_), .B2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT87), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n225_), .B(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(G204gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G197gat), .ZN(new_n229_));
  OR2_X1    g028(.A1(new_n229_), .A2(KEYINPUT93), .ZN(new_n230_));
  INV_X1    g029(.A(G197gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(G204gat), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n229_), .A2(KEYINPUT93), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n230_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G211gat), .B(G218gat), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT21), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n234_), .A2(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(new_n235_), .B1(new_n234_), .B2(KEYINPUT21), .ZN(new_n239_));
  AOI21_X1  g038(.A(new_n236_), .B1(new_n229_), .B2(new_n232_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT92), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n238_), .B1(new_n239_), .B2(new_n241_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n203_), .B1(new_n227_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G226gat), .A2(G233gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT19), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(G183gat), .A2(G190gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n205_), .B1(new_n210_), .B2(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT95), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n217_), .A2(new_n249_), .ZN(new_n250_));
  AOI21_X1  g049(.A(new_n213_), .B1(new_n217_), .B2(new_n249_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT26), .B(G190gat), .ZN(new_n252_));
  XNOR2_X1  g051(.A(KEYINPUT25), .B(G183gat), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n250_), .A2(new_n251_), .B1(new_n252_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT96), .ZN(new_n255_));
  AND2_X1   g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n214_), .B1(new_n254_), .B2(new_n255_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n248_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n243_), .B(new_n246_), .C1(new_n242_), .C2(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n242_), .ZN(new_n260_));
  OAI211_X1 g059(.A(KEYINPUT20), .B(new_n260_), .C1(new_n227_), .C2(new_n242_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(new_n245_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n259_), .A2(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G8gat), .B(G36gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT18), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G64gat), .B(G92gat), .ZN(new_n266_));
  XOR2_X1   g065(.A(new_n265_), .B(new_n266_), .Z(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n263_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT27), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n269_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n271_), .A2(KEYINPUT99), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT99), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n269_), .A2(new_n273_), .A3(new_n270_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n272_), .A2(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n242_), .B(KEYINPUT94), .ZN(new_n276_));
  OR2_X1    g075(.A1(new_n276_), .A2(new_n258_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n243_), .A2(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n245_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(new_n245_), .B2(new_n261_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n268_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n281_), .B(KEYINPUT27), .C1(new_n263_), .C2(new_n268_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n275_), .A2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G228gat), .A2(G233gat), .ZN(new_n284_));
  XOR2_X1   g083(.A(new_n284_), .B(KEYINPUT91), .Z(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G141gat), .A2(G148gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT89), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT2), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(G141gat), .ZN(new_n291_));
  INV_X1    g090(.A(G148gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  OR3_X1    g092(.A1(new_n293_), .A2(KEYINPUT90), .A3(KEYINPUT3), .ZN(new_n294_));
  NAND3_X1  g093(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n293_), .B1(KEYINPUT90), .B2(KEYINPUT3), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n290_), .A2(new_n294_), .A3(new_n295_), .A4(new_n296_), .ZN(new_n297_));
  XOR2_X1   g096(.A(G155gat), .B(G162gat), .Z(new_n298_));
  INV_X1    g097(.A(KEYINPUT1), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n301_));
  AND3_X1   g100(.A1(new_n288_), .A2(new_n293_), .A3(new_n301_), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n297_), .A2(new_n298_), .B1(new_n300_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT29), .ZN(new_n304_));
  OR2_X1    g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n286_), .B1(new_n305_), .B2(new_n242_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n305_), .A2(new_n286_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n306_), .B1(new_n276_), .B2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G22gat), .B(G50gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n303_), .A2(new_n304_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT28), .ZN(new_n312_));
  XOR2_X1   g111(.A(G78gat), .B(G106gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  OR2_X1    g113(.A1(new_n310_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n310_), .A2(new_n314_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G227gat), .A2(G233gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(G15gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n227_), .B(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT31), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G71gat), .B(G99gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n322_), .B(G43gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(KEYINPUT88), .B(KEYINPUT30), .ZN(new_n324_));
  XNOR2_X1  g123(.A(new_n323_), .B(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G127gat), .B(G134gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G113gat), .B(G120gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n325_), .B(new_n328_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n321_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n321_), .A2(new_n329_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(G225gat), .A2(G233gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n303_), .B(new_n328_), .Z(new_n334_));
  NAND2_X1  g133(.A1(new_n334_), .A2(KEYINPUT4), .ZN(new_n335_));
  OR3_X1    g134(.A1(new_n303_), .A2(KEYINPUT4), .A3(new_n328_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n333_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G1gat), .B(G29gat), .ZN(new_n338_));
  INV_X1    g137(.A(G85gat), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n338_), .B(new_n339_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(KEYINPUT0), .B(G57gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n333_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n334_), .A2(new_n343_), .ZN(new_n344_));
  OR3_X1    g143(.A1(new_n337_), .A2(new_n342_), .A3(new_n344_), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n342_), .B1(new_n337_), .B2(new_n344_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n332_), .A2(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n283_), .A2(new_n317_), .A3(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT100), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n283_), .A2(KEYINPUT100), .A3(new_n317_), .A4(new_n348_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n317_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n347_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n275_), .A2(new_n353_), .A3(new_n354_), .A4(new_n282_), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n267_), .A2(KEYINPUT32), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n280_), .A2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n357_), .B(new_n347_), .C1(new_n263_), .C2(new_n356_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n335_), .A2(new_n333_), .A3(new_n336_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n342_), .B1(new_n334_), .B2(new_n343_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT97), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363_));
  OR2_X1    g162(.A1(new_n346_), .A2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n346_), .A2(new_n363_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n362_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n358_), .B1(new_n366_), .B2(new_n269_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n367_), .A2(KEYINPUT98), .A3(new_n317_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n317_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT98), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n355_), .A2(new_n368_), .A3(new_n371_), .ZN(new_n372_));
  AOI22_X1  g171(.A1(new_n351_), .A2(new_n352_), .B1(new_n372_), .B2(new_n332_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT73), .ZN(new_n374_));
  NAND2_X1  g173(.A1(G99gat), .A2(G106gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT6), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT6), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n377_), .A2(G99gat), .A3(G106gat), .ZN(new_n378_));
  AND3_X1   g177(.A1(new_n376_), .A2(new_n378_), .A3(KEYINPUT70), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT70), .B1(new_n376_), .B2(new_n378_), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(G99gat), .ZN(new_n382_));
  INV_X1    g181(.A(G106gat), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT68), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT7), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT7), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT68), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n384_), .B1(new_n386_), .B2(new_n388_), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n382_), .A2(new_n383_), .B1(new_n387_), .B2(KEYINPUT68), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT71), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n384_), .A2(new_n388_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT71), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT68), .B(KEYINPUT7), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n392_), .B(new_n393_), .C1(new_n394_), .C2(new_n384_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n381_), .A2(new_n391_), .A3(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G92gat), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n339_), .A2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(G85gat), .A2(G92gat), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(KEYINPUT72), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n401_), .A2(KEYINPUT8), .ZN(new_n402_));
  AOI21_X1  g201(.A(KEYINPUT72), .B1(new_n396_), .B2(new_n400_), .ZN(new_n403_));
  OAI21_X1  g202(.A(new_n374_), .B1(new_n402_), .B2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n396_), .A2(new_n400_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT72), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  NAND4_X1  g206(.A1(new_n407_), .A2(KEYINPUT73), .A3(KEYINPUT8), .A4(new_n401_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT8), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n376_), .A2(new_n378_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT66), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n392_), .B1(new_n394_), .B2(new_n384_), .ZN(new_n412_));
  OAI211_X1 g211(.A(new_n409_), .B(new_n400_), .C1(new_n411_), .C2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT69), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n404_), .A2(new_n408_), .A3(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(KEYINPUT10), .B(G99gat), .Z(new_n416_));
  AOI21_X1  g215(.A(new_n411_), .B1(new_n383_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n398_), .ZN(new_n418_));
  INV_X1    g217(.A(KEYINPUT9), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n418_), .A2(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(KEYINPUT65), .ZN(new_n421_));
  INV_X1    g220(.A(new_n399_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n422_), .B1(new_n418_), .B2(new_n419_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n417_), .B1(new_n421_), .B2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT67), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n415_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(G29gat), .B(G36gat), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n429_), .B(KEYINPUT80), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G43gat), .B(G50gat), .ZN(new_n431_));
  XOR2_X1   g230(.A(new_n430_), .B(new_n431_), .Z(new_n432_));
  INV_X1    g231(.A(KEYINPUT35), .ZN(new_n433_));
  XNOR2_X1  g232(.A(KEYINPUT79), .B(KEYINPUT34), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G232gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n434_), .B(new_n435_), .ZN(new_n436_));
  AOI22_X1  g235(.A1(new_n428_), .A2(new_n432_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT81), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n432_), .B(KEYINPUT15), .ZN(new_n439_));
  AND3_X1   g238(.A1(new_n427_), .A2(new_n438_), .A3(new_n439_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n438_), .B1(new_n427_), .B2(new_n439_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n437_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n436_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n442_), .A2(KEYINPUT35), .A3(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(G190gat), .B(G218gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(G134gat), .B(G162gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n447_), .A2(KEYINPUT36), .ZN(new_n448_));
  OAI221_X1 g247(.A(new_n437_), .B1(new_n433_), .B2(new_n436_), .C1(new_n440_), .C2(new_n441_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n444_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  XOR2_X1   g249(.A(new_n447_), .B(KEYINPUT36), .Z(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n452_), .B1(new_n444_), .B2(new_n449_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT37), .B1(new_n450_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n444_), .A2(new_n449_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(new_n451_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT37), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n444_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n456_), .A2(new_n457_), .A3(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n454_), .A2(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(G127gat), .B(G155gat), .Z(new_n462_));
  XNOR2_X1  g261(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n463_));
  XNOR2_X1  g262(.A(new_n462_), .B(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G183gat), .B(G211gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n466_), .A2(KEYINPUT17), .ZN(new_n467_));
  XOR2_X1   g266(.A(G1gat), .B(G8gat), .Z(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT82), .ZN(new_n469_));
  INV_X1    g268(.A(G8gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n202_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(G15gat), .ZN(new_n473_));
  INV_X1    g272(.A(G22gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G15gat), .A2(G22gat), .ZN(new_n476_));
  AOI22_X1  g275(.A1(new_n472_), .A2(KEYINPUT14), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  OR2_X1    g276(.A1(new_n469_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n469_), .A2(new_n477_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n478_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(G231gat), .A2(G233gat), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n480_), .B(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G57gat), .B(G64gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT11), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n484_), .B(KEYINPUT74), .ZN(new_n485_));
  XOR2_X1   g284(.A(G71gat), .B(G78gat), .Z(new_n486_));
  OAI21_X1  g285(.A(new_n486_), .B1(KEYINPUT11), .B2(new_n483_), .ZN(new_n487_));
  OR2_X1    g286(.A1(new_n485_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n487_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(new_n482_), .B(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n467_), .B1(new_n491_), .B2(KEYINPUT75), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n492_), .B1(KEYINPUT75), .B2(new_n491_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n466_), .B(KEYINPUT17), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n494_), .B(KEYINPUT84), .Z(new_n495_));
  OR2_X1    g294(.A1(new_n495_), .A2(new_n491_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  NOR3_X1   g296(.A1(new_n373_), .A2(new_n461_), .A3(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT13), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G230gat), .A2(G233gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT64), .ZN(new_n501_));
  INV_X1    g300(.A(new_n501_), .ZN(new_n502_));
  AND3_X1   g301(.A1(new_n415_), .A2(new_n426_), .A3(new_n490_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n490_), .B1(new_n415_), .B2(new_n426_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n502_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G120gat), .B(G148gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n506_), .B(KEYINPUT5), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G176gat), .B(G204gat), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n507_), .B(new_n508_), .Z(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT75), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n490_), .A2(new_n511_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n488_), .A2(KEYINPUT75), .A3(new_n489_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(KEYINPUT12), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n427_), .A2(new_n515_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n516_), .B1(KEYINPUT12), .B2(new_n504_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n415_), .A2(new_n426_), .A3(new_n490_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n518_), .A2(new_n501_), .ZN(new_n519_));
  OAI211_X1 g318(.A(new_n505_), .B(new_n510_), .C1(new_n517_), .C2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT77), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n519_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n490_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n427_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT12), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n523_), .A2(new_n527_), .A3(new_n516_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n528_), .A2(KEYINPUT77), .A3(new_n505_), .A4(new_n510_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n522_), .A2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT12), .B1(new_n427_), .B2(new_n524_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n514_), .B1(new_n415_), .B2(new_n426_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n531_), .A2(new_n519_), .A3(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n505_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT76), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT76), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n536_), .B(new_n505_), .C1(new_n517_), .C2(new_n519_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n535_), .A2(new_n509_), .A3(new_n537_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n530_), .A2(new_n538_), .A3(KEYINPUT78), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT78), .B1(new_n530_), .B2(new_n538_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n499_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n530_), .A2(new_n538_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT78), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n530_), .A2(new_n538_), .A3(KEYINPUT78), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n544_), .A2(KEYINPUT13), .A3(new_n545_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n541_), .A2(new_n546_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n439_), .A2(new_n479_), .A3(new_n478_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n480_), .A2(new_n432_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(G229gat), .A2(G233gat), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n548_), .A2(new_n549_), .A3(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n480_), .B(new_n432_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n550_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n551_), .A2(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(G113gat), .B(G141gat), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G169gat), .B(G197gat), .ZN(new_n557_));
  XOR2_X1   g356(.A(new_n556_), .B(new_n557_), .Z(new_n558_));
  XNOR2_X1  g357(.A(new_n555_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n547_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AND4_X1   g361(.A1(new_n202_), .A2(new_n498_), .A3(new_n562_), .A4(new_n347_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n563_), .A2(KEYINPUT101), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(KEYINPUT101), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(new_n565_), .A3(KEYINPUT38), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT102), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT38), .B1(new_n564_), .B2(new_n565_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n456_), .A2(new_n458_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  NOR3_X1   g370(.A1(new_n373_), .A2(new_n571_), .A3(new_n497_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n562_), .ZN(new_n573_));
  OAI21_X1  g372(.A(G1gat), .B1(new_n573_), .B2(new_n354_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n574_), .B(KEYINPUT103), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n569_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n568_), .A2(new_n576_), .ZN(G1324gat));
  NOR2_X1   g376(.A1(new_n573_), .A2(new_n283_), .ZN(new_n578_));
  OR3_X1    g377(.A1(new_n578_), .A2(KEYINPUT39), .A3(new_n470_), .ZN(new_n579_));
  OAI21_X1  g378(.A(KEYINPUT39), .B1(new_n578_), .B2(new_n470_), .ZN(new_n580_));
  AND2_X1   g379(.A1(new_n498_), .A2(new_n562_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n283_), .A2(G8gat), .ZN(new_n582_));
  AOI22_X1  g381(.A1(new_n579_), .A2(new_n580_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n584_));
  XOR2_X1   g383(.A(new_n583_), .B(new_n584_), .Z(G1325gat));
  OAI21_X1  g384(.A(G15gat), .B1(new_n573_), .B2(new_n332_), .ZN(new_n586_));
  XOR2_X1   g385(.A(new_n586_), .B(KEYINPUT41), .Z(new_n587_));
  INV_X1    g386(.A(new_n332_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n581_), .A2(new_n473_), .A3(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n587_), .A2(new_n589_), .ZN(G1326gat));
  OAI21_X1  g389(.A(G22gat), .B1(new_n573_), .B2(new_n317_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT42), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n581_), .A2(new_n474_), .A3(new_n353_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(G1327gat));
  NOR2_X1   g393(.A1(new_n373_), .A2(new_n570_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n497_), .ZN(new_n596_));
  NOR2_X1   g395(.A1(new_n561_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n598_), .B(KEYINPUT106), .ZN(new_n599_));
  AOI21_X1  g398(.A(G29gat), .B1(new_n599_), .B2(new_n347_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n373_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n601_), .A2(new_n461_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(new_n602_), .ZN(new_n604_));
  NOR2_X1   g403(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n605_));
  OAI22_X1  g404(.A1(new_n373_), .A2(new_n460_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n603_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(new_n597_), .ZN(new_n608_));
  INV_X1    g407(.A(KEYINPUT44), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n608_), .A2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n607_), .A2(KEYINPUT44), .A3(new_n597_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n347_), .A2(G29gat), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n600_), .B1(new_n613_), .B2(new_n614_), .ZN(G1328gat));
  OAI21_X1  g414(.A(G36gat), .B1(new_n612_), .B2(new_n283_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n598_), .B(KEYINPUT106), .Z(new_n618_));
  INV_X1    g417(.A(new_n283_), .ZN(new_n619_));
  INV_X1    g418(.A(G36gat), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n617_), .B1(new_n618_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n617_), .ZN(new_n623_));
  NAND4_X1  g422(.A1(new_n599_), .A2(new_n620_), .A3(new_n619_), .A4(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n616_), .A2(new_n622_), .A3(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT46), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n616_), .A2(new_n622_), .A3(new_n624_), .A4(KEYINPUT46), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(new_n628_), .ZN(G1329gat));
  NOR2_X1   g428(.A1(new_n618_), .A2(new_n332_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n588_), .A2(G43gat), .ZN(new_n631_));
  OAI22_X1  g430(.A1(new_n630_), .A2(G43gat), .B1(new_n612_), .B2(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g432(.A(G50gat), .B1(new_n599_), .B2(new_n353_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n353_), .A2(G50gat), .ZN(new_n635_));
  AOI21_X1  g434(.A(new_n634_), .B1(new_n613_), .B2(new_n635_), .ZN(G1331gat));
  NOR2_X1   g435(.A1(new_n547_), .A2(new_n560_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n572_), .A2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT108), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  OAI21_X1  g439(.A(G57gat), .B1(new_n640_), .B2(new_n354_), .ZN(new_n641_));
  AND2_X1   g440(.A1(new_n498_), .A2(new_n637_), .ZN(new_n642_));
  INV_X1    g441(.A(G57gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n642_), .A2(new_n643_), .A3(new_n347_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n644_), .ZN(G1332gat));
  INV_X1    g444(.A(G64gat), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n642_), .A2(new_n646_), .A3(new_n619_), .ZN(new_n647_));
  OAI21_X1  g446(.A(G64gat), .B1(new_n640_), .B2(new_n283_), .ZN(new_n648_));
  AND2_X1   g447(.A1(new_n648_), .A2(KEYINPUT48), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n648_), .A2(KEYINPUT48), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n647_), .B1(new_n649_), .B2(new_n650_), .ZN(G1333gat));
  INV_X1    g450(.A(G71gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n642_), .A2(new_n652_), .A3(new_n588_), .ZN(new_n653_));
  OAI21_X1  g452(.A(G71gat), .B1(new_n640_), .B2(new_n332_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n654_), .A2(KEYINPUT49), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(KEYINPUT49), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n655_), .B2(new_n656_), .ZN(G1334gat));
  INV_X1    g456(.A(G78gat), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n642_), .A2(new_n658_), .A3(new_n353_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G78gat), .B1(new_n640_), .B2(new_n317_), .ZN(new_n660_));
  XOR2_X1   g459(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n660_), .A2(new_n662_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n659_), .B1(new_n663_), .B2(new_n664_), .ZN(G1335gat));
  NAND2_X1  g464(.A1(new_n637_), .A2(new_n497_), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n373_), .A2(new_n666_), .A3(new_n570_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT110), .Z(new_n668_));
  AOI21_X1  g467(.A(G85gat), .B1(new_n668_), .B2(new_n347_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n666_), .B(KEYINPUT111), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n607_), .A2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT112), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n354_), .A2(new_n339_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n669_), .B1(new_n672_), .B2(new_n673_), .ZN(G1336gat));
  AOI21_X1  g473(.A(G92gat), .B1(new_n668_), .B2(new_n619_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n283_), .A2(new_n397_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n672_), .B2(new_n676_), .ZN(G1337gat));
  NAND3_X1  g476(.A1(new_n668_), .A2(new_n416_), .A3(new_n588_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n671_), .A2(new_n332_), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n678_), .B1(new_n679_), .B2(new_n382_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g480(.A1(new_n668_), .A2(new_n383_), .A3(new_n353_), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n607_), .A2(new_n670_), .A3(new_n353_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(G106gat), .ZN(new_n684_));
  AND2_X1   g483(.A1(new_n684_), .A2(KEYINPUT52), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(KEYINPUT52), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n687_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g487(.A1(new_n560_), .A2(new_n497_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n541_), .A2(new_n546_), .A3(new_n460_), .A4(new_n689_), .ZN(new_n690_));
  OR2_X1    g489(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(KEYINPUT113), .A2(KEYINPUT54), .ZN(new_n693_));
  XOR2_X1   g492(.A(new_n693_), .B(KEYINPUT114), .Z(new_n694_));
  INV_X1    g493(.A(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n690_), .A2(new_n691_), .A3(new_n694_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n559_), .B1(new_n522_), .B2(new_n529_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT115), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n700_), .B1(new_n517_), .B2(new_n519_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n701_), .A2(KEYINPUT55), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT55), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n528_), .A2(new_n700_), .A3(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n502_), .B1(new_n517_), .B2(new_n503_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n702_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  AND3_X1   g505(.A1(new_n706_), .A2(KEYINPUT56), .A3(new_n509_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT56), .B1(new_n706_), .B2(new_n509_), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT116), .B(new_n699_), .C1(new_n707_), .C2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n555_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n548_), .A2(new_n549_), .A3(new_n553_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n558_), .B1(new_n552_), .B2(new_n550_), .ZN(new_n712_));
  AOI22_X1  g511(.A1(new_n710_), .A2(new_n558_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n713_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n709_), .A2(new_n714_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n532_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n716_));
  AOI21_X1  g515(.A(KEYINPUT115), .B1(new_n716_), .B2(new_n523_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n705_), .B1(new_n717_), .B2(new_n703_), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n701_), .A2(KEYINPUT55), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n509_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT56), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n706_), .A2(KEYINPUT56), .A3(new_n509_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(KEYINPUT116), .B1(new_n724_), .B2(new_n699_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n570_), .B1(new_n715_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT57), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT57), .B(new_n570_), .C1(new_n715_), .C2(new_n725_), .ZN(new_n729_));
  AND2_X1   g528(.A1(new_n530_), .A2(new_n713_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n724_), .A2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT58), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n460_), .B1(new_n731_), .B2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n724_), .A2(KEYINPUT58), .A3(new_n730_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n728_), .A2(new_n729_), .A3(new_n735_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n698_), .B1(new_n736_), .B2(new_n497_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  NOR4_X1   g537(.A1(new_n619_), .A2(new_n332_), .A3(new_n353_), .A4(new_n354_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  INV_X1    g540(.A(G113gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(new_n560_), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT117), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT59), .B1(new_n738_), .B2(new_n744_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(new_n745_), .B(new_n740_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(new_n560_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n747_), .B2(new_n742_), .ZN(G1340gat));
  INV_X1    g547(.A(G120gat), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n749_), .B1(new_n547_), .B2(KEYINPUT60), .ZN(new_n750_));
  OAI211_X1 g549(.A(new_n741_), .B(new_n750_), .C1(KEYINPUT60), .C2(new_n749_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n547_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n746_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n751_), .B1(new_n753_), .B2(new_n749_), .ZN(G1341gat));
  AND2_X1   g553(.A1(new_n746_), .A2(new_n596_), .ZN(new_n755_));
  INV_X1    g554(.A(G127gat), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n596_), .A2(new_n756_), .ZN(new_n757_));
  OAI22_X1  g556(.A1(new_n755_), .A2(new_n756_), .B1(new_n740_), .B2(new_n757_), .ZN(G1342gat));
  INV_X1    g557(.A(G134gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n741_), .A2(new_n759_), .A3(new_n571_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n746_), .A2(new_n461_), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n760_), .B1(new_n761_), .B2(new_n759_), .ZN(G1343gat));
  NOR2_X1   g561(.A1(new_n737_), .A2(new_n588_), .ZN(new_n763_));
  NAND4_X1  g562(.A1(new_n763_), .A2(new_n353_), .A3(new_n347_), .A4(new_n283_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n764_), .A2(new_n559_), .ZN(new_n765_));
  XNOR2_X1  g564(.A(new_n765_), .B(new_n291_), .ZN(G1344gat));
  NOR2_X1   g565(.A1(new_n764_), .A2(new_n547_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(new_n292_), .ZN(G1345gat));
  NOR2_X1   g567(.A1(new_n764_), .A2(new_n497_), .ZN(new_n769_));
  XOR2_X1   g568(.A(KEYINPUT61), .B(G155gat), .Z(new_n770_));
  XNOR2_X1  g569(.A(new_n769_), .B(new_n770_), .ZN(G1346gat));
  OAI21_X1  g570(.A(G162gat), .B1(new_n764_), .B2(new_n460_), .ZN(new_n772_));
  OR2_X1    g571(.A1(new_n570_), .A2(G162gat), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n772_), .B1(new_n764_), .B2(new_n773_), .ZN(G1347gat));
  NAND3_X1  g573(.A1(new_n619_), .A2(new_n317_), .A3(new_n348_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n737_), .A2(new_n775_), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  NOR3_X1   g576(.A1(new_n777_), .A2(KEYINPUT118), .A3(new_n559_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n778_), .A2(new_n215_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT62), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT118), .B1(new_n777_), .B2(new_n559_), .ZN(new_n781_));
  AND3_X1   g580(.A1(new_n779_), .A2(new_n780_), .A3(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n780_), .B1(new_n779_), .B2(new_n781_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT119), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n737_), .B2(new_n775_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n775_), .ZN(new_n786_));
  AOI22_X1  g585(.A1(new_n726_), .A2(new_n727_), .B1(new_n734_), .B2(new_n733_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n596_), .B1(new_n787_), .B2(new_n729_), .ZN(new_n788_));
  OAI211_X1 g587(.A(KEYINPUT119), .B(new_n786_), .C1(new_n788_), .C2(new_n698_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  XNOR2_X1  g590(.A(KEYINPUT22), .B(G169gat), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n560_), .A2(new_n792_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT120), .ZN(new_n794_));
  OAI22_X1  g593(.A1(new_n782_), .A2(new_n783_), .B1(new_n791_), .B2(new_n794_), .ZN(G1348gat));
  NAND3_X1  g594(.A1(new_n776_), .A2(G176gat), .A3(new_n752_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n790_), .A2(new_n752_), .ZN(new_n797_));
  AOI21_X1  g596(.A(KEYINPUT121), .B1(new_n797_), .B2(new_n216_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n547_), .B1(new_n785_), .B2(new_n789_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT121), .ZN(new_n800_));
  NOR3_X1   g599(.A1(new_n799_), .A2(new_n800_), .A3(G176gat), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n796_), .B1(new_n798_), .B2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT122), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT122), .ZN(new_n804_));
  OAI211_X1 g603(.A(new_n804_), .B(new_n796_), .C1(new_n798_), .C2(new_n801_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n803_), .A2(new_n805_), .ZN(G1349gat));
  NOR2_X1   g605(.A1(new_n777_), .A2(new_n497_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n497_), .A2(new_n253_), .ZN(new_n808_));
  OAI22_X1  g607(.A1(new_n807_), .A2(G183gat), .B1(new_n791_), .B2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT123), .ZN(G1350gat));
  NAND3_X1  g609(.A1(new_n790_), .A2(new_n252_), .A3(new_n571_), .ZN(new_n811_));
  INV_X1    g610(.A(G190gat), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n790_), .B2(new_n461_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n813_), .A2(KEYINPUT124), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(KEYINPUT124), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n811_), .B1(new_n814_), .B2(new_n815_), .ZN(G1351gat));
  NAND4_X1  g615(.A1(new_n763_), .A2(new_n353_), .A3(new_n354_), .A4(new_n619_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(new_n559_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(KEYINPUT125), .B(G197gat), .ZN(new_n819_));
  XNOR2_X1  g618(.A(new_n818_), .B(new_n819_), .ZN(G1352gat));
  NOR2_X1   g619(.A1(new_n817_), .A2(new_n547_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(new_n228_), .ZN(G1353gat));
  INV_X1    g621(.A(KEYINPUT126), .ZN(new_n823_));
  NOR2_X1   g622(.A1(new_n817_), .A2(new_n497_), .ZN(new_n824_));
  XOR2_X1   g623(.A(KEYINPUT63), .B(G211gat), .Z(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n827_), .B1(new_n817_), .B2(new_n497_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n823_), .B1(new_n826_), .B2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(new_n823_), .B2(new_n826_), .ZN(G1354gat));
  OAI21_X1  g629(.A(G218gat), .B1(new_n817_), .B2(new_n460_), .ZN(new_n831_));
  OR2_X1    g630(.A1(new_n570_), .A2(G218gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n817_), .B2(new_n832_), .ZN(G1355gat));
endmodule


