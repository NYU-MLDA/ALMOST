//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n896_, new_n897_, new_n898_, new_n899_,
    new_n901_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n943_, new_n944_, new_n945_, new_n946_, new_n948_,
    new_n949_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n959_, new_n960_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_;
  XOR2_X1   g000(.A(KEYINPUT10), .B(G99gat), .Z(new_n202_));
  INV_X1    g001(.A(G106gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G85gat), .B(G92gat), .Z(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT9), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT6), .ZN(new_n208_));
  INV_X1    g007(.A(G85gat), .ZN(new_n209_));
  INV_X1    g008(.A(G92gat), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n209_), .A2(new_n210_), .A3(KEYINPUT9), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n204_), .A2(new_n206_), .A3(new_n208_), .A4(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G57gat), .B(G64gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT11), .ZN(new_n214_));
  XOR2_X1   g013(.A(G71gat), .B(G78gat), .Z(new_n215_));
  OR2_X1    g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n213_), .A2(KEYINPUT11), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n214_), .A2(new_n215_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n216_), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT8), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT6), .ZN(new_n221_));
  XNOR2_X1  g020(.A(new_n207_), .B(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n208_), .A2(KEYINPUT65), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G99gat), .A2(G106gat), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT7), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n225_), .A3(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n220_), .B1(new_n228_), .B2(new_n205_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n226_), .B(new_n230_), .ZN(new_n231_));
  NOR2_X1   g030(.A1(new_n231_), .A2(new_n222_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n220_), .A2(KEYINPUT64), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n220_), .A2(KEYINPUT64), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n205_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  OAI211_X1 g035(.A(new_n212_), .B(new_n219_), .C1(new_n229_), .C2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n212_), .B1(new_n229_), .B2(new_n236_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n219_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n243_), .A2(G230gat), .A3(G233gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G230gat), .A2(G233gat), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n237_), .A2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n219_), .B(new_n247_), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(KEYINPUT12), .A3(new_n240_), .ZN(new_n249_));
  INV_X1    g048(.A(KEYINPUT12), .ZN(new_n250_));
  AOI21_X1  g049(.A(KEYINPUT68), .B1(new_n242_), .B2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n252_));
  AOI211_X1 g051(.A(new_n252_), .B(KEYINPUT12), .C1(new_n240_), .C2(new_n241_), .ZN(new_n253_));
  OAI211_X1 g052(.A(new_n246_), .B(new_n249_), .C1(new_n251_), .C2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n244_), .A2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(G120gat), .B(G148gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT5), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G176gat), .B(G204gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n257_), .B(new_n258_), .Z(new_n259_));
  NAND2_X1  g058(.A1(new_n255_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n259_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n244_), .A2(new_n254_), .A3(new_n261_), .ZN(new_n262_));
  AND2_X1   g061(.A1(new_n260_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(KEYINPUT13), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(new_n262_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT13), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n264_), .A2(new_n267_), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT69), .ZN(new_n269_));
  XOR2_X1   g068(.A(G29gat), .B(G36gat), .Z(new_n270_));
  XOR2_X1   g069(.A(G43gat), .B(G50gat), .Z(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT15), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n240_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n274_), .A2(KEYINPUT70), .ZN(new_n275_));
  NAND2_X1  g074(.A1(G232gat), .A2(G233gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT34), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n275_), .A2(KEYINPUT35), .A3(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n278_), .B1(KEYINPUT35), .B2(new_n277_), .ZN(new_n279_));
  INV_X1    g078(.A(new_n205_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n231_), .B1(KEYINPUT65), .B2(new_n208_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n280_), .B1(new_n281_), .B2(new_n224_), .ZN(new_n282_));
  OAI22_X1  g081(.A1(new_n282_), .A2(new_n220_), .B1(new_n232_), .B2(new_n235_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(new_n272_), .A3(new_n212_), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n279_), .A2(new_n274_), .A3(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n274_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G190gat), .B(G218gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G134gat), .B(G162gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  AOI22_X1  g088(.A1(new_n278_), .A2(new_n286_), .B1(KEYINPUT36), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n285_), .A2(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n289_), .A2(KEYINPUT36), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  OAI211_X1 g092(.A(new_n285_), .B(new_n290_), .C1(KEYINPUT36), .C2(new_n289_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT37), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT37), .B1(new_n293_), .B2(new_n294_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  XOR2_X1   g098(.A(G127gat), .B(G155gat), .Z(new_n300_));
  XNOR2_X1  g099(.A(KEYINPUT74), .B(KEYINPUT16), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n300_), .B(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G183gat), .B(G211gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT17), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G1gat), .B(G8gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(KEYINPUT71), .B(G1gat), .ZN(new_n308_));
  INV_X1    g107(.A(G8gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT14), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT72), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G15gat), .B(G22gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n311_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n315_));
  OAI21_X1  g114(.A(new_n307_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n310_), .A2(new_n312_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT72), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n318_), .A2(new_n313_), .A3(new_n306_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n316_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT73), .ZN(new_n321_));
  AND2_X1   g120(.A1(G231gat), .A2(G233gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI21_X1  g123(.A(new_n305_), .B1(new_n324_), .B2(new_n219_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n325_), .B1(new_n219_), .B2(new_n324_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n304_), .A2(KEYINPUT17), .ZN(new_n327_));
  INV_X1    g126(.A(new_n248_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n327_), .B1(new_n323_), .B2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n329_), .B1(new_n328_), .B2(new_n323_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n326_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n299_), .A2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n269_), .A2(new_n333_), .ZN(new_n334_));
  XNOR2_X1  g133(.A(new_n334_), .B(KEYINPUT75), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT90), .ZN(new_n336_));
  XNOR2_X1  g135(.A(G22gat), .B(G50gat), .ZN(new_n337_));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n338_));
  INV_X1    g137(.A(G141gat), .ZN(new_n339_));
  INV_X1    g138(.A(G148gat), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n338_), .A2(new_n339_), .A3(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G141gat), .A2(G148gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT2), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n341_), .A2(new_n344_), .A3(new_n345_), .A4(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT85), .ZN(new_n348_));
  AND2_X1   g147(.A1(G155gat), .A2(G162gat), .ZN(new_n349_));
  NOR2_X1   g148(.A1(G155gat), .A2(G162gat), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n348_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(G155gat), .ZN(new_n352_));
  INV_X1    g151(.A(G162gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G155gat), .A2(G162gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(KEYINPUT85), .A3(new_n355_), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n347_), .A2(new_n351_), .A3(new_n356_), .ZN(new_n357_));
  XOR2_X1   g156(.A(G141gat), .B(G148gat), .Z(new_n358_));
  NAND2_X1  g157(.A1(new_n355_), .A2(KEYINPUT1), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(new_n354_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n355_), .A2(KEYINPUT1), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n358_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  AND2_X1   g161(.A1(new_n357_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT28), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n363_), .A2(new_n364_), .A3(new_n365_), .ZN(new_n366_));
  AND4_X1   g165(.A1(new_n344_), .A2(new_n341_), .A3(new_n345_), .A4(new_n346_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n351_), .A2(new_n356_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n362_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT28), .B1(new_n369_), .B2(KEYINPUT29), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n337_), .B1(new_n366_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n366_), .A2(new_n370_), .A3(new_n337_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT87), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n375_), .B1(new_n369_), .B2(KEYINPUT29), .ZN(new_n376_));
  INV_X1    g175(.A(G218gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(G211gat), .ZN(new_n378_));
  INV_X1    g177(.A(G211gat), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(G218gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(G197gat), .A2(G204gat), .ZN(new_n382_));
  NOR2_X1   g181(.A1(G197gat), .A2(G204gat), .ZN(new_n383_));
  NOR2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n381_), .B1(KEYINPUT21), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT89), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G197gat), .B(G204gat), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT21), .ZN(new_n388_));
  AOI21_X1  g187(.A(KEYINPUT88), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  OAI211_X1 g188(.A(KEYINPUT88), .B(new_n388_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  OAI211_X1 g190(.A(new_n385_), .B(new_n386_), .C1(new_n389_), .C2(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n381_), .A2(new_n384_), .A3(KEYINPUT21), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n395_), .B1(new_n384_), .B2(KEYINPUT21), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(new_n390_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n386_), .B1(new_n397_), .B2(new_n385_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n376_), .B1(new_n394_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT86), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G228gat), .A2(G233gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n385_), .B1(new_n389_), .B2(new_n391_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n403_), .A2(KEYINPUT89), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(new_n393_), .A3(new_n392_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT86), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n405_), .A2(new_n406_), .A3(new_n376_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n400_), .A2(new_n402_), .A3(new_n407_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n402_), .B1(new_n400_), .B2(new_n407_), .ZN(new_n409_));
  OAI211_X1 g208(.A(new_n336_), .B(new_n374_), .C1(new_n408_), .C2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n407_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n406_), .B1(new_n405_), .B2(new_n376_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n401_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n373_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n336_), .B1(new_n414_), .B2(new_n371_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n400_), .A2(new_n402_), .A3(new_n407_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n372_), .A2(KEYINPUT90), .A3(new_n373_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n413_), .A2(new_n415_), .A3(new_n416_), .A4(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n410_), .A2(new_n418_), .ZN(new_n419_));
  XOR2_X1   g218(.A(G78gat), .B(G106gat), .Z(new_n420_));
  INV_X1    g219(.A(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n410_), .A2(new_n418_), .A3(new_n420_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(G134gat), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(G127gat), .ZN(new_n426_));
  INV_X1    g225(.A(G127gat), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(G134gat), .ZN(new_n428_));
  AOI21_X1  g227(.A(KEYINPUT82), .B1(new_n426_), .B2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n426_), .A2(new_n428_), .A3(KEYINPUT82), .ZN(new_n431_));
  XNOR2_X1  g230(.A(G113gat), .B(G120gat), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n432_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n431_), .ZN(new_n435_));
  OAI21_X1  g234(.A(new_n434_), .B1(new_n435_), .B2(new_n429_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n433_), .A2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n363_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT93), .ZN(new_n439_));
  NAND4_X1  g238(.A1(new_n369_), .A2(new_n439_), .A3(new_n433_), .A4(new_n436_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(new_n440_), .A3(KEYINPUT4), .ZN(new_n441_));
  INV_X1    g240(.A(new_n437_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT4), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n442_), .A2(new_n439_), .A3(new_n443_), .A4(new_n369_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G225gat), .A2(G233gat), .ZN(new_n446_));
  INV_X1    g245(.A(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n449_), .B(G85gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(KEYINPUT0), .B(G57gat), .ZN(new_n451_));
  XOR2_X1   g250(.A(new_n450_), .B(new_n451_), .Z(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n442_), .A2(new_n369_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n447_), .B1(new_n454_), .B2(new_n438_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n448_), .A2(new_n453_), .A3(new_n456_), .ZN(new_n457_));
  AOI21_X1  g256(.A(new_n446_), .B1(new_n441_), .B2(new_n444_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n452_), .B1(new_n458_), .B2(new_n455_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G183gat), .A2(G190gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT23), .ZN(new_n462_));
  OR2_X1    g261(.A1(G183gat), .A2(G190gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT81), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT79), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT22), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n466_), .B1(new_n467_), .B2(G169gat), .ZN(new_n468_));
  AOI21_X1  g267(.A(G176gat), .B1(new_n467_), .B2(G169gat), .ZN(new_n469_));
  INV_X1    g268(.A(G169gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n470_), .A2(KEYINPUT79), .A3(KEYINPUT22), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n468_), .A2(new_n469_), .A3(KEYINPUT80), .A4(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G169gat), .A2(G176gat), .ZN(new_n473_));
  AND2_X1   g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n468_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT80), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n465_), .B1(new_n474_), .B2(new_n477_), .ZN(new_n478_));
  AND4_X1   g277(.A1(new_n465_), .A2(new_n477_), .A3(new_n473_), .A4(new_n472_), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n464_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NOR2_X1   g279(.A1(new_n394_), .A2(new_n398_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n473_), .A2(KEYINPUT24), .ZN(new_n482_));
  NOR2_X1   g281(.A1(G169gat), .A2(G176gat), .ZN(new_n483_));
  MUX2_X1   g282(.A(new_n482_), .B(KEYINPUT24), .S(new_n483_), .Z(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT25), .B(G183gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT78), .ZN(new_n486_));
  INV_X1    g285(.A(G190gat), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT26), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  OR2_X1    g287(.A1(new_n487_), .A2(KEYINPUT26), .ZN(new_n489_));
  OAI211_X1 g288(.A(new_n485_), .B(new_n488_), .C1(new_n489_), .C2(new_n486_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n484_), .A2(new_n462_), .A3(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n480_), .A2(new_n481_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G226gat), .A2(G233gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT19), .ZN(new_n494_));
  INV_X1    g293(.A(new_n494_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT20), .ZN(new_n496_));
  XNOR2_X1  g295(.A(KEYINPUT26), .B(G190gat), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n485_), .A2(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n498_), .A2(new_n462_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(new_n484_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n470_), .A2(KEYINPUT22), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n467_), .A2(G169gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n503_), .A2(KEYINPUT91), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n503_), .A2(KEYINPUT91), .ZN(new_n506_));
  AOI21_X1  g305(.A(G176gat), .B1(new_n505_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n464_), .A2(new_n473_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n500_), .B1(new_n507_), .B2(new_n508_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n496_), .B1(new_n405_), .B2(new_n509_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n492_), .A2(new_n495_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n508_), .ZN(new_n512_));
  INV_X1    g311(.A(G176gat), .ZN(new_n513_));
  INV_X1    g312(.A(new_n506_), .ZN(new_n514_));
  OAI21_X1  g313(.A(new_n513_), .B1(new_n514_), .B2(new_n504_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n512_), .A2(new_n515_), .B1(new_n484_), .B2(new_n499_), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n496_), .B1(new_n481_), .B2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n464_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n477_), .A2(new_n473_), .A3(new_n472_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT81), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n474_), .A2(new_n465_), .A3(new_n477_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n518_), .B1(new_n520_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n491_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n405_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n495_), .B1(new_n517_), .B2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n511_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G8gat), .B(G36gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n527_), .B(KEYINPUT18), .ZN(new_n528_));
  XNOR2_X1  g327(.A(G64gat), .B(G92gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n528_), .B(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(KEYINPUT32), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n460_), .B1(new_n526_), .B2(new_n532_), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n522_), .A2(new_n405_), .A3(new_n523_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT20), .B1(new_n481_), .B2(new_n516_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n494_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n517_), .A2(new_n524_), .A3(new_n495_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n532_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT96), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT96), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n536_), .A2(new_n540_), .A3(new_n537_), .A4(new_n532_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n533_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n424_), .A2(new_n542_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n517_), .A2(new_n524_), .A3(new_n495_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n495_), .B1(new_n492_), .B2(new_n510_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n544_), .A2(new_n545_), .A3(new_n530_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n531_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n547_));
  OR3_X1    g346(.A1(new_n546_), .A2(new_n547_), .A3(KEYINPUT92), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n454_), .A2(new_n438_), .A3(new_n447_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n453_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT95), .ZN(new_n551_));
  OAI22_X1  g350(.A1(new_n550_), .A2(new_n551_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n552_));
  AOI21_X1  g351(.A(new_n552_), .B1(new_n551_), .B2(new_n550_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n459_), .A2(KEYINPUT94), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT33), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n459_), .A2(KEYINPUT94), .A3(KEYINPUT33), .ZN(new_n557_));
  AOI21_X1  g356(.A(new_n553_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  OAI21_X1  g357(.A(KEYINPUT92), .B1(new_n546_), .B2(new_n547_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n548_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n543_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(KEYINPUT27), .ZN(new_n562_));
  OAI21_X1  g361(.A(new_n562_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n530_), .B1(new_n511_), .B2(new_n525_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n536_), .A2(new_n531_), .A3(new_n537_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n564_), .A2(KEYINPUT27), .A3(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT97), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n460_), .A2(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n457_), .A2(KEYINPUT97), .A3(new_n459_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n424_), .B1(new_n567_), .B2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n437_), .B(KEYINPUT31), .ZN(new_n573_));
  XNOR2_X1  g372(.A(G71gat), .B(G99gat), .ZN(new_n574_));
  INV_X1    g373(.A(G43gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n574_), .B(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n576_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n576_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n480_), .A2(new_n491_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(G227gat), .A2(G233gat), .ZN(new_n580_));
  INV_X1    g379(.A(G15gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n582_), .B(KEYINPUT30), .ZN(new_n583_));
  AND3_X1   g382(.A1(new_n577_), .A2(new_n579_), .A3(new_n583_), .ZN(new_n584_));
  AOI21_X1  g383(.A(new_n583_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n585_));
  OAI21_X1  g384(.A(new_n573_), .B1(new_n584_), .B2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT83), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT83), .B(new_n573_), .C1(new_n584_), .C2(new_n585_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n577_), .A2(new_n579_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n583_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n573_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n577_), .A2(new_n579_), .A3(new_n583_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(KEYINPUT84), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n593_), .A2(KEYINPUT84), .A3(new_n594_), .A4(new_n595_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n590_), .A2(new_n600_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n561_), .A2(new_n572_), .A3(new_n602_), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n422_), .A2(new_n423_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n571_), .B1(new_n590_), .B2(new_n600_), .ZN(new_n605_));
  AND3_X1   g404(.A1(new_n564_), .A2(KEYINPUT27), .A3(new_n565_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n530_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n607_));
  AOI21_X1  g406(.A(KEYINPUT27), .B1(new_n607_), .B2(new_n565_), .ZN(new_n608_));
  NOR3_X1   g407(.A1(new_n606_), .A2(new_n608_), .A3(KEYINPUT98), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT98), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n610_), .B1(new_n563_), .B2(new_n566_), .ZN(new_n611_));
  OAI211_X1 g410(.A(new_n604_), .B(new_n605_), .C1(new_n609_), .C2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(KEYINPUT99), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT99), .ZN(new_n614_));
  OAI21_X1  g413(.A(KEYINPUT98), .B1(new_n606_), .B2(new_n608_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n563_), .A2(new_n610_), .A3(new_n566_), .ZN(new_n616_));
  AOI21_X1  g415(.A(new_n424_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(new_n614_), .B1(new_n617_), .B2(new_n605_), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n603_), .B1(new_n613_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT76), .ZN(new_n620_));
  INV_X1    g419(.A(new_n272_), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n316_), .A2(new_n621_), .A3(new_n319_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n621_), .B1(new_n316_), .B2(new_n319_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n620_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n624_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n626_), .A2(KEYINPUT76), .A3(new_n622_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(G229gat), .A2(G233gat), .ZN(new_n628_));
  INV_X1    g427(.A(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n625_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT15), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n272_), .B(new_n631_), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n626_), .B(new_n628_), .C1(new_n632_), .C2(new_n320_), .ZN(new_n633_));
  XNOR2_X1  g432(.A(G113gat), .B(G141gat), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G169gat), .B(G197gat), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n634_), .B(new_n635_), .Z(new_n636_));
  NAND3_X1  g435(.A1(new_n630_), .A2(new_n633_), .A3(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n636_), .B1(new_n630_), .B2(new_n633_), .ZN(new_n639_));
  OAI21_X1  g438(.A(KEYINPUT77), .B1(new_n638_), .B2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n639_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT77), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n641_), .A2(new_n642_), .A3(new_n637_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  AND3_X1   g443(.A1(new_n335_), .A2(new_n619_), .A3(new_n644_), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n645_), .A2(new_n571_), .A3(new_n308_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT38), .ZN(new_n647_));
  INV_X1    g446(.A(new_n644_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n268_), .A2(new_n648_), .A3(new_n331_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT100), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n612_), .A2(KEYINPUT99), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n617_), .A2(new_n614_), .A3(new_n605_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n601_), .B1(new_n543_), .B2(new_n560_), .ZN(new_n653_));
  AOI22_X1  g452(.A1(new_n651_), .A2(new_n652_), .B1(new_n653_), .B2(new_n572_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n295_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n650_), .A2(new_n656_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT101), .ZN(new_n658_));
  INV_X1    g457(.A(new_n571_), .ZN(new_n659_));
  OAI21_X1  g458(.A(G1gat), .B1(new_n658_), .B2(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n647_), .A2(new_n660_), .ZN(G1324gat));
  NAND2_X1  g460(.A1(new_n615_), .A2(new_n616_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n645_), .A2(new_n309_), .A3(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(G8gat), .B1(new_n657_), .B2(new_n662_), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n665_), .B(KEYINPUT39), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n664_), .A2(new_n666_), .ZN(new_n667_));
  XOR2_X1   g466(.A(new_n667_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g467(.A(G15gat), .B1(new_n658_), .B2(new_n602_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT41), .Z(new_n670_));
  NAND3_X1  g469(.A1(new_n645_), .A2(new_n581_), .A3(new_n601_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(G1326gat));
  INV_X1    g471(.A(G22gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n645_), .A2(new_n673_), .A3(new_n424_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G22gat), .B1(new_n658_), .B2(new_n604_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n675_), .A2(KEYINPUT42), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(KEYINPUT42), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n674_), .B1(new_n676_), .B2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT102), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  OAI211_X1 g479(.A(KEYINPUT102), .B(new_n674_), .C1(new_n676_), .C2(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1327gat));
  NAND2_X1  g481(.A1(new_n655_), .A2(new_n331_), .ZN(new_n683_));
  NOR4_X1   g482(.A1(new_n654_), .A2(new_n648_), .A3(new_n268_), .A4(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(G29gat), .B1(new_n684_), .B2(new_n571_), .ZN(new_n685_));
  INV_X1    g484(.A(KEYINPUT44), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n268_), .A2(new_n332_), .A3(new_n648_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(KEYINPUT43), .B1(new_n654_), .B2(new_n299_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT43), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n297_), .A2(new_n298_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n619_), .A2(new_n690_), .A3(new_n691_), .ZN(new_n692_));
  AOI21_X1  g491(.A(new_n688_), .B1(new_n689_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n686_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  AOI211_X1 g494(.A(KEYINPUT103), .B(new_n688_), .C1(new_n689_), .C2(new_n692_), .ZN(new_n696_));
  OAI21_X1  g495(.A(KEYINPUT104), .B1(new_n695_), .B2(new_n696_), .ZN(new_n697_));
  NOR3_X1   g496(.A1(new_n654_), .A2(KEYINPUT43), .A3(new_n299_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n690_), .B1(new_n619_), .B2(new_n691_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n687_), .B1(new_n698_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT103), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT104), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n689_), .A2(new_n692_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n703_), .A2(new_n694_), .A3(new_n687_), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n701_), .A2(new_n702_), .A3(new_n686_), .A4(new_n704_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n697_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n693_), .A2(KEYINPUT44), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n708_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n571_), .A2(G29gat), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n685_), .B1(new_n709_), .B2(new_n710_), .ZN(G1328gat));
  INV_X1    g510(.A(G36gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n684_), .A2(new_n712_), .A3(new_n663_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT45), .Z(new_n714_));
  NAND3_X1  g513(.A1(new_n706_), .A2(new_n663_), .A3(new_n707_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n715_), .B2(G36gat), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT105), .B(KEYINPUT46), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n716_), .B(new_n718_), .ZN(G1329gat));
  NAND2_X1  g518(.A1(new_n601_), .A2(G43gat), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n684_), .A2(new_n601_), .ZN(new_n721_));
  OAI22_X1  g520(.A1(new_n708_), .A2(new_n720_), .B1(G43gat), .B2(new_n721_), .ZN(new_n722_));
  XNOR2_X1  g521(.A(new_n722_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g522(.A(G50gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n684_), .A2(new_n724_), .A3(new_n424_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n707_), .A2(new_n424_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT44), .B1(new_n700_), .B2(KEYINPUT103), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n702_), .B1(new_n728_), .B2(new_n704_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n695_), .A2(KEYINPUT104), .A3(new_n696_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n727_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT106), .B1(new_n731_), .B2(G50gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n726_), .B1(new_n697_), .B2(new_n705_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n724_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n725_), .B1(new_n732_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(KEYINPUT107), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n738_));
  OAI211_X1 g537(.A(new_n738_), .B(new_n725_), .C1(new_n732_), .C2(new_n735_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n737_), .A2(new_n739_), .ZN(G1331gat));
  INV_X1    g539(.A(new_n268_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n333_), .A2(new_n741_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n654_), .A2(new_n644_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  OR3_X1    g543(.A1(new_n744_), .A2(G57gat), .A3(new_n659_), .ZN(new_n745_));
  NAND4_X1  g544(.A1(new_n656_), .A2(new_n269_), .A3(new_n648_), .A4(new_n332_), .ZN(new_n746_));
  OAI21_X1  g545(.A(G57gat), .B1(new_n746_), .B2(new_n659_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n745_), .A2(new_n747_), .ZN(G1332gat));
  OAI21_X1  g547(.A(G64gat), .B1(new_n746_), .B2(new_n662_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT48), .ZN(new_n750_));
  OR2_X1    g549(.A1(new_n662_), .A2(G64gat), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n744_), .B2(new_n751_), .ZN(G1333gat));
  OAI21_X1  g551(.A(G71gat), .B1(new_n746_), .B2(new_n602_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT49), .ZN(new_n754_));
  OR2_X1    g553(.A1(new_n602_), .A2(G71gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n744_), .B2(new_n755_), .ZN(G1334gat));
  OAI21_X1  g555(.A(G78gat), .B1(new_n746_), .B2(new_n604_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT50), .ZN(new_n758_));
  OR2_X1    g557(.A1(new_n604_), .A2(G78gat), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n758_), .B1(new_n744_), .B2(new_n759_), .ZN(G1335gat));
  NAND4_X1  g559(.A1(new_n703_), .A2(new_n648_), .A3(new_n268_), .A4(new_n331_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761_), .B2(new_n659_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n269_), .ZN(new_n763_));
  NOR4_X1   g562(.A1(new_n763_), .A2(new_n654_), .A3(new_n644_), .A4(new_n683_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n209_), .A3(new_n571_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n762_), .A2(new_n765_), .ZN(G1336gat));
  OAI21_X1  g565(.A(G92gat), .B1(new_n761_), .B2(new_n662_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n764_), .A2(new_n210_), .A3(new_n663_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(G1337gat));
  OAI21_X1  g568(.A(G99gat), .B1(new_n761_), .B2(new_n602_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n764_), .A2(new_n202_), .A3(new_n601_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR2_X1   g572(.A1(new_n761_), .A2(new_n604_), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n774_), .A2(KEYINPUT109), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n203_), .B1(new_n774_), .B2(KEYINPUT109), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(KEYINPUT52), .A3(new_n776_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n764_), .A2(new_n203_), .A3(new_n424_), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n778_), .B(KEYINPUT108), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n777_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n775_), .A2(new_n776_), .ZN(new_n783_));
  OAI211_X1 g582(.A(new_n781_), .B(new_n782_), .C1(KEYINPUT52), .C2(new_n783_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(KEYINPUT52), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT53), .B1(new_n785_), .B2(new_n780_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  INV_X1    g586(.A(new_n249_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n219_), .B1(new_n283_), .B2(new_n212_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n252_), .B1(new_n789_), .B2(KEYINPUT12), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n242_), .A2(KEYINPUT68), .A3(new_n250_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n788_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n245_), .B1(new_n792_), .B2(new_n239_), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n254_), .A2(new_n794_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n793_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT112), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n254_), .A2(new_n797_), .A3(new_n794_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n797_), .B1(new_n254_), .B2(new_n794_), .ZN(new_n799_));
  INV_X1    g598(.A(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n796_), .A2(new_n798_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n259_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT56), .ZN(new_n803_));
  NOR3_X1   g602(.A1(new_n799_), .A2(new_n793_), .A3(new_n795_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n261_), .B1(new_n804_), .B2(new_n798_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n320_), .A2(new_n632_), .ZN(new_n808_));
  OR3_X1    g607(.A1(new_n808_), .A2(KEYINPUT114), .A3(new_n624_), .ZN(new_n809_));
  OAI21_X1  g608(.A(KEYINPUT114), .B1(new_n808_), .B2(new_n624_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n809_), .A2(new_n629_), .A3(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n636_), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n625_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT115), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n811_), .A2(new_n816_), .A3(new_n812_), .A4(new_n813_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n815_), .A2(new_n637_), .A3(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n262_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n803_), .A2(new_n807_), .A3(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT58), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n299_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n821_), .A2(new_n822_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n826_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n825_), .A2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n806_), .B1(new_n805_), .B2(KEYINPUT113), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n802_), .A2(new_n830_), .A3(KEYINPUT56), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n644_), .A2(new_n262_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT111), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n832_), .A2(new_n833_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n644_), .A2(KEYINPUT111), .A3(new_n262_), .ZN(new_n835_));
  NAND4_X1  g634(.A1(new_n829_), .A2(new_n831_), .A3(new_n834_), .A4(new_n835_), .ZN(new_n836_));
  OR2_X1    g635(.A1(new_n263_), .A2(new_n818_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n295_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(KEYINPUT116), .B(KEYINPUT57), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n655_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT118), .ZN(new_n843_));
  AND3_X1   g642(.A1(new_n842_), .A2(new_n843_), .A3(KEYINPUT57), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n843_), .B1(new_n842_), .B2(KEYINPUT57), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n828_), .B(new_n841_), .C1(new_n844_), .C2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n331_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n741_), .A2(new_n299_), .A3(new_n648_), .A4(new_n332_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n847_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT59), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n617_), .A2(new_n571_), .A3(new_n601_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n852_), .A2(new_n853_), .A3(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n644_), .A2(G113gat), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(KEYINPUT120), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT119), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n844_), .A2(new_n845_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n821_), .A2(new_n822_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n861_), .A2(new_n824_), .A3(new_n691_), .ZN(new_n862_));
  INV_X1    g661(.A(new_n826_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n823_), .A2(new_n824_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n840_), .ZN(new_n866_));
  OAI22_X1  g665(.A1(new_n864_), .A2(new_n865_), .B1(new_n842_), .B2(new_n866_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n859_), .B1(new_n860_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869_));
  OAI21_X1  g668(.A(KEYINPUT118), .B1(new_n839_), .B2(new_n869_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n842_), .A2(new_n843_), .A3(KEYINPUT57), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  AOI22_X1  g671(.A1(new_n825_), .A2(new_n827_), .B1(new_n839_), .B2(new_n840_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(new_n873_), .A3(KEYINPUT119), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n868_), .A2(new_n331_), .A3(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n854_), .B1(new_n875_), .B2(new_n851_), .ZN(new_n876_));
  OAI211_X1 g675(.A(new_n856_), .B(new_n858_), .C1(new_n876_), .C2(new_n853_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(G113gat), .B1(new_n876_), .B2(new_n644_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n878_), .A2(new_n879_), .ZN(G1340gat));
  OAI21_X1  g679(.A(new_n856_), .B1(new_n876_), .B2(new_n853_), .ZN(new_n881_));
  OAI21_X1  g680(.A(G120gat), .B1(new_n881_), .B2(new_n763_), .ZN(new_n882_));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n741_), .B2(KEYINPUT60), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n876_), .B(new_n884_), .C1(KEYINPUT60), .C2(new_n883_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n882_), .A2(new_n885_), .ZN(G1341gat));
  OAI21_X1  g685(.A(G127gat), .B1(new_n881_), .B2(new_n331_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n876_), .A2(new_n427_), .A3(new_n332_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1342gat));
  NOR2_X1   g688(.A1(new_n299_), .A2(new_n425_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(KEYINPUT121), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n856_), .B(new_n891_), .C1(new_n876_), .C2(new_n853_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(G134gat), .B1(new_n876_), .B2(new_n655_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1343gat));
  NOR2_X1   g694(.A1(new_n604_), .A2(new_n601_), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n896_), .A2(new_n571_), .A3(new_n662_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n897_), .B1(new_n875_), .B2(new_n851_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(new_n644_), .ZN(new_n899_));
  XNOR2_X1  g698(.A(new_n899_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g699(.A1(new_n898_), .A2(new_n269_), .ZN(new_n901_));
  XNOR2_X1  g700(.A(new_n901_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g701(.A1(new_n898_), .A2(new_n332_), .ZN(new_n903_));
  XNOR2_X1  g702(.A(KEYINPUT61), .B(G155gat), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n903_), .B(new_n904_), .ZN(G1346gat));
  INV_X1    g704(.A(KEYINPUT122), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n353_), .B1(new_n898_), .B2(new_n691_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n655_), .A2(new_n353_), .ZN(new_n908_));
  AOI211_X1 g707(.A(new_n897_), .B(new_n908_), .C1(new_n875_), .C2(new_n851_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n906_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n898_), .A2(new_n353_), .A3(new_n655_), .ZN(new_n911_));
  AOI211_X1 g710(.A(new_n299_), .B(new_n897_), .C1(new_n875_), .C2(new_n851_), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n911_), .B(KEYINPUT122), .C1(new_n912_), .C2(new_n353_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n913_), .ZN(G1347gat));
  NOR2_X1   g713(.A1(new_n662_), .A2(new_n571_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n601_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n916_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n852_), .A2(new_n604_), .A3(new_n644_), .A4(new_n917_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n514_), .A2(new_n504_), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n918_), .A2(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(KEYINPUT123), .B1(new_n918_), .B2(G169gat), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT62), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n332_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n924_));
  OAI211_X1 g723(.A(new_n604_), .B(new_n917_), .C1(new_n924_), .C2(new_n850_), .ZN(new_n925_));
  OAI21_X1  g724(.A(G169gat), .B1(new_n925_), .B2(new_n648_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT123), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n926_), .A2(new_n927_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n918_), .A2(KEYINPUT123), .A3(G169gat), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n928_), .A2(new_n929_), .A3(KEYINPUT62), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n923_), .A2(new_n930_), .ZN(G1348gat));
  INV_X1    g730(.A(KEYINPUT124), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n925_), .A2(new_n741_), .ZN(new_n933_));
  NOR2_X1   g732(.A1(new_n933_), .A2(G176gat), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n875_), .A2(new_n851_), .ZN(new_n935_));
  NOR3_X1   g734(.A1(new_n763_), .A2(new_n513_), .A3(new_n916_), .ZN(new_n936_));
  AND3_X1   g735(.A1(new_n935_), .A2(new_n604_), .A3(new_n936_), .ZN(new_n937_));
  OAI21_X1  g736(.A(new_n932_), .B1(new_n934_), .B2(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n424_), .B1(new_n875_), .B2(new_n851_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n939_), .A2(new_n936_), .ZN(new_n940_));
  OAI211_X1 g739(.A(new_n940_), .B(KEYINPUT124), .C1(G176gat), .C2(new_n933_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n938_), .A2(new_n941_), .ZN(G1349gat));
  NOR2_X1   g741(.A1(new_n916_), .A2(new_n331_), .ZN(new_n943_));
  AOI21_X1  g742(.A(G183gat), .B1(new_n939_), .B2(new_n943_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n424_), .B1(new_n847_), .B2(new_n851_), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n916_), .A2(new_n485_), .A3(new_n331_), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n944_), .B1(new_n945_), .B2(new_n946_), .ZN(G1350gat));
  OAI21_X1  g746(.A(G190gat), .B1(new_n925_), .B2(new_n299_), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n655_), .A2(new_n497_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n925_), .B2(new_n949_), .ZN(G1351gat));
  NAND2_X1  g749(.A1(KEYINPUT125), .A2(G197gat), .ZN(new_n951_));
  XOR2_X1   g750(.A(new_n951_), .B(KEYINPUT126), .Z(new_n952_));
  AND2_X1   g751(.A1(new_n915_), .A2(new_n896_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n935_), .A2(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(new_n954_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n644_), .B1(KEYINPUT125), .B2(G197gat), .ZN(new_n956_));
  INV_X1    g755(.A(new_n956_), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n952_), .B1(new_n955_), .B2(new_n957_), .ZN(new_n958_));
  INV_X1    g757(.A(new_n952_), .ZN(new_n959_));
  NOR3_X1   g758(.A1(new_n954_), .A2(new_n956_), .A3(new_n959_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(new_n958_), .A2(new_n960_), .ZN(G1352gat));
  XOR2_X1   g760(.A(KEYINPUT127), .B(G204gat), .Z(new_n962_));
  NAND3_X1  g761(.A1(new_n955_), .A2(new_n269_), .A3(new_n962_), .ZN(new_n963_));
  NOR2_X1   g762(.A1(new_n954_), .A2(new_n763_), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n965_));
  NOR2_X1   g764(.A1(new_n965_), .A2(G204gat), .ZN(new_n966_));
  OAI21_X1  g765(.A(new_n963_), .B1(new_n964_), .B2(new_n966_), .ZN(G1353gat));
  XNOR2_X1  g766(.A(KEYINPUT63), .B(G211gat), .ZN(new_n968_));
  NOR3_X1   g767(.A1(new_n954_), .A2(new_n331_), .A3(new_n968_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n955_), .A2(new_n332_), .ZN(new_n970_));
  NOR2_X1   g769(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n971_));
  AOI21_X1  g770(.A(new_n969_), .B1(new_n970_), .B2(new_n971_), .ZN(G1354gat));
  OAI21_X1  g771(.A(G218gat), .B1(new_n954_), .B2(new_n299_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n655_), .A2(new_n377_), .ZN(new_n974_));
  OAI21_X1  g773(.A(new_n973_), .B1(new_n954_), .B2(new_n974_), .ZN(G1355gat));
endmodule


