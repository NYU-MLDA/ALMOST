//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 0 0 1 0 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n759_, new_n760_, new_n761_, new_n762_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n783_, new_n784_, new_n785_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n895_, new_n896_, new_n897_, new_n899_,
    new_n900_, new_n902_, new_n903_, new_n904_, new_n905_, new_n906_,
    new_n907_, new_n908_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n917_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_;
  AOI21_X1  g000(.A(G176gat), .B1(KEYINPUT82), .B2(KEYINPUT22), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G169gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(G183gat), .A2(G190gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT23), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NAND3_X1  g005(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n207_));
  OAI211_X1 g006(.A(new_n206_), .B(new_n207_), .C1(G183gat), .C2(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n203_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(KEYINPUT26), .B(G190gat), .ZN(new_n210_));
  INV_X1    g009(.A(G183gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(KEYINPUT80), .A3(KEYINPUT25), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT80), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT25), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n213_), .B1(new_n214_), .B2(G183gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n210_), .A2(new_n212_), .A3(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT81), .ZN(new_n217_));
  OAI21_X1  g016(.A(G183gat), .B1(new_n217_), .B2(KEYINPUT25), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n214_), .A2(KEYINPUT81), .ZN(new_n219_));
  NOR2_X1   g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n216_), .A2(new_n220_), .ZN(new_n221_));
  NOR3_X1   g020(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n223_));
  INV_X1    g022(.A(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(G169gat), .A2(G176gat), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n222_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n204_), .A2(KEYINPUT23), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n205_), .A2(G183gat), .A3(G190gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n226_), .A2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n209_), .B1(new_n221_), .B2(new_n230_), .ZN(new_n231_));
  XOR2_X1   g030(.A(KEYINPUT83), .B(KEYINPUT30), .Z(new_n232_));
  XNOR2_X1  g031(.A(new_n231_), .B(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n233_), .B(KEYINPUT84), .Z(new_n234_));
  XNOR2_X1  g033(.A(G71gat), .B(G99gat), .ZN(new_n235_));
  INV_X1    g034(.A(G43gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(new_n235_), .B(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G227gat), .A2(G233gat), .ZN(new_n238_));
  INV_X1    g037(.A(G15gat), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n237_), .B(new_n240_), .ZN(new_n241_));
  NOR2_X1   g040(.A1(new_n234_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n233_), .A2(KEYINPUT84), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n242_), .B1(new_n243_), .B2(new_n241_), .ZN(new_n244_));
  INV_X1    g043(.A(G134gat), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G127gat), .ZN(new_n246_));
  INV_X1    g045(.A(G127gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n247_), .A2(G134gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(G120gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G113gat), .ZN(new_n251_));
  INV_X1    g050(.A(G113gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(G120gat), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n251_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n249_), .A2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n246_), .A2(new_n248_), .A3(new_n251_), .A4(new_n253_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(KEYINPUT85), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n249_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT85), .ZN(new_n259_));
  NAND4_X1  g058(.A1(new_n258_), .A2(new_n259_), .A3(new_n251_), .A4(new_n253_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n257_), .A2(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n261_), .B(KEYINPUT31), .ZN(new_n262_));
  OR2_X1    g061(.A1(new_n244_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n244_), .A2(new_n262_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(G8gat), .B(G36gat), .Z(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT18), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G64gat), .B(G92gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n267_), .B(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT95), .B(KEYINPUT19), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G226gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n271_), .B(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT20), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT90), .ZN(new_n275_));
  AND2_X1   g074(.A1(KEYINPUT88), .A2(G197gat), .ZN(new_n276_));
  NOR2_X1   g075(.A1(KEYINPUT88), .A2(G197gat), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n276_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT89), .ZN(new_n279_));
  INV_X1    g078(.A(G197gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n279_), .B1(new_n280_), .B2(G204gat), .ZN(new_n281_));
  INV_X1    g080(.A(G204gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n278_), .A2(G204gat), .B1(new_n281_), .B2(new_n283_), .ZN(new_n284_));
  XOR2_X1   g083(.A(G211gat), .B(G218gat), .Z(new_n285_));
  NAND2_X1  g084(.A1(new_n285_), .A2(KEYINPUT21), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n275_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n281_), .A2(new_n283_), .ZN(new_n288_));
  OR2_X1    g087(.A1(KEYINPUT88), .A2(G197gat), .ZN(new_n289_));
  NAND2_X1  g088(.A1(KEYINPUT88), .A2(G197gat), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n289_), .A2(G204gat), .A3(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n288_), .A2(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G211gat), .B(G218gat), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT21), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n292_), .A2(KEYINPUT90), .A3(new_n295_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n288_), .A2(new_n291_), .A3(new_n294_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n289_), .A2(new_n282_), .A3(new_n290_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n294_), .B1(G197gat), .B2(G204gat), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n285_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  AOI22_X1  g099(.A1(new_n287_), .A2(new_n296_), .B1(new_n297_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n230_), .ZN(new_n302_));
  OR2_X1    g101(.A1(new_n218_), .A2(new_n219_), .ZN(new_n303_));
  NAND4_X1  g102(.A1(new_n303_), .A2(new_n212_), .A3(new_n210_), .A4(new_n215_), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n302_), .A2(new_n304_), .B1(new_n208_), .B2(new_n203_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n274_), .B1(new_n301_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n300_), .A2(new_n297_), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n292_), .A2(KEYINPUT90), .A3(new_n295_), .ZN(new_n308_));
  AOI21_X1  g107(.A(KEYINPUT90), .B1(new_n292_), .B2(new_n295_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n307_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n225_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT22), .B(G169gat), .ZN(new_n312_));
  INV_X1    g111(.A(G176gat), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n314_), .A2(new_n208_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT25), .B(G183gat), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n210_), .A2(new_n316_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n317_));
  AND2_X1   g116(.A1(new_n317_), .A2(new_n226_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n310_), .B1(new_n315_), .B2(new_n318_), .ZN(new_n319_));
  AOI21_X1  g118(.A(new_n273_), .B1(new_n306_), .B2(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(KEYINPUT20), .B1(new_n301_), .B2(new_n305_), .ZN(new_n321_));
  AOI22_X1  g120(.A1(new_n317_), .A2(new_n226_), .B1(new_n314_), .B2(new_n208_), .ZN(new_n322_));
  OAI211_X1 g121(.A(new_n322_), .B(new_n307_), .C1(new_n308_), .C2(new_n309_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n273_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n321_), .A2(new_n324_), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n270_), .B1(new_n320_), .B2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n273_), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT20), .B1(new_n310_), .B2(new_n231_), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n301_), .A2(new_n322_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n327_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n274_), .B1(new_n310_), .B2(new_n231_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n331_), .A2(new_n273_), .A3(new_n323_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n269_), .A3(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n326_), .A2(KEYINPUT96), .A3(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT96), .ZN(new_n335_));
  OAI211_X1 g134(.A(new_n335_), .B(new_n270_), .C1(new_n320_), .C2(new_n325_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT97), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT97), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n334_), .A2(new_n339_), .A3(new_n336_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G141gat), .ZN(new_n342_));
  INV_X1    g141(.A(G148gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(new_n343_), .A3(KEYINPUT3), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(G141gat), .B2(G148gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT2), .ZN(new_n350_));
  AOI22_X1  g149(.A1(new_n348_), .A2(KEYINPUT86), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT86), .ZN(new_n352_));
  NAND4_X1  g151(.A1(new_n352_), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n347_), .A2(new_n351_), .A3(new_n353_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G155gat), .B(G162gat), .Z(new_n355_));
  INV_X1    g154(.A(KEYINPUT1), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n342_), .A2(new_n343_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n358_), .A2(new_n349_), .A3(new_n359_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n354_), .A2(new_n355_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n361_));
  OR3_X1    g160(.A1(new_n261_), .A2(new_n361_), .A3(KEYINPUT4), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT98), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n366_), .B1(new_n261_), .B2(new_n361_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n354_), .A2(new_n355_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n357_), .A2(new_n360_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n257_), .A2(new_n260_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(KEYINPUT98), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n367_), .A2(new_n372_), .ZN(new_n373_));
  AND2_X1   g172(.A1(new_n255_), .A2(new_n256_), .ZN(new_n374_));
  OR2_X1    g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  NAND4_X1  g174(.A1(new_n373_), .A2(KEYINPUT99), .A3(KEYINPUT4), .A4(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n370_), .A2(new_n374_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(new_n367_), .B2(new_n372_), .ZN(new_n379_));
  AOI21_X1  g178(.A(KEYINPUT99), .B1(new_n379_), .B2(KEYINPUT4), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n365_), .B1(new_n377_), .B2(new_n380_), .ZN(new_n381_));
  AND2_X1   g180(.A1(new_n379_), .A2(new_n363_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G85gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT0), .B(G57gat), .ZN(new_n386_));
  XOR2_X1   g185(.A(new_n385_), .B(new_n386_), .Z(new_n387_));
  AND2_X1   g186(.A1(new_n387_), .A2(KEYINPUT33), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n381_), .A2(new_n383_), .A3(new_n388_), .ZN(new_n389_));
  AND3_X1   g188(.A1(new_n370_), .A2(KEYINPUT98), .A3(new_n371_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT98), .B1(new_n370_), .B2(new_n371_), .ZN(new_n391_));
  OAI211_X1 g190(.A(KEYINPUT4), .B(new_n375_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT99), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n394_), .A2(new_n376_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n362_), .A2(new_n363_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n395_), .A2(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n387_), .B1(new_n379_), .B2(new_n364_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n387_), .ZN(new_n400_));
  AOI211_X1 g199(.A(new_n382_), .B(new_n400_), .C1(new_n395_), .C2(new_n365_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n389_), .B(new_n399_), .C1(new_n401_), .C2(KEYINPUT33), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT100), .B1(new_n341_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n389_), .A2(new_n399_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n382_), .B1(new_n395_), .B2(new_n365_), .ZN(new_n405_));
  AOI21_X1  g204(.A(KEYINPUT33), .B1(new_n405_), .B2(new_n387_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n404_), .A2(new_n406_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n334_), .A2(new_n339_), .A3(new_n336_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n339_), .B1(new_n334_), .B2(new_n336_), .ZN(new_n409_));
  NOR2_X1   g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT100), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n407_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n269_), .A2(KEYINPUT32), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n330_), .A2(new_n332_), .A3(new_n413_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n306_), .A2(new_n319_), .A3(new_n273_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n301_), .A2(KEYINPUT91), .ZN(new_n416_));
  INV_X1    g215(.A(KEYINPUT91), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n310_), .A2(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n416_), .A2(new_n418_), .A3(new_n322_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n273_), .B1(new_n419_), .B2(new_n331_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT101), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n415_), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(new_n421_), .B2(new_n420_), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n405_), .A2(new_n387_), .ZN(new_n424_));
  OAI221_X1 g223(.A(new_n414_), .B1(new_n423_), .B2(new_n413_), .C1(new_n424_), .C2(new_n401_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n403_), .A2(new_n412_), .A3(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT102), .ZN(new_n427_));
  OR3_X1    g226(.A1(new_n370_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n428_));
  OAI21_X1  g227(.A(KEYINPUT28), .B1(new_n370_), .B2(KEYINPUT29), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n428_), .A2(new_n429_), .ZN(new_n430_));
  XNOR2_X1  g229(.A(G22gat), .B(G50gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n430_), .B(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n370_), .A2(KEYINPUT29), .ZN(new_n433_));
  INV_X1    g232(.A(G233gat), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT87), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n435_), .A2(G228gat), .ZN(new_n436_));
  INV_X1    g235(.A(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n435_), .A2(G228gat), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n434_), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n310_), .A2(new_n433_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  NOR2_X1   g241(.A1(new_n310_), .A2(new_n417_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n287_), .A2(new_n296_), .ZN(new_n444_));
  AOI21_X1  g243(.A(KEYINPUT91), .B1(new_n444_), .B2(new_n307_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n433_), .B1(new_n443_), .B2(new_n445_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n442_), .B1(new_n446_), .B2(new_n439_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(G78gat), .B(G106gat), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n433_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n451_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n441_), .B1(new_n452_), .B2(new_n440_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n448_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n432_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n450_), .A2(new_n432_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n448_), .B1(new_n447_), .B2(KEYINPUT92), .ZN(new_n458_));
  OAI211_X1 g257(.A(KEYINPUT92), .B(new_n441_), .C1(new_n452_), .C2(new_n440_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NOR3_X1   g259(.A1(new_n458_), .A2(KEYINPUT93), .A3(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT93), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT92), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n449_), .B1(new_n453_), .B2(new_n463_), .ZN(new_n464_));
  AOI21_X1  g263(.A(new_n462_), .B1(new_n464_), .B2(new_n459_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n457_), .B1(new_n461_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT94), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(KEYINPUT93), .B1(new_n458_), .B2(new_n460_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n464_), .A2(new_n462_), .A3(new_n459_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(KEYINPUT94), .A3(new_n457_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n455_), .B1(new_n468_), .B2(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n426_), .A2(new_n427_), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n455_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT94), .B1(new_n471_), .B2(new_n457_), .ZN(new_n476_));
  AOI211_X1 g275(.A(new_n467_), .B(new_n456_), .C1(new_n469_), .C2(new_n470_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  OAI211_X1 g277(.A(KEYINPUT27), .B(new_n333_), .C1(new_n423_), .C2(new_n269_), .ZN(new_n479_));
  OR2_X1    g278(.A1(new_n337_), .A2(KEYINPUT27), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n424_), .A2(new_n401_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n478_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n474_), .A2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n427_), .B1(new_n426_), .B2(new_n473_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n265_), .B1(new_n485_), .B2(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT103), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n478_), .A2(new_n481_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n483_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n265_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(KEYINPUT103), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n493_), .B(new_n265_), .C1(new_n485_), .C2(new_n486_), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n488_), .A2(new_n492_), .A3(new_n494_), .ZN(new_n495_));
  XOR2_X1   g294(.A(G15gat), .B(G22gat), .Z(new_n496_));
  NAND2_X1  g295(.A1(G1gat), .A2(G8gat), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(KEYINPUT14), .B2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(new_n498_), .B(KEYINPUT75), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n499_), .B(KEYINPUT76), .ZN(new_n500_));
  XOR2_X1   g299(.A(G1gat), .B(G8gat), .Z(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT76), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n499_), .B(new_n503_), .ZN(new_n504_));
  INV_X1    g303(.A(new_n501_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n502_), .A2(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(G29gat), .B(G36gat), .Z(new_n508_));
  XOR2_X1   g307(.A(G43gat), .B(G50gat), .Z(new_n509_));
  OR2_X1    g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n509_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT78), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n507_), .A2(new_n514_), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n502_), .A2(new_n506_), .A3(new_n513_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n518_), .B(KEYINPUT79), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  AOI21_X1  g320(.A(new_n521_), .B1(new_n507_), .B2(new_n514_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n512_), .B(KEYINPUT15), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n502_), .A2(new_n506_), .A3(new_n523_), .ZN(new_n524_));
  AOI22_X1  g323(.A1(new_n517_), .A2(new_n519_), .B1(new_n522_), .B2(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(G113gat), .B(G141gat), .Z(new_n526_));
  XNOR2_X1  g325(.A(G169gat), .B(G197gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  XNOR2_X1  g327(.A(new_n525_), .B(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G120gat), .B(G148gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT5), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  NAND2_X1  g332(.A1(G230gat), .A2(G233gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT64), .Z(new_n535_));
  AND2_X1   g334(.A1(G85gat), .A2(G92gat), .ZN(new_n536_));
  NOR2_X1   g335(.A1(G85gat), .A2(G92gat), .ZN(new_n537_));
  NOR3_X1   g336(.A1(new_n536_), .A2(new_n537_), .A3(KEYINPUT8), .ZN(new_n538_));
  NAND2_X1  g337(.A1(G99gat), .A2(G106gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT6), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT67), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(G99gat), .ZN(new_n543_));
  INV_X1    g342(.A(G106gat), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n543_), .A2(new_n544_), .A3(KEYINPUT68), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(KEYINPUT7), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n538_), .B1(new_n542_), .B2(new_n546_), .ZN(new_n547_));
  OR2_X1    g346(.A1(new_n545_), .A2(KEYINPUT7), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(KEYINPUT7), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n540_), .A3(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT69), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n536_), .A2(new_n537_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n550_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT8), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n551_), .B1(new_n550_), .B2(new_n552_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n547_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n557_), .A2(KEYINPUT11), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n557_), .A2(KEYINPUT11), .ZN(new_n559_));
  XOR2_X1   g358(.A(G71gat), .B(G78gat), .Z(new_n560_));
  NAND3_X1  g359(.A1(new_n558_), .A2(new_n559_), .A3(new_n560_), .ZN(new_n561_));
  OR2_X1    g360(.A1(new_n559_), .A2(new_n560_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n542_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT66), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n536_), .B1(new_n565_), .B2(KEYINPUT9), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n565_), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n566_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(KEYINPUT10), .B(G99gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n569_), .B(KEYINPUT65), .ZN(new_n570_));
  OAI211_X1 g369(.A(new_n564_), .B(new_n568_), .C1(G106gat), .C2(new_n570_), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n556_), .A2(new_n563_), .A3(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n563_), .B1(new_n556_), .B2(new_n571_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT12), .ZN(new_n575_));
  NOR3_X1   g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n575_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  OAI21_X1  g377(.A(new_n535_), .B1(new_n576_), .B2(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n574_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n535_), .B1(new_n580_), .B2(new_n572_), .ZN(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT70), .B1(new_n579_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n535_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n580_), .A2(KEYINPUT12), .A3(new_n572_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n584_), .B1(new_n585_), .B2(new_n577_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT70), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n586_), .A2(new_n587_), .A3(new_n581_), .ZN(new_n588_));
  OAI21_X1  g387(.A(new_n533_), .B1(new_n583_), .B2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n533_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n579_), .A2(new_n590_), .A3(new_n582_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n589_), .A2(KEYINPUT71), .A3(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT71), .ZN(new_n593_));
  OAI211_X1 g392(.A(new_n593_), .B(new_n533_), .C1(new_n583_), .C2(new_n588_), .ZN(new_n594_));
  AND2_X1   g393(.A1(new_n592_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT13), .ZN(new_n596_));
  OR3_X1    g395(.A1(new_n595_), .A2(KEYINPUT72), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(KEYINPUT72), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n596_), .A2(KEYINPUT72), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n595_), .A2(new_n598_), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n597_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(G190gat), .B(G218gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(G134gat), .B(G162gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT36), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n556_), .A2(new_n571_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n523_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT34), .ZN(new_n612_));
  INV_X1    g411(.A(new_n512_), .ZN(new_n613_));
  OAI221_X1 g412(.A(new_n610_), .B1(KEYINPUT35), .B2(new_n612_), .C1(new_n613_), .C2(new_n609_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(KEYINPUT35), .ZN(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  OR2_X1    g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n616_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT73), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n608_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n617_), .A2(KEYINPUT73), .A3(new_n618_), .A4(new_n607_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n621_), .A2(new_n622_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n619_), .A2(KEYINPUT36), .A3(new_n606_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT74), .B(KEYINPUT37), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n625_), .B(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(G231gat), .A2(G233gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n563_), .B(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n507_), .A2(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(G127gat), .B(G155gat), .Z(new_n633_));
  XNOR2_X1  g432(.A(new_n633_), .B(KEYINPUT16), .ZN(new_n634_));
  XNOR2_X1  g433(.A(G183gat), .B(G211gat), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT17), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n502_), .A2(new_n506_), .A3(new_n630_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n632_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT77), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n632_), .A2(new_n639_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n636_), .B(KEYINPUT17), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n641_), .A2(new_n644_), .ZN(new_n645_));
  NOR2_X1   g444(.A1(new_n628_), .A2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n495_), .A2(new_n529_), .A3(new_n603_), .A4(new_n646_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n647_), .A2(G1gat), .A3(new_n483_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n649_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n650_), .A2(KEYINPUT38), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT38), .B1(new_n650_), .B2(new_n651_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n529_), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n602_), .A2(new_n654_), .A3(new_n645_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n625_), .B(KEYINPUT105), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n495_), .A2(new_n655_), .A3(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(G1gat), .B1(new_n657_), .B2(new_n483_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT106), .ZN(new_n659_));
  OR3_X1    g458(.A1(new_n652_), .A2(new_n653_), .A3(new_n659_), .ZN(G1324gat));
  INV_X1    g459(.A(new_n647_), .ZN(new_n661_));
  INV_X1    g460(.A(G8gat), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n662_), .A3(new_n481_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT39), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n657_), .A2(new_n482_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n662_), .B1(new_n665_), .B2(KEYINPUT107), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT107), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n667_), .B1(new_n657_), .B2(new_n482_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n664_), .B1(new_n666_), .B2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n494_), .A2(new_n492_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n426_), .A2(new_n473_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT102), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n672_), .A2(new_n484_), .A3(new_n474_), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n493_), .B1(new_n673_), .B2(new_n265_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n670_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n656_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND4_X1  g476(.A1(new_n677_), .A2(KEYINPUT107), .A3(new_n481_), .A4(new_n655_), .ZN(new_n678_));
  AND4_X1   g477(.A1(new_n664_), .A2(new_n678_), .A3(new_n668_), .A4(G8gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n663_), .B1(new_n669_), .B2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(KEYINPUT108), .B(KEYINPUT40), .ZN(new_n681_));
  INV_X1    g480(.A(new_n681_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(new_n683_));
  OAI211_X1 g482(.A(new_n663_), .B(new_n681_), .C1(new_n669_), .C2(new_n679_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1325gat));
  OAI21_X1  g484(.A(G15gat), .B1(new_n657_), .B2(new_n265_), .ZN(new_n686_));
  XOR2_X1   g485(.A(new_n686_), .B(KEYINPUT41), .Z(new_n687_));
  INV_X1    g486(.A(new_n265_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n661_), .A2(new_n239_), .A3(new_n688_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n687_), .A2(new_n689_), .ZN(G1326gat));
  OAI21_X1  g489(.A(G22gat), .B1(new_n657_), .B2(new_n473_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT42), .ZN(new_n692_));
  OR3_X1    g491(.A1(new_n647_), .A2(G22gat), .A3(new_n473_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT109), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(G1327gat));
  NOR2_X1   g495(.A1(new_n675_), .A2(new_n654_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n645_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n625_), .ZN(new_n699_));
  NOR3_X1   g498(.A1(new_n602_), .A2(new_n698_), .A3(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n697_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(G29gat), .B1(new_n702_), .B2(new_n490_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n628_), .B1(new_n670_), .B2(new_n674_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(KEYINPUT43), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n495_), .A2(new_n706_), .A3(new_n628_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  NOR3_X1   g507(.A1(new_n602_), .A2(new_n654_), .A3(new_n698_), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT44), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711_));
  INV_X1    g510(.A(new_n709_), .ZN(new_n712_));
  AOI211_X1 g511(.A(new_n711_), .B(new_n712_), .C1(new_n705_), .C2(new_n707_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n710_), .A2(new_n713_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n490_), .A2(G29gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n703_), .B1(new_n714_), .B2(new_n715_), .ZN(G1328gat));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n717_));
  INV_X1    g516(.A(G36gat), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n718_), .B1(new_n714_), .B2(new_n481_), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n697_), .A2(new_n718_), .A3(new_n481_), .A4(new_n700_), .ZN(new_n720_));
  XOR2_X1   g519(.A(KEYINPUT110), .B(KEYINPUT45), .Z(new_n721_));
  XNOR2_X1  g520(.A(new_n720_), .B(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n717_), .B1(new_n719_), .B2(new_n723_), .ZN(new_n724_));
  NOR3_X1   g523(.A1(new_n710_), .A2(new_n713_), .A3(new_n482_), .ZN(new_n725_));
  OAI211_X1 g524(.A(KEYINPUT46), .B(new_n722_), .C1(new_n725_), .C2(new_n718_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1329gat));
  AOI21_X1  g526(.A(G43gat), .B1(new_n702_), .B2(new_n688_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n265_), .A2(new_n236_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n728_), .B1(new_n714_), .B2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n731_));
  NOR2_X1   g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(new_n731_), .ZN(new_n733_));
  AOI211_X1 g532(.A(new_n733_), .B(new_n728_), .C1(new_n714_), .C2(new_n729_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1330gat));
  AOI21_X1  g534(.A(G50gat), .B1(new_n702_), .B2(new_n478_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n478_), .A2(G50gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n736_), .B1(new_n714_), .B2(new_n737_), .ZN(G1331gat));
  NAND2_X1  g537(.A1(new_n602_), .A2(new_n646_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT112), .ZN(new_n740_));
  NOR2_X1   g539(.A1(new_n675_), .A2(new_n529_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT113), .Z(new_n743_));
  AOI21_X1  g542(.A(G57gat), .B1(new_n743_), .B2(new_n490_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n529_), .A2(new_n645_), .ZN(new_n745_));
  AND2_X1   g544(.A1(new_n602_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n677_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(G57gat), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n749_), .B1(new_n490_), .B2(KEYINPUT114), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(KEYINPUT114), .B2(new_n749_), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n744_), .B1(new_n748_), .B2(new_n751_), .ZN(G1332gat));
  INV_X1    g551(.A(G64gat), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n743_), .A2(new_n753_), .A3(new_n481_), .ZN(new_n754_));
  OAI21_X1  g553(.A(G64gat), .B1(new_n747_), .B2(new_n482_), .ZN(new_n755_));
  XOR2_X1   g554(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n754_), .A2(new_n757_), .ZN(G1333gat));
  INV_X1    g557(.A(G71gat), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n743_), .A2(new_n759_), .A3(new_n688_), .ZN(new_n760_));
  OAI21_X1  g559(.A(G71gat), .B1(new_n747_), .B2(new_n265_), .ZN(new_n761_));
  XNOR2_X1  g560(.A(new_n761_), .B(KEYINPUT49), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1334gat));
  INV_X1    g562(.A(G78gat), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n743_), .A2(new_n764_), .A3(new_n478_), .ZN(new_n765_));
  OAI21_X1  g564(.A(G78gat), .B1(new_n747_), .B2(new_n473_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT50), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(G1335gat));
  NAND4_X1  g567(.A1(new_n741_), .A2(new_n602_), .A3(new_n645_), .A4(new_n625_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(G85gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n770_), .A2(new_n771_), .A3(new_n490_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n708_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n603_), .A2(new_n529_), .A3(new_n698_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  NOR3_X1   g574(.A1(new_n773_), .A2(new_n483_), .A3(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n776_), .B2(new_n771_), .ZN(G1336gat));
  AOI21_X1  g576(.A(G92gat), .B1(new_n770_), .B2(new_n481_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n773_), .A2(new_n775_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n481_), .A2(G92gat), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT116), .ZN(new_n781_));
  AOI21_X1  g580(.A(new_n778_), .B1(new_n779_), .B2(new_n781_), .ZN(G1337gat));
  OR3_X1    g581(.A1(new_n769_), .A2(new_n265_), .A3(new_n570_), .ZN(new_n783_));
  NOR3_X1   g582(.A1(new_n773_), .A2(new_n265_), .A3(new_n775_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n783_), .B1(new_n784_), .B2(new_n543_), .ZN(new_n785_));
  XNOR2_X1  g584(.A(new_n785_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g585(.A1(new_n770_), .A2(new_n544_), .A3(new_n478_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n708_), .A2(new_n478_), .A3(new_n774_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(KEYINPUT52), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n544_), .B1(new_n789_), .B2(KEYINPUT52), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n788_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n790_), .B1(new_n788_), .B2(new_n791_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n787_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n794_));
  XNOR2_X1  g593(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n794_), .A2(new_n796_), .ZN(new_n797_));
  OAI211_X1 g596(.A(new_n787_), .B(new_n795_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(G1339gat));
  NAND3_X1  g598(.A1(new_n489_), .A2(new_n688_), .A3(new_n490_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n800_), .A2(KEYINPUT59), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n528_), .B1(new_n517_), .B2(new_n520_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n515_), .A2(new_n524_), .A3(new_n521_), .ZN(new_n803_));
  AOI22_X1  g602(.A1(new_n525_), .A2(new_n528_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n587_), .B1(new_n586_), .B2(new_n581_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n579_), .A2(KEYINPUT70), .A3(new_n582_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n590_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n591_), .A2(KEYINPUT71), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n804_), .B(new_n594_), .C1(new_n807_), .C2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT121), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n579_), .A2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n586_), .A2(KEYINPUT55), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n585_), .A2(new_n584_), .A3(new_n577_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT120), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n585_), .A2(KEYINPUT120), .A3(new_n584_), .A4(new_n577_), .ZN(new_n817_));
  NAND4_X1  g616(.A1(new_n812_), .A2(new_n813_), .A3(new_n816_), .A4(new_n817_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n818_), .A2(KEYINPUT56), .A3(new_n533_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT56), .B1(new_n818_), .B2(new_n533_), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n529_), .B(new_n591_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT121), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n592_), .A2(new_n822_), .A3(new_n594_), .A4(new_n804_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n810_), .A2(new_n821_), .A3(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(new_n699_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n824_), .A2(KEYINPUT57), .A3(new_n699_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n591_), .B(new_n804_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830_));
  OR2_X1    g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n829_), .A2(new_n830_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n628_), .A2(new_n831_), .A3(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n827_), .A2(new_n828_), .A3(new_n833_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n834_), .A2(new_n645_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT119), .ZN(new_n836_));
  XNOR2_X1  g635(.A(new_n745_), .B(new_n836_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n625_), .B(new_n626_), .ZN(new_n838_));
  NAND4_X1  g637(.A1(new_n597_), .A2(new_n837_), .A3(new_n601_), .A4(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n839_), .B(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n801_), .B1(new_n835_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n834_), .A2(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n827_), .A2(new_n833_), .A3(KEYINPUT122), .A4(new_n828_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n645_), .A3(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n839_), .B(KEYINPUT54), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n800_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n842_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(G113gat), .B1(new_n850_), .B2(new_n654_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n848_), .A2(new_n252_), .A3(new_n529_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(G1340gat));
  OAI211_X1 g652(.A(new_n602_), .B(new_n842_), .C1(new_n848_), .C2(new_n849_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n250_), .B1(new_n603_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n848_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n250_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n855_), .A2(KEYINPUT123), .A3(new_n857_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1341gat));
  OAI21_X1  g661(.A(G127gat), .B1(new_n850_), .B2(new_n645_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n848_), .A2(new_n247_), .A3(new_n698_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(G1342gat));
  OAI21_X1  g664(.A(G134gat), .B1(new_n850_), .B2(new_n838_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n848_), .A2(new_n245_), .A3(new_n676_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(G1343gat));
  NAND2_X1  g667(.A1(new_n846_), .A2(new_n847_), .ZN(new_n869_));
  NOR4_X1   g668(.A1(new_n688_), .A2(new_n473_), .A3(new_n483_), .A4(new_n481_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n869_), .A2(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n654_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(new_n342_), .ZN(G1344gat));
  NOR2_X1   g672(.A1(new_n871_), .A2(new_n603_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT124), .B(G148gat), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n874_), .B(new_n875_), .ZN(G1345gat));
  NOR2_X1   g675(.A1(new_n871_), .A2(new_n645_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT61), .B(G155gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  OAI21_X1  g678(.A(G162gat), .B1(new_n871_), .B2(new_n838_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n656_), .A2(G162gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n871_), .B2(new_n881_), .ZN(G1347gat));
  NOR2_X1   g681(.A1(new_n841_), .A2(new_n835_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n491_), .A2(new_n481_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(new_n473_), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n883_), .A2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(G169gat), .B1(new_n887_), .B2(new_n654_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n888_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n888_), .A2(new_n889_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n883_), .A2(new_n886_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n892_), .A2(new_n312_), .A3(new_n529_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n890_), .A2(new_n891_), .A3(new_n893_), .ZN(G1348gat));
  AOI21_X1  g693(.A(G176gat), .B1(new_n892_), .B2(new_n602_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n478_), .B1(new_n846_), .B2(new_n847_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n603_), .A2(new_n313_), .A3(new_n884_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n895_), .B1(new_n896_), .B2(new_n897_), .ZN(G1349gat));
  NOR3_X1   g697(.A1(new_n887_), .A2(new_n316_), .A3(new_n645_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n896_), .A2(new_n698_), .A3(new_n885_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n211_), .B2(new_n900_), .ZN(G1350gat));
  NAND3_X1  g700(.A1(new_n892_), .A2(new_n210_), .A3(new_n676_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n887_), .A2(new_n838_), .ZN(new_n903_));
  INV_X1    g702(.A(G190gat), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n902_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT125), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n907_), .B(new_n902_), .C1(new_n903_), .C2(new_n904_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(G1351gat));
  NOR4_X1   g708(.A1(new_n688_), .A2(new_n473_), .A3(new_n490_), .A4(new_n482_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n869_), .A2(new_n910_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n911_), .A2(new_n654_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n280_), .A2(KEYINPUT126), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n280_), .A2(KEYINPUT126), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n912_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n915_), .B1(new_n912_), .B2(new_n914_), .ZN(G1352gat));
  NOR2_X1   g715(.A1(new_n911_), .A2(new_n603_), .ZN(new_n917_));
  XNOR2_X1  g716(.A(new_n917_), .B(new_n282_), .ZN(G1353gat));
  INV_X1    g717(.A(new_n911_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT127), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n645_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n919_), .A2(new_n920_), .A3(new_n921_), .ZN(new_n922_));
  AOI21_X1  g721(.A(new_n920_), .B1(new_n919_), .B2(new_n921_), .ZN(new_n923_));
  OAI22_X1  g722(.A1(new_n922_), .A2(new_n923_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n919_), .A2(new_n921_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(KEYINPUT127), .ZN(new_n926_));
  NOR2_X1   g725(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n919_), .A2(new_n920_), .A3(new_n921_), .ZN(new_n928_));
  NAND3_X1  g727(.A1(new_n926_), .A2(new_n927_), .A3(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n924_), .A2(new_n929_), .ZN(G1354gat));
  OR3_X1    g729(.A1(new_n911_), .A2(G218gat), .A3(new_n656_), .ZN(new_n931_));
  OAI21_X1  g730(.A(G218gat), .B1(new_n911_), .B2(new_n838_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(G1355gat));
endmodule


