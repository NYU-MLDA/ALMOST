//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n915_, new_n916_, new_n918_,
    new_n919_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n945_,
    new_n946_, new_n947_, new_n949_, new_n950_;
  NOR2_X1   g000(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n202_));
  AND2_X1   g001(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n203_));
  AND2_X1   g002(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n205_));
  OAI22_X1  g004(.A1(new_n202_), .A2(new_n203_), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT82), .ZN(new_n207_));
  XNOR2_X1  g006(.A(KEYINPUT25), .B(G183gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(KEYINPUT26), .B(G190gat), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n207_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G183gat), .A2(G190gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT23), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(G183gat), .A3(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n214_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(G169gat), .ZN(new_n218_));
  INV_X1    g017(.A(G176gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n220_), .A2(KEYINPUT24), .A3(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT24), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n217_), .A2(new_n222_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT83), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT22), .B1(new_n227_), .B2(new_n218_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT22), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(KEYINPUT83), .A3(G169gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(new_n219_), .A3(new_n230_), .ZN(new_n231_));
  OR2_X1    g030(.A1(G183gat), .A2(G190gat), .ZN(new_n232_));
  AOI22_X1  g031(.A1(new_n217_), .A2(new_n232_), .B1(G169gat), .B2(G176gat), .ZN(new_n233_));
  AOI22_X1  g032(.A1(new_n212_), .A2(new_n226_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  XNOR2_X1  g035(.A(G15gat), .B(G43gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G227gat), .A2(G233gat), .ZN(new_n238_));
  XNOR2_X1  g037(.A(new_n237_), .B(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n236_), .B(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G120gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G127gat), .A2(G134gat), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G127gat), .A2(G134gat), .ZN(new_n244_));
  NOR3_X1   g043(.A1(new_n243_), .A2(new_n244_), .A3(G113gat), .ZN(new_n245_));
  INV_X1    g044(.A(G113gat), .ZN(new_n246_));
  INV_X1    g045(.A(G127gat), .ZN(new_n247_));
  INV_X1    g046(.A(G134gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n246_), .B1(new_n249_), .B2(new_n242_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n241_), .B1(new_n245_), .B2(new_n250_), .ZN(new_n251_));
  OAI21_X1  g050(.A(G113gat), .B1(new_n243_), .B2(new_n244_), .ZN(new_n252_));
  NAND3_X1  g051(.A1(new_n249_), .A2(new_n246_), .A3(new_n242_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(G120gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n251_), .A2(new_n254_), .ZN(new_n255_));
  XOR2_X1   g054(.A(G71gat), .B(G99gat), .Z(new_n256_));
  XNOR2_X1  g055(.A(new_n256_), .B(KEYINPUT30), .ZN(new_n257_));
  XOR2_X1   g056(.A(new_n255_), .B(new_n257_), .Z(new_n258_));
  XOR2_X1   g057(.A(new_n240_), .B(new_n258_), .Z(new_n259_));
  AND2_X1   g058(.A1(G211gat), .A2(G218gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(G211gat), .A2(G218gat), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(G197gat), .ZN(new_n263_));
  AND2_X1   g062(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n264_));
  NOR2_X1   g063(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT21), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(G197gat), .B2(G204gat), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n262_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(G197gat), .B1(new_n264_), .B2(new_n265_), .ZN(new_n270_));
  INV_X1    g069(.A(G204gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(G197gat), .ZN(new_n272_));
  INV_X1    g071(.A(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n270_), .A2(new_n267_), .A3(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n270_), .A2(new_n273_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n276_), .A2(KEYINPUT21), .A3(new_n262_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n275_), .A2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(KEYINPUT94), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n218_), .A2(KEYINPUT22), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n229_), .A2(G169gat), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n279_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n229_), .A2(G169gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n218_), .A2(KEYINPUT22), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(KEYINPUT94), .ZN(new_n285_));
  AOI21_X1  g084(.A(G176gat), .B1(new_n282_), .B2(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n217_), .A2(new_n232_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n221_), .B(KEYINPUT93), .ZN(new_n289_));
  INV_X1    g088(.A(new_n289_), .ZN(new_n290_));
  NOR3_X1   g089(.A1(new_n286_), .A2(new_n288_), .A3(new_n290_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n203_), .A2(new_n202_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n205_), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT91), .ZN(new_n294_));
  NAND2_X1  g093(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT91), .B1(new_n204_), .B2(new_n205_), .ZN(new_n297_));
  AOI21_X1  g096(.A(new_n292_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT92), .ZN(new_n299_));
  AND3_X1   g098(.A1(new_n221_), .A2(new_n299_), .A3(KEYINPUT24), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n299_), .B1(new_n221_), .B2(KEYINPUT24), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n300_), .A2(new_n301_), .A3(new_n223_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n217_), .A2(new_n225_), .ZN(new_n303_));
  NOR3_X1   g102(.A1(new_n298_), .A2(new_n302_), .A3(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n278_), .B1(new_n291_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G226gat), .A2(G233gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n306_), .B(KEYINPUT19), .Z(new_n307_));
  XOR2_X1   g106(.A(new_n307_), .B(KEYINPUT90), .Z(new_n308_));
  XNOR2_X1  g107(.A(G211gat), .B(G218gat), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n270_), .B2(new_n273_), .ZN(new_n310_));
  AOI22_X1  g109(.A1(KEYINPUT21), .A2(new_n310_), .B1(new_n269_), .B2(new_n274_), .ZN(new_n311_));
  NOR2_X1   g110(.A1(new_n206_), .A2(KEYINPUT82), .ZN(new_n312_));
  AOI21_X1  g111(.A(new_n210_), .B1(new_n208_), .B2(new_n209_), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n226_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n233_), .A2(new_n231_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n311_), .A2(new_n314_), .A3(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n305_), .A2(KEYINPUT20), .A3(new_n308_), .A4(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT98), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n296_), .A2(new_n297_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(new_n208_), .ZN(new_n320_));
  OR3_X1    g119(.A1(new_n300_), .A2(new_n301_), .A3(new_n223_), .ZN(new_n321_));
  NAND4_X1  g120(.A1(new_n320_), .A2(new_n321_), .A3(new_n217_), .A4(new_n225_), .ZN(new_n322_));
  INV_X1    g121(.A(new_n285_), .ZN(new_n323_));
  AOI21_X1  g122(.A(KEYINPUT94), .B1(new_n283_), .B2(new_n284_), .ZN(new_n324_));
  OAI21_X1  g123(.A(new_n219_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(new_n287_), .A3(new_n289_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n322_), .A2(new_n311_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n315_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n217_), .A2(new_n222_), .A3(new_n225_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n329_), .B1(new_n207_), .B2(new_n211_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n278_), .B1(new_n328_), .B2(new_n330_), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n327_), .A2(new_n331_), .A3(KEYINPUT20), .ZN(new_n332_));
  INV_X1    g131(.A(new_n307_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n332_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT20), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n335_), .B1(new_n234_), .B2(new_n311_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT98), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n336_), .A2(new_n305_), .A3(new_n337_), .A4(new_n308_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n318_), .A2(new_n334_), .A3(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(KEYINPUT95), .B(KEYINPUT18), .Z(new_n340_));
  XNOR2_X1  g139(.A(G8gat), .B(G36gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n340_), .B(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G64gat), .B(G92gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n339_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n308_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n314_), .A2(new_n315_), .ZN(new_n348_));
  OAI21_X1  g147(.A(KEYINPUT20), .B1(new_n348_), .B2(new_n278_), .ZN(new_n349_));
  AOI21_X1  g148(.A(new_n311_), .B1(new_n322_), .B2(new_n326_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n347_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND4_X1  g150(.A1(new_n327_), .A2(new_n331_), .A3(KEYINPUT20), .A4(new_n307_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n351_), .A2(new_n352_), .A3(new_n344_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n346_), .A2(KEYINPUT27), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT100), .ZN(new_n355_));
  AND4_X1   g154(.A1(KEYINPUT20), .A2(new_n327_), .A3(new_n331_), .A4(new_n307_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n308_), .B1(new_n336_), .B2(new_n305_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n345_), .B1(new_n356_), .B2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n353_), .ZN(new_n359_));
  XOR2_X1   g158(.A(KEYINPUT99), .B(KEYINPUT27), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n355_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n362_));
  AOI211_X1 g161(.A(KEYINPUT100), .B(new_n360_), .C1(new_n358_), .C2(new_n353_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n354_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G225gat), .A2(G233gat), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(G141gat), .A2(G148gat), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT3), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n367_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(G141gat), .A2(G148gat), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT2), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n369_), .A2(new_n372_), .A3(new_n373_), .A4(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G155gat), .A2(G162gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n375_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n370_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n381_), .A2(new_n367_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT85), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n378_), .A2(new_n384_), .A3(KEYINPUT1), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n384_), .B1(new_n378_), .B2(KEYINPUT1), .ZN(new_n386_));
  NOR2_X1   g185(.A1(new_n385_), .A2(new_n386_), .ZN(new_n387_));
  AND2_X1   g186(.A1(G155gat), .A2(G162gat), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT1), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n376_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n383_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n255_), .B1(new_n380_), .B2(new_n391_), .ZN(new_n392_));
  OAI21_X1  g191(.A(KEYINPUT85), .B1(new_n388_), .B2(new_n389_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n378_), .A2(new_n384_), .A3(KEYINPUT1), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n390_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(new_n382_), .ZN(new_n396_));
  NAND4_X1  g195(.A1(new_n396_), .A2(new_n254_), .A3(new_n251_), .A4(new_n379_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n366_), .B1(new_n392_), .B2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n392_), .A2(KEYINPUT4), .A3(new_n397_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(KEYINPUT96), .ZN(new_n400_));
  OR2_X1    g199(.A1(new_n392_), .A2(KEYINPUT4), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT96), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n392_), .A2(new_n402_), .A3(KEYINPUT4), .A4(new_n397_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n400_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n398_), .B1(new_n404_), .B2(new_n366_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(G85gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT0), .ZN(new_n408_));
  OR2_X1    g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n408_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n409_), .A2(G57gat), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(G57gat), .B1(new_n409_), .B2(new_n410_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n411_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n405_), .A2(new_n414_), .ZN(new_n415_));
  AOI211_X1 g214(.A(new_n398_), .B(new_n413_), .C1(new_n404_), .C2(new_n366_), .ZN(new_n416_));
  NOR2_X1   g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n396_), .A2(new_n379_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT29), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n421_));
  INV_X1    g220(.A(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n419_), .A2(new_n420_), .A3(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n421_), .B1(new_n418_), .B2(KEYINPUT29), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G22gat), .B(G50gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(new_n425_), .B(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G228gat), .A2(G233gat), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n278_), .B(new_n429_), .C1(new_n419_), .C2(new_n420_), .ZN(new_n430_));
  AOI21_X1  g229(.A(new_n420_), .B1(new_n396_), .B2(new_n379_), .ZN(new_n431_));
  OAI211_X1 g230(.A(G228gat), .B(G233gat), .C1(new_n431_), .C2(new_n311_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G78gat), .B(G106gat), .ZN(new_n433_));
  XOR2_X1   g232(.A(new_n433_), .B(KEYINPUT88), .Z(new_n434_));
  INV_X1    g233(.A(new_n434_), .ZN(new_n435_));
  NAND4_X1  g234(.A1(new_n430_), .A2(new_n432_), .A3(KEYINPUT89), .A4(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n430_), .A2(new_n432_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n437_), .A2(new_n434_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT89), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n437_), .B2(new_n433_), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n428_), .B(new_n436_), .C1(new_n438_), .C2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n425_), .B(new_n426_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n435_), .B1(new_n430_), .B2(new_n432_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n442_), .B1(new_n438_), .B2(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n441_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n417_), .A2(new_n445_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n364_), .A2(new_n446_), .ZN(new_n447_));
  NAND4_X1  g246(.A1(new_n400_), .A2(new_n365_), .A3(new_n401_), .A4(new_n403_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n392_), .A2(new_n366_), .A3(new_n397_), .ZN(new_n449_));
  AND3_X1   g248(.A1(new_n448_), .A2(new_n414_), .A3(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n450_), .A2(new_n359_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n404_), .A2(new_n366_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n398_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n454_), .A2(KEYINPUT33), .A3(new_n413_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT33), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n456_), .B1(new_n405_), .B2(new_n414_), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n451_), .A2(new_n455_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n344_), .A2(KEYINPUT32), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n351_), .A2(new_n352_), .A3(new_n459_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT97), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n339_), .A2(new_n460_), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  OR2_X1    g262(.A1(new_n461_), .A2(new_n462_), .ZN(new_n464_));
  OAI211_X1 g263(.A(new_n463_), .B(new_n464_), .C1(new_n415_), .C2(new_n416_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n445_), .B1(new_n458_), .B2(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n259_), .B1(new_n447_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(KEYINPUT101), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT101), .ZN(new_n469_));
  OAI211_X1 g268(.A(new_n469_), .B(new_n259_), .C1(new_n447_), .C2(new_n466_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n468_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT102), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n364_), .A2(new_n472_), .ZN(new_n473_));
  OAI211_X1 g272(.A(KEYINPUT102), .B(new_n354_), .C1(new_n362_), .C2(new_n363_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n445_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n473_), .A2(new_n474_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT103), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n259_), .ZN(new_n479_));
  NAND4_X1  g278(.A1(new_n473_), .A2(KEYINPUT103), .A3(new_n474_), .A4(new_n475_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n478_), .A2(new_n417_), .A3(new_n479_), .A4(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n471_), .A2(new_n481_), .ZN(new_n482_));
  XNOR2_X1  g281(.A(G29gat), .B(G36gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n483_), .B(KEYINPUT74), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(G43gat), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT74), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n483_), .B(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(G43gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n487_), .A2(new_n488_), .ZN(new_n489_));
  AOI21_X1  g288(.A(G50gat), .B1(new_n485_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n485_), .A2(new_n489_), .A3(G50gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n491_), .A2(KEYINPUT15), .A3(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT15), .ZN(new_n494_));
  INV_X1    g293(.A(new_n492_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n494_), .B1(new_n495_), .B2(new_n490_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n493_), .A2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n498_));
  INV_X1    g297(.A(G85gat), .ZN(new_n499_));
  INV_X1    g298(.A(G92gat), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT64), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT9), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT9), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT64), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n501_), .A2(new_n503_), .A3(new_n505_), .ZN(new_n506_));
  AND2_X1   g305(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n507_));
  NOR2_X1   g306(.A1(KEYINPUT65), .A2(G92gat), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n507_), .A2(new_n508_), .A3(new_n499_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n498_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT66), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G99gat), .A2(G106gat), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT6), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n512_), .B(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  XOR2_X1   g314(.A(KEYINPUT10), .B(G99gat), .Z(new_n516_));
  INV_X1    g315(.A(G106gat), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND4_X1  g317(.A1(new_n510_), .A2(new_n511_), .A3(new_n515_), .A4(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n510_), .A2(new_n515_), .A3(new_n518_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT66), .ZN(new_n521_));
  XOR2_X1   g320(.A(G85gat), .B(G92gat), .Z(new_n522_));
  OR3_X1    g321(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n523_));
  OAI21_X1  g322(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n522_), .B1(new_n514_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n526_), .A2(KEYINPUT8), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT8), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n528_), .B(new_n522_), .C1(new_n514_), .C2(new_n525_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n527_), .A2(KEYINPUT70), .A3(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT70), .B1(new_n527_), .B2(new_n529_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n519_), .B(new_n521_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT75), .B1(new_n497_), .B2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G232gat), .A2(G233gat), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT72), .Z(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT34), .ZN(new_n536_));
  OR2_X1    g335(.A1(new_n536_), .A2(KEYINPUT35), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n527_), .A2(new_n529_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n521_), .A2(new_n538_), .A3(new_n519_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n539_), .A2(KEYINPUT67), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT67), .ZN(new_n541_));
  NAND4_X1  g340(.A1(new_n521_), .A2(new_n538_), .A3(new_n541_), .A4(new_n519_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n540_), .A2(new_n542_), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(new_n492_), .A3(new_n491_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n533_), .A2(new_n537_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n536_), .A2(KEYINPUT35), .ZN(new_n546_));
  XOR2_X1   g345(.A(new_n546_), .B(KEYINPUT73), .Z(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n545_), .A2(new_n548_), .ZN(new_n549_));
  NAND4_X1  g348(.A1(new_n533_), .A2(new_n544_), .A3(new_n537_), .A4(new_n547_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G190gat), .B(G218gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n552_), .B(new_n248_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(G162gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n554_), .B(KEYINPUT36), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n551_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT36), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n554_), .A2(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n559_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n557_), .A2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n482_), .A2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT106), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT13), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G230gat), .A2(G233gat), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G57gat), .B(G64gat), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT11), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G71gat), .B(G78gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n570_), .B(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n569_), .A2(KEYINPUT11), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n575_), .B1(new_n540_), .B2(new_n542_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT68), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n540_), .A2(new_n575_), .A3(new_n542_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT69), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n568_), .B1(new_n577_), .B2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT12), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n576_), .B1(new_n581_), .B2(new_n578_), .ZN(new_n582_));
  NAND3_X1  g381(.A1(new_n532_), .A2(KEYINPUT12), .A3(new_n575_), .ZN(new_n583_));
  NAND3_X1  g382(.A1(new_n582_), .A2(new_n567_), .A3(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G120gat), .B(G148gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT5), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(G176gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(new_n271_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n580_), .A2(new_n584_), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n589_), .B1(new_n580_), .B2(new_n584_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n566_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(KEYINPUT13), .A3(new_n590_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n593_), .A2(new_n595_), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G15gat), .B(G22gat), .ZN(new_n597_));
  INV_X1    g396(.A(G1gat), .ZN(new_n598_));
  INV_X1    g397(.A(G8gat), .ZN(new_n599_));
  OAI21_X1  g398(.A(KEYINPUT14), .B1(new_n598_), .B2(new_n599_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n597_), .A2(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(G1gat), .B(G8gat), .ZN(new_n602_));
  XOR2_X1   g401(.A(new_n601_), .B(new_n602_), .Z(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n497_), .A2(new_n604_), .ZN(new_n605_));
  NOR3_X1   g404(.A1(new_n495_), .A2(new_n604_), .A3(new_n490_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G229gat), .A2(G233gat), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n605_), .A2(new_n607_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n608_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n603_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n610_), .B1(new_n611_), .B2(new_n606_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT80), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT80), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n614_), .B(new_n610_), .C1(new_n611_), .C2(new_n606_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n609_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(G113gat), .B(G141gat), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(KEYINPUT81), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n618_), .B(new_n218_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(new_n263_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n616_), .B(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n596_), .A2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(G231gat), .A2(G233gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n625_), .B(KEYINPUT77), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n603_), .B(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(new_n575_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(G127gat), .B(G155gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n629_), .B(KEYINPUT16), .ZN(new_n630_));
  INV_X1    g429(.A(G183gat), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  XNOR2_X1  g431(.A(new_n632_), .B(G211gat), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT17), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n628_), .A2(new_n635_), .ZN(new_n636_));
  XNOR2_X1  g435(.A(new_n636_), .B(KEYINPUT78), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n633_), .A2(new_n634_), .ZN(new_n638_));
  OR3_X1    g437(.A1(new_n628_), .A2(new_n638_), .A3(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT79), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n482_), .A2(KEYINPUT106), .A3(new_n562_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n565_), .A2(new_n624_), .A3(new_n642_), .A4(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G1gat), .B1(new_n644_), .B2(new_n417_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n557_), .A2(KEYINPUT37), .A3(new_n560_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT37), .ZN(new_n647_));
  INV_X1    g446(.A(new_n560_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n556_), .A2(KEYINPUT76), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n556_), .A2(KEYINPUT76), .ZN(new_n650_));
  NAND4_X1  g449(.A1(new_n549_), .A2(new_n550_), .A3(new_n649_), .A4(new_n650_), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n647_), .B1(new_n648_), .B2(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n646_), .A2(new_n652_), .ZN(new_n653_));
  AOI211_X1 g452(.A(new_n641_), .B(new_n653_), .C1(new_n471_), .C2(new_n481_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n596_), .B(KEYINPUT71), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n622_), .A3(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT104), .ZN(new_n657_));
  INV_X1    g456(.A(new_n417_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n657_), .A2(new_n598_), .A3(new_n658_), .ZN(new_n659_));
  OR2_X1    g458(.A1(new_n659_), .A2(KEYINPUT105), .ZN(new_n660_));
  INV_X1    g459(.A(KEYINPUT38), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(KEYINPUT105), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n660_), .A2(new_n661_), .A3(new_n662_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n661_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n645_), .B1(new_n663_), .B2(new_n664_), .ZN(G1324gat));
  NAND2_X1  g464(.A1(new_n473_), .A2(new_n474_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n657_), .A2(new_n599_), .A3(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n666_), .ZN(new_n668_));
  OAI21_X1  g467(.A(G8gat), .B1(new_n644_), .B2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT107), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT39), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT107), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n672_), .B(G8gat), .C1(new_n644_), .C2(new_n668_), .ZN(new_n673_));
  AND3_X1   g472(.A1(new_n670_), .A2(new_n671_), .A3(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n671_), .B1(new_n670_), .B2(new_n673_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n667_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT40), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n676_), .B(new_n677_), .ZN(G1325gat));
  OAI21_X1  g477(.A(G15gat), .B1(new_n644_), .B2(new_n259_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT41), .Z(new_n680_));
  INV_X1    g479(.A(G15gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n657_), .A2(new_n681_), .A3(new_n479_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(G1326gat));
  OAI21_X1  g482(.A(G22gat), .B1(new_n644_), .B2(new_n475_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT42), .ZN(new_n685_));
  INV_X1    g484(.A(G22gat), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n657_), .A2(new_n686_), .A3(new_n445_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n685_), .A2(new_n687_), .ZN(G1327gat));
  NOR2_X1   g487(.A1(new_n642_), .A2(new_n562_), .ZN(new_n689_));
  AND3_X1   g488(.A1(new_n482_), .A2(new_n624_), .A3(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(G29gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n690_), .A2(new_n691_), .A3(new_n658_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n482_), .A2(new_n653_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n693_), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n648_), .A2(new_n651_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(KEYINPUT37), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n648_), .B(new_n647_), .C1(new_n551_), .C2(new_n556_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n698_), .B1(new_n471_), .B2(new_n481_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT43), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n699_), .A2(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT108), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(new_n699_), .B2(new_n700_), .ZN(new_n703_));
  NAND3_X1  g502(.A1(new_n694_), .A2(new_n701_), .A3(new_n703_), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n704_), .A2(new_n624_), .A3(new_n641_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT109), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n705_), .A2(new_n706_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n707_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n704_), .A2(new_n624_), .A3(new_n641_), .A4(new_n709_), .ZN(new_n710_));
  AND3_X1   g509(.A1(new_n708_), .A2(new_n658_), .A3(new_n710_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n692_), .B1(new_n711_), .B2(new_n691_), .ZN(G1328gat));
  NAND3_X1  g511(.A1(new_n708_), .A2(new_n666_), .A3(new_n710_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(G36gat), .ZN(new_n714_));
  INV_X1    g513(.A(G36gat), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n690_), .A2(new_n666_), .A3(new_n715_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(new_n716_), .B(KEYINPUT45), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n714_), .A2(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT46), .B1(new_n718_), .B2(KEYINPUT110), .ZN(new_n719_));
  INV_X1    g518(.A(new_n717_), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n720_), .B1(new_n713_), .B2(G36gat), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT46), .ZN(new_n723_));
  NOR3_X1   g522(.A1(new_n721_), .A2(new_n722_), .A3(new_n723_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n719_), .A2(new_n724_), .ZN(G1329gat));
  NAND3_X1  g524(.A1(new_n690_), .A2(new_n488_), .A3(new_n479_), .ZN(new_n726_));
  AND3_X1   g525(.A1(new_n708_), .A2(new_n479_), .A3(new_n710_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(new_n488_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT47), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n728_), .B(new_n729_), .ZN(G1330gat));
  INV_X1    g529(.A(G50gat), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n690_), .A2(new_n731_), .A3(new_n445_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n708_), .A2(new_n445_), .A3(new_n710_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n732_), .B1(new_n733_), .B2(new_n731_), .ZN(G1331gat));
  AND3_X1   g533(.A1(new_n654_), .A2(new_n623_), .A3(new_n596_), .ZN(new_n735_));
  AOI21_X1  g534(.A(G57gat), .B1(new_n735_), .B2(new_n658_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n565_), .A2(new_n642_), .A3(new_n643_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n655_), .A2(new_n622_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n739_), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n658_), .A2(G57gat), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n736_), .B1(new_n740_), .B2(new_n741_), .ZN(G1332gat));
  OAI21_X1  g541(.A(G64gat), .B1(new_n739_), .B2(new_n668_), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT48), .ZN(new_n744_));
  INV_X1    g543(.A(G64gat), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n735_), .A2(new_n745_), .A3(new_n666_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n739_), .B2(new_n259_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT49), .ZN(new_n749_));
  INV_X1    g548(.A(G71gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n735_), .A2(new_n750_), .A3(new_n479_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n749_), .A2(new_n751_), .ZN(G1334gat));
  OAI21_X1  g551(.A(G78gat), .B1(new_n739_), .B2(new_n475_), .ZN(new_n753_));
  XNOR2_X1  g552(.A(new_n753_), .B(KEYINPUT50), .ZN(new_n754_));
  INV_X1    g553(.A(G78gat), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n735_), .A2(new_n755_), .A3(new_n445_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n754_), .A2(new_n756_), .ZN(G1335gat));
  AND3_X1   g556(.A1(new_n738_), .A2(new_n482_), .A3(new_n689_), .ZN(new_n758_));
  AOI21_X1  g557(.A(G85gat), .B1(new_n758_), .B2(new_n658_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n596_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n760_), .A2(new_n622_), .A3(new_n642_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n704_), .A2(new_n761_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT111), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(KEYINPUT111), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n417_), .B1(new_n763_), .B2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n759_), .B1(new_n765_), .B2(G85gat), .ZN(G1336gat));
  NAND2_X1  g565(.A1(new_n763_), .A2(new_n764_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n668_), .A2(new_n508_), .A3(new_n507_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT112), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n758_), .A2(new_n666_), .ZN(new_n770_));
  AOI22_X1  g569(.A1(new_n767_), .A2(new_n769_), .B1(new_n500_), .B2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT113), .ZN(G1337gat));
  NAND3_X1  g571(.A1(new_n758_), .A2(new_n516_), .A3(new_n479_), .ZN(new_n773_));
  XNOR2_X1  g572(.A(new_n773_), .B(KEYINPUT114), .ZN(new_n774_));
  OAI21_X1  g573(.A(G99gat), .B1(new_n762_), .B2(new_n259_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT115), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777_));
  OAI211_X1 g576(.A(new_n774_), .B(new_n775_), .C1(new_n776_), .C2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n777_), .ZN(new_n779_));
  XNOR2_X1  g578(.A(new_n778_), .B(new_n779_), .ZN(G1338gat));
  XNOR2_X1  g579(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n704_), .A2(new_n445_), .A3(new_n761_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT116), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n782_), .A2(new_n783_), .A3(G106gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n782_), .B2(G106gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(KEYINPUT52), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n782_), .A2(G106gat), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(KEYINPUT116), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n782_), .A2(new_n783_), .A3(G106gat), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n788_), .A2(new_n789_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n786_), .A2(new_n791_), .ZN(new_n792_));
  AND3_X1   g591(.A1(new_n758_), .A2(new_n517_), .A3(new_n445_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n781_), .B1(new_n792_), .B2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n781_), .ZN(new_n796_));
  AOI211_X1 g595(.A(new_n796_), .B(new_n793_), .C1(new_n786_), .C2(new_n791_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n795_), .A2(new_n797_), .ZN(G1339gat));
  INV_X1    g597(.A(KEYINPUT54), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n653_), .A2(new_n622_), .A3(new_n641_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n799_), .B1(new_n800_), .B2(new_n760_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n698_), .A2(new_n642_), .A3(new_n623_), .ZN(new_n802_));
  NOR3_X1   g601(.A1(new_n802_), .A2(new_n596_), .A3(KEYINPUT54), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n616_), .A2(new_n621_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n608_), .B1(new_n611_), .B2(new_n606_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n605_), .A2(new_n610_), .A3(new_n607_), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n807_), .A2(new_n621_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n805_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n567_), .B1(new_n582_), .B2(new_n583_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT55), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n584_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n578_), .A2(new_n581_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n543_), .A2(new_n574_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n813_), .A2(new_n583_), .A3(new_n814_), .ZN(new_n815_));
  NOR3_X1   g614(.A1(new_n815_), .A2(new_n811_), .A3(new_n568_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n812_), .A2(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT56), .B1(new_n818_), .B2(new_n588_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT56), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n820_), .B(new_n589_), .C1(new_n812_), .C2(new_n817_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n590_), .B(new_n809_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT58), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n698_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  OAI21_X1  g623(.A(KEYINPUT119), .B1(new_n822_), .B2(new_n823_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n811_), .B1(new_n815_), .B2(new_n568_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n815_), .A2(new_n568_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n826_), .A2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n588_), .B1(new_n828_), .B2(new_n816_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n820_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n818_), .A2(KEYINPUT56), .A3(new_n588_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n591_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n832_), .A2(new_n833_), .A3(KEYINPUT58), .A4(new_n809_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n824_), .A2(new_n825_), .A3(new_n834_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n622_), .A2(new_n590_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n836_), .B1(new_n819_), .B2(new_n821_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n594_), .A2(new_n590_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(new_n809_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n561_), .B1(new_n837_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT118), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT57), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT57), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n830_), .A2(new_n831_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n844_), .A2(new_n836_), .B1(new_n838_), .B2(new_n809_), .ZN(new_n845_));
  OAI211_X1 g644(.A(KEYINPUT118), .B(new_n843_), .C1(new_n845_), .C2(new_n561_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n835_), .A2(new_n842_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n804_), .B1(new_n847_), .B2(new_n641_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n417_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n478_), .A2(new_n480_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(new_n479_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n849_), .A2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(G113gat), .B1(new_n854_), .B2(new_n622_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n856_));
  AND3_X1   g655(.A1(new_n849_), .A2(new_n852_), .A3(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT120), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n860_), .B1(new_n849_), .B2(new_n852_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n623_), .B1(new_n858_), .B2(new_n862_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n855_), .B1(new_n863_), .B2(G113gat), .ZN(G1340gat));
  AOI21_X1  g663(.A(KEYINPUT60), .B1(new_n596_), .B2(new_n241_), .ZN(new_n865_));
  OR3_X1    g664(.A1(new_n853_), .A2(KEYINPUT60), .A3(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n655_), .ZN(new_n867_));
  OAI221_X1 g666(.A(new_n867_), .B1(new_n853_), .B2(new_n865_), .C1(new_n857_), .C2(new_n861_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n866_), .B1(new_n869_), .B2(new_n241_), .ZN(G1341gat));
  AOI21_X1  g669(.A(G127gat), .B1(new_n854_), .B2(new_n642_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n641_), .B1(new_n858_), .B2(new_n862_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n871_), .B1(new_n872_), .B2(G127gat), .ZN(G1342gat));
  AOI21_X1  g672(.A(G134gat), .B1(new_n854_), .B2(new_n561_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n698_), .B1(new_n858_), .B2(new_n862_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(G134gat), .ZN(G1343gat));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n479_), .A2(new_n475_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NOR2_X1   g678(.A1(new_n879_), .A2(new_n666_), .ZN(new_n880_));
  AND3_X1   g679(.A1(new_n849_), .A2(new_n877_), .A3(new_n880_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n877_), .B1(new_n849_), .B2(new_n880_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n622_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(KEYINPUT122), .B(G141gat), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n883_), .B(new_n884_), .ZN(G1344gat));
  OAI21_X1  g684(.A(new_n867_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g686(.A(KEYINPUT61), .B(G155gat), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(KEYINPUT123), .ZN(new_n889_));
  OR2_X1    g688(.A1(new_n881_), .A2(new_n882_), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n889_), .B1(new_n890_), .B2(new_n642_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n642_), .B(new_n889_), .C1(new_n881_), .C2(new_n882_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1346gat));
  AOI21_X1  g693(.A(G162gat), .B1(new_n890_), .B2(new_n561_), .ZN(new_n895_));
  OAI211_X1 g694(.A(G162gat), .B(new_n653_), .C1(new_n881_), .C2(new_n882_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n895_), .A2(new_n897_), .ZN(G1347gat));
  XOR2_X1   g697(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n848_), .A2(new_n445_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n668_), .A2(new_n658_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(new_n479_), .ZN(new_n903_));
  XOR2_X1   g702(.A(new_n903_), .B(KEYINPUT124), .Z(new_n904_));
  NAND2_X1  g703(.A1(new_n901_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n623_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n900_), .B1(new_n906_), .B2(new_n218_), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n908_));
  OAI211_X1 g707(.A(G169gat), .B(new_n899_), .C1(new_n905_), .C2(new_n623_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(G1348gat));
  NOR3_X1   g709(.A1(new_n905_), .A2(new_n219_), .A3(new_n655_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n905_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n596_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n911_), .B1(new_n219_), .B2(new_n913_), .ZN(G1349gat));
  NOR2_X1   g713(.A1(new_n905_), .A2(new_n641_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(new_n208_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n916_), .B1(new_n915_), .B2(new_n631_), .ZN(G1350gat));
  OAI21_X1  g716(.A(G190gat), .B1(new_n905_), .B2(new_n698_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n561_), .A2(new_n319_), .ZN(new_n919_));
  OAI21_X1  g718(.A(new_n918_), .B1(new_n905_), .B2(new_n919_), .ZN(G1351gat));
  NAND2_X1  g719(.A1(new_n847_), .A2(new_n641_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n804_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NAND3_X1  g722(.A1(new_n923_), .A2(new_n878_), .A3(new_n902_), .ZN(new_n924_));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n879_), .B1(new_n921_), .B2(new_n922_), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n927_), .A2(KEYINPUT126), .A3(new_n902_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(new_n622_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(G197gat), .ZN(G1352gat));
  INV_X1    g730(.A(new_n265_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(KEYINPUT87), .A2(G204gat), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n932_), .A2(new_n933_), .ZN(new_n934_));
  AOI21_X1  g733(.A(KEYINPUT126), .B1(new_n927_), .B2(new_n902_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n902_), .ZN(new_n936_));
  NOR4_X1   g735(.A1(new_n848_), .A2(new_n925_), .A3(new_n879_), .A4(new_n936_), .ZN(new_n937_));
  OAI211_X1 g736(.A(new_n934_), .B(new_n867_), .C1(new_n935_), .C2(new_n937_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n655_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n938_), .B1(new_n939_), .B2(new_n271_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n940_), .A2(KEYINPUT127), .ZN(new_n941_));
  INV_X1    g740(.A(KEYINPUT127), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n938_), .A2(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n941_), .A2(new_n943_), .ZN(G1353gat));
  AOI21_X1  g743(.A(new_n641_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n945_));
  NOR3_X1   g744(.A1(new_n945_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n946_));
  XOR2_X1   g745(.A(KEYINPUT63), .B(G211gat), .Z(new_n947_));
  AOI21_X1  g746(.A(new_n946_), .B1(new_n945_), .B2(new_n947_), .ZN(G1354gat));
  AOI21_X1  g747(.A(G218gat), .B1(new_n929_), .B2(new_n561_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n698_), .B1(new_n926_), .B2(new_n928_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(G218gat), .B2(new_n950_), .ZN(G1355gat));
endmodule


