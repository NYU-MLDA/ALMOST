//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n649_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n713_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n726_, new_n727_,
    new_n728_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n874_, new_n875_,
    new_n877_, new_n879_, new_n880_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n907_, new_n908_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT0), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n204_), .B(G57gat), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G127gat), .B(G134gat), .ZN(new_n207_));
  INV_X1    g006(.A(G113gat), .ZN(new_n208_));
  XNOR2_X1  g007(.A(new_n207_), .B(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(G120gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT4), .ZN(new_n211_));
  OR2_X1    g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NOR2_X1   g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  NOR2_X1   g013(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n215_));
  XNOR2_X1  g014(.A(new_n214_), .B(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT2), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  NAND3_X1  g018(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n220_));
  NAND2_X1  g019(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n222_));
  OAI211_X1 g021(.A(new_n212_), .B(new_n213_), .C1(new_n216_), .C2(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n213_), .A2(KEYINPUT1), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n213_), .A2(KEYINPUT1), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n212_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(new_n214_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n217_), .A3(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n223_), .A2(new_n228_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n210_), .A2(new_n211_), .A3(new_n229_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n210_), .B(new_n229_), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n230_), .B1(new_n231_), .B2(new_n211_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(G225gat), .A2(G233gat), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n231_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n235_), .A2(new_n233_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n206_), .B1(new_n234_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n234_), .A2(new_n206_), .A3(new_n236_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G228gat), .A2(G233gat), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT91), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n242_), .B1(new_n229_), .B2(KEYINPUT29), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT29), .ZN(new_n244_));
  AOI211_X1 g043(.A(KEYINPUT91), .B(new_n244_), .C1(new_n223_), .C2(new_n228_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n241_), .B1(new_n243_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(G197gat), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n247_), .A2(KEYINPUT92), .A3(G204gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(G204gat), .ZN(new_n249_));
  INV_X1    g048(.A(G204gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(G197gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n249_), .A2(new_n251_), .ZN(new_n252_));
  OAI211_X1 g051(.A(KEYINPUT21), .B(new_n248_), .C1(new_n252_), .C2(KEYINPUT92), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT93), .ZN(new_n254_));
  XOR2_X1   g053(.A(G211gat), .B(G218gat), .Z(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n252_), .A2(KEYINPUT21), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n254_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(KEYINPUT21), .A3(new_n252_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT94), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n258_), .A2(KEYINPUT94), .A3(new_n259_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n246_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G22gat), .B(G50gat), .ZN(new_n266_));
  INV_X1    g065(.A(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n229_), .A2(KEYINPUT29), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n241_), .B1(new_n260_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n265_), .A2(new_n267_), .A3(new_n270_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n266_), .B1(new_n264_), .B2(new_n269_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(new_n229_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G78gat), .B(G106gat), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n244_), .A3(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n275_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n277_), .B1(new_n229_), .B2(KEYINPUT29), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  XOR2_X1   g078(.A(KEYINPUT90), .B(KEYINPUT28), .Z(new_n280_));
  AND2_X1   g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NOR2_X1   g080(.A1(new_n279_), .A2(new_n280_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n273_), .A2(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n271_), .A2(new_n272_), .A3(new_n283_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n210_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT88), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT23), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n289_), .A2(G183gat), .A3(G190gat), .ZN(new_n290_));
  INV_X1    g089(.A(G183gat), .ZN(new_n291_));
  INV_X1    g090(.A(G190gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(KEYINPUT23), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  AND2_X1   g092(.A1(new_n293_), .A2(KEYINPUT85), .ZN(new_n294_));
  NOR2_X1   g093(.A1(new_n293_), .A2(KEYINPUT85), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n290_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT24), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299_));
  MUX2_X1   g098(.A(new_n298_), .B(KEYINPUT24), .S(new_n299_), .Z(new_n300_));
  NOR2_X1   g099(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(KEYINPUT84), .B(G190gat), .Z(new_n302_));
  AOI21_X1  g101(.A(new_n301_), .B1(new_n302_), .B2(KEYINPUT26), .ZN(new_n303_));
  XOR2_X1   g102(.A(KEYINPUT25), .B(G183gat), .Z(new_n304_));
  OAI211_X1 g103(.A(new_n296_), .B(new_n300_), .C1(new_n303_), .C2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(G176gat), .ZN(new_n306_));
  INV_X1    g105(.A(G169gat), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT22), .B1(new_n307_), .B2(KEYINPUT86), .ZN(new_n308_));
  OR2_X1    g107(.A1(new_n307_), .A2(KEYINPUT22), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n306_), .B(new_n308_), .C1(new_n309_), .C2(KEYINPUT86), .ZN(new_n310_));
  INV_X1    g109(.A(new_n293_), .ZN(new_n311_));
  OR2_X1    g110(.A1(new_n290_), .A2(KEYINPUT87), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n290_), .A2(KEYINPUT87), .ZN(new_n313_));
  AOI21_X1  g112(.A(new_n311_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n302_), .A2(G183gat), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n297_), .B(new_n310_), .C1(new_n314_), .C2(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT30), .ZN(new_n317_));
  AND3_X1   g116(.A1(new_n305_), .A2(new_n316_), .A3(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n317_), .B1(new_n305_), .B2(new_n316_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n288_), .B1(new_n318_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT31), .ZN(new_n321_));
  XOR2_X1   g120(.A(G15gat), .B(G43gat), .Z(new_n322_));
  XNOR2_X1  g121(.A(G71gat), .B(G99gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G227gat), .A2(G233gat), .ZN(new_n325_));
  XOR2_X1   g124(.A(new_n324_), .B(new_n325_), .Z(new_n326_));
  NAND3_X1  g125(.A1(new_n320_), .A2(new_n321_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(new_n321_), .B1(new_n320_), .B2(new_n326_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n287_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n320_), .A2(new_n326_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(KEYINPUT31), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(new_n210_), .A3(new_n327_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n318_), .A2(new_n319_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(new_n288_), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n330_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n335_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n285_), .B(new_n286_), .C1(new_n336_), .C2(new_n337_), .ZN(new_n338_));
  NOR3_X1   g137(.A1(new_n328_), .A2(new_n329_), .A3(new_n287_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n210_), .B1(new_n332_), .B2(new_n327_), .ZN(new_n340_));
  OAI22_X1  g139(.A1(new_n339_), .A2(new_n340_), .B1(new_n288_), .B2(new_n334_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n330_), .A2(new_n333_), .A3(new_n335_), .ZN(new_n342_));
  AND3_X1   g141(.A1(new_n271_), .A2(new_n272_), .A3(new_n283_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n283_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n341_), .B(new_n342_), .C1(new_n343_), .C2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n240_), .B1(new_n338_), .B2(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n347_), .B(KEYINPUT95), .Z(new_n348_));
  XOR2_X1   g147(.A(new_n348_), .B(KEYINPUT19), .Z(new_n349_));
  INV_X1    g148(.A(KEYINPUT20), .ZN(new_n350_));
  INV_X1    g149(.A(new_n304_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT26), .B(G190gat), .ZN(new_n352_));
  AND2_X1   g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n300_), .ZN(new_n354_));
  OR3_X1    g153(.A1(new_n353_), .A2(new_n354_), .A3(new_n314_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n291_), .A2(new_n292_), .ZN(new_n356_));
  AOI22_X1  g155(.A1(new_n296_), .A2(new_n356_), .B1(G169gat), .B2(G176gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(KEYINPUT22), .B(G169gat), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(new_n306_), .ZN(new_n359_));
  AND3_X1   g158(.A1(new_n357_), .A2(KEYINPUT96), .A3(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(KEYINPUT96), .B1(new_n357_), .B2(new_n359_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n355_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n350_), .B1(new_n362_), .B2(new_n260_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n305_), .A2(new_n316_), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n262_), .A2(new_n263_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n349_), .B1(new_n363_), .B2(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT18), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G64gat), .ZN(new_n371_));
  INV_X1    g170(.A(G92gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT97), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n262_), .A2(new_n263_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n374_), .B1(new_n375_), .B2(new_n364_), .ZN(new_n376_));
  AOI211_X1 g175(.A(KEYINPUT97), .B(new_n365_), .C1(new_n262_), .C2(new_n263_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n376_), .A2(new_n377_), .ZN(new_n378_));
  OAI211_X1 g177(.A(KEYINPUT20), .B(new_n349_), .C1(new_n362_), .C2(new_n260_), .ZN(new_n379_));
  OAI211_X1 g178(.A(new_n368_), .B(new_n373_), .C1(new_n378_), .C2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n373_), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n258_), .A2(KEYINPUT94), .A3(new_n259_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT94), .B1(new_n258_), .B2(new_n259_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n364_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(KEYINPUT97), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n375_), .A2(new_n374_), .A3(new_n364_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n379_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n381_), .B1(new_n387_), .B2(new_n367_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n380_), .A2(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT27), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT100), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n363_), .A2(new_n349_), .A3(new_n366_), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  XOR2_X1   g193(.A(KEYINPUT98), .B(KEYINPUT20), .Z(new_n395_));
  INV_X1    g194(.A(new_n260_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n357_), .A2(new_n359_), .ZN(new_n397_));
  AND2_X1   g196(.A1(new_n397_), .A2(new_n355_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n395_), .B1(new_n396_), .B2(new_n398_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n399_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n349_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n394_), .B1(new_n400_), .B2(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(new_n402_), .A2(new_n373_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n380_), .A2(KEYINPUT27), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n392_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n399_), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n406_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n393_), .B1(new_n407_), .B2(new_n349_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n408_), .A2(new_n381_), .ZN(new_n409_));
  NAND4_X1  g208(.A1(new_n409_), .A2(KEYINPUT100), .A3(KEYINPUT27), .A4(new_n380_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n346_), .A2(new_n391_), .A3(new_n405_), .A4(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n233_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n235_), .A2(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n413_), .B1(new_n232_), .B2(new_n412_), .ZN(new_n414_));
  OAI21_X1  g213(.A(KEYINPUT33), .B1(new_n414_), .B2(new_n206_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n415_), .A2(new_n239_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n234_), .A2(KEYINPUT33), .A3(new_n206_), .A4(new_n236_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n416_), .A2(new_n380_), .A3(new_n388_), .A4(new_n417_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n239_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n420_), .A2(new_n237_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n373_), .A2(KEYINPUT32), .ZN(new_n422_));
  OAI21_X1  g221(.A(KEYINPUT99), .B1(new_n402_), .B2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT99), .ZN(new_n424_));
  INV_X1    g223(.A(new_n422_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n408_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n421_), .B1(new_n423_), .B2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n387_), .A2(new_n367_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n428_), .A2(new_n422_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n419_), .B1(new_n427_), .B2(new_n429_), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n336_), .A2(new_n337_), .ZN(new_n431_));
  NOR2_X1   g230(.A1(new_n343_), .A2(new_n344_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  OAI21_X1  g232(.A(new_n411_), .B1(new_n430_), .B2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(KEYINPUT78), .B(G15gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(G22gat), .ZN(new_n436_));
  INV_X1    g235(.A(G1gat), .ZN(new_n437_));
  INV_X1    g236(.A(G8gat), .ZN(new_n438_));
  OAI21_X1  g237(.A(KEYINPUT14), .B1(new_n437_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n436_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT79), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XOR2_X1   g241(.A(G1gat), .B(G8gat), .Z(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n440_), .B(KEYINPUT79), .ZN(new_n445_));
  INV_X1    g244(.A(new_n443_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G29gat), .B(G36gat), .ZN(new_n449_));
  INV_X1    g248(.A(G43gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(G50gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT15), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n448_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(G229gat), .A2(G233gat), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n444_), .A2(new_n447_), .A3(new_n453_), .ZN(new_n459_));
  INV_X1    g258(.A(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n457_), .A2(new_n458_), .A3(new_n460_), .ZN(new_n461_));
  AND2_X1   g260(.A1(new_n444_), .A2(new_n447_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n462_), .A2(new_n453_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(KEYINPUT82), .A3(new_n460_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n458_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT82), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n462_), .A2(new_n453_), .ZN(new_n467_));
  OAI21_X1  g266(.A(new_n466_), .B1(new_n467_), .B2(new_n459_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(new_n465_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n461_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(G113gat), .B(G141gat), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(new_n307_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(new_n247_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n470_), .A2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n473_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n461_), .A2(new_n469_), .A3(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n474_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n434_), .A2(KEYINPUT101), .A3(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(KEYINPUT101), .B1(new_n434_), .B2(new_n477_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(G230gat), .A2(G233gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(KEYINPUT64), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G85gat), .B(G92gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT65), .B(KEYINPUT9), .ZN(new_n485_));
  XNOR2_X1  g284(.A(KEYINPUT10), .B(G99gat), .ZN(new_n486_));
  OAI22_X1  g285(.A1(new_n484_), .A2(new_n485_), .B1(new_n486_), .B2(G106gat), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT66), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT66), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n491_), .A2(KEYINPUT6), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G99gat), .A2(G106gat), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n490_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n493_), .B1(new_n490_), .B2(new_n492_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G85gat), .A2(G92gat), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n488_), .B(new_n496_), .C1(KEYINPUT9), .C2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n490_), .A2(new_n492_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n493_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n502_));
  INV_X1    g301(.A(new_n502_), .ZN(new_n503_));
  NOR3_X1   g302(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n490_), .A2(new_n492_), .A3(new_n493_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n501_), .A2(new_n505_), .A3(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT8), .ZN(new_n508_));
  INV_X1    g307(.A(new_n484_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n510_));
  AOI21_X1  g309(.A(new_n508_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n498_), .B1(new_n510_), .B2(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G71gat), .B(G78gat), .Z(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G57gat), .B(G64gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT11), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n514_), .A2(new_n516_), .ZN(new_n517_));
  OR2_X1    g316(.A1(new_n515_), .A2(KEYINPUT11), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n513_), .A2(KEYINPUT11), .A3(new_n515_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n517_), .A2(new_n518_), .A3(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n512_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n520_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n498_), .B(new_n522_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n483_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n524_));
  XOR2_X1   g323(.A(new_n524_), .B(KEYINPUT67), .Z(new_n525_));
  NAND2_X1  g324(.A1(new_n520_), .A2(KEYINPUT12), .ZN(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n498_), .B(KEYINPUT68), .C1(new_n510_), .C2(new_n511_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT7), .ZN(new_n530_));
  INV_X1    g329(.A(G99gat), .ZN(new_n531_));
  INV_X1    g330(.A(G106gat), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n533_), .A2(new_n502_), .ZN(new_n534_));
  NOR3_X1   g333(.A1(new_n494_), .A2(new_n495_), .A3(new_n534_), .ZN(new_n535_));
  OAI21_X1  g334(.A(KEYINPUT8), .B1(new_n535_), .B2(new_n484_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n507_), .A2(new_n508_), .A3(new_n509_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  AOI21_X1  g337(.A(KEYINPUT68), .B1(new_n538_), .B2(new_n498_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n527_), .B1(new_n529_), .B2(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT12), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n497_), .A2(KEYINPUT9), .ZN(new_n542_));
  NOR4_X1   g341(.A1(new_n487_), .A2(new_n542_), .A3(new_n495_), .A4(new_n494_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n543_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n541_), .B1(new_n544_), .B2(new_n522_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT69), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n540_), .A2(new_n546_), .ZN(new_n547_));
  OAI211_X1 g346(.A(KEYINPUT69), .B(new_n527_), .C1(new_n529_), .C2(new_n539_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n523_), .A2(new_n483_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(KEYINPUT70), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT70), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n523_), .A2(new_n551_), .A3(new_n483_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n550_), .A2(new_n552_), .ZN(new_n553_));
  NAND3_X1  g352(.A1(new_n547_), .A2(new_n548_), .A3(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n525_), .A2(new_n554_), .ZN(new_n555_));
  XOR2_X1   g354(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n556_));
  XNOR2_X1  g355(.A(G120gat), .B(G148gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G176gat), .B(G204gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n558_), .B(new_n559_), .ZN(new_n560_));
  OR2_X1    g359(.A1(new_n555_), .A2(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n555_), .A2(new_n560_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  XOR2_X1   g362(.A(KEYINPUT72), .B(KEYINPUT13), .Z(new_n564_));
  NOR2_X1   g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n566_));
  AOI21_X1  g365(.A(new_n566_), .B1(new_n561_), .B2(new_n562_), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n481_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n544_), .A2(new_n453_), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n571_), .B(KEYINPUT75), .Z(new_n572_));
  OAI21_X1  g371(.A(new_n454_), .B1(new_n539_), .B2(new_n529_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(new_n574_));
  XOR2_X1   g373(.A(KEYINPUT74), .B(KEYINPUT35), .Z(new_n575_));
  NAND2_X1  g374(.A1(G232gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT73), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT34), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n574_), .A2(new_n575_), .A3(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n575_), .ZN(new_n580_));
  OR2_X1    g379(.A1(new_n578_), .A2(new_n575_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n572_), .A2(new_n573_), .A3(new_n580_), .A4(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n579_), .A2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(KEYINPUT77), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT76), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(G134gat), .ZN(new_n587_));
  INV_X1    g386(.A(G162gat), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(new_n589_), .B(KEYINPUT36), .Z(new_n590_));
  INV_X1    g389(.A(KEYINPUT77), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n579_), .A2(new_n582_), .A3(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n584_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n589_), .A2(KEYINPUT36), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n583_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n593_), .A2(new_n596_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT37), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n583_), .A2(new_n590_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n596_), .A2(KEYINPUT37), .A3(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(KEYINPUT80), .B(KEYINPUT81), .Z(new_n603_));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n448_), .B(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(new_n522_), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G127gat), .B(G155gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT16), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(new_n291_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n610_), .B(G211gat), .ZN(new_n611_));
  INV_X1    g410(.A(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n607_), .B1(KEYINPUT17), .B2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT17), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n611_), .B(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n607_), .A2(new_n615_), .ZN(new_n616_));
  NOR2_X1   g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n602_), .A2(new_n617_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n570_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n240_), .B(KEYINPUT102), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n437_), .A3(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n617_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n597_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n434_), .A2(new_n627_), .A3(new_n477_), .A4(new_n569_), .ZN(new_n628_));
  OAI21_X1  g427(.A(G1gat), .B1(new_n628_), .B2(new_n421_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n622_), .A2(new_n623_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n624_), .A2(new_n629_), .A3(new_n630_), .ZN(G1324gat));
  NAND3_X1  g430(.A1(new_n405_), .A2(new_n391_), .A3(new_n410_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G8gat), .B1(new_n628_), .B2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT39), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n438_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n635_), .B1(new_n619_), .B2(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT40), .Z(G1325gat));
  OAI21_X1  g437(.A(G15gat), .B1(new_n628_), .B2(new_n431_), .ZN(new_n639_));
  XOR2_X1   g438(.A(new_n639_), .B(KEYINPUT41), .Z(new_n640_));
  OR2_X1    g439(.A1(new_n431_), .A2(G15gat), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n640_), .B1(new_n619_), .B2(new_n641_), .ZN(G1326gat));
  OAI21_X1  g441(.A(G22gat), .B1(new_n628_), .B2(new_n432_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n644_));
  XNOR2_X1  g443(.A(new_n643_), .B(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT104), .ZN(new_n646_));
  OAI21_X1  g445(.A(new_n646_), .B1(new_n432_), .B2(G22gat), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n620_), .A2(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n432_), .A2(new_n646_), .A3(G22gat), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(G1327gat));
  INV_X1    g449(.A(KEYINPUT107), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT44), .ZN(new_n652_));
  OAI211_X1 g451(.A(new_n617_), .B(new_n477_), .C1(new_n565_), .C2(new_n567_), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(KEYINPUT105), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n338_), .A2(new_n345_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n655_), .A2(new_n421_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n632_), .A2(new_n656_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n402_), .A2(KEYINPUT99), .A3(new_n422_), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n424_), .B1(new_n408_), .B2(new_n425_), .ZN(new_n659_));
  OAI211_X1 g458(.A(new_n240_), .B(new_n429_), .C1(new_n658_), .C2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n433_), .B1(new_n660_), .B2(new_n418_), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n602_), .B1(new_n657_), .B2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n662_), .A2(KEYINPUT43), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT43), .ZN(new_n664_));
  OAI211_X1 g463(.A(new_n664_), .B(new_n602_), .C1(new_n657_), .C2(new_n661_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n654_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n652_), .B1(new_n666_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n665_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n664_), .B1(new_n434_), .B2(new_n602_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  OAI211_X1 g470(.A(KEYINPUT106), .B(KEYINPUT44), .C1(new_n671_), .C2(new_n654_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n668_), .A2(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n621_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n651_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n673_), .A2(KEYINPUT107), .A3(new_n621_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(G29gat), .A3(new_n677_), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n625_), .A2(new_n597_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n481_), .A2(KEYINPUT108), .A3(new_n569_), .A4(new_n679_), .ZN(new_n680_));
  OAI211_X1 g479(.A(new_n569_), .B(new_n679_), .C1(new_n479_), .C2(new_n480_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT108), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n680_), .A2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  OR2_X1    g484(.A1(new_n421_), .A2(G29gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n678_), .B1(new_n685_), .B2(new_n686_), .ZN(G1328gat));
  INV_X1    g486(.A(KEYINPUT46), .ZN(new_n688_));
  INV_X1    g487(.A(KEYINPUT109), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n673_), .B2(new_n632_), .ZN(new_n690_));
  AOI211_X1 g489(.A(KEYINPUT109), .B(new_n633_), .C1(new_n668_), .C2(new_n672_), .ZN(new_n691_));
  INV_X1    g490(.A(G36gat), .ZN(new_n692_));
  NOR3_X1   g491(.A1(new_n690_), .A2(new_n691_), .A3(new_n692_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n680_), .A2(new_n692_), .A3(new_n683_), .A4(new_n632_), .ZN(new_n694_));
  XNOR2_X1  g493(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n688_), .B1(new_n693_), .B2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n690_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n691_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n698_), .A2(new_n699_), .A3(G36gat), .ZN(new_n700_));
  INV_X1    g499(.A(new_n695_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n694_), .B(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n700_), .A2(new_n702_), .A3(KEYINPUT46), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n697_), .A2(new_n703_), .ZN(G1329gat));
  OAI21_X1  g503(.A(G43gat), .B1(new_n674_), .B2(new_n431_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n431_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n684_), .A2(new_n450_), .A3(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n708_), .B(new_n709_), .ZN(G1330gat));
  OAI21_X1  g509(.A(G50gat), .B1(new_n674_), .B2(new_n432_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n432_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n684_), .A2(new_n452_), .A3(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(G1331gat));
  AND4_X1   g513(.A1(new_n474_), .A2(new_n434_), .A3(new_n476_), .A4(new_n568_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(new_n627_), .ZN(new_n716_));
  INV_X1    g515(.A(G57gat), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n716_), .A2(new_n717_), .A3(new_n421_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n715_), .A2(new_n621_), .A3(new_n618_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n717_), .B2(new_n719_), .ZN(G1332gat));
  OAI21_X1  g519(.A(G64gat), .B1(new_n716_), .B2(new_n633_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT48), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n715_), .A2(new_n618_), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n633_), .A2(G64gat), .ZN(new_n724_));
  OAI21_X1  g523(.A(new_n722_), .B1(new_n723_), .B2(new_n724_), .ZN(G1333gat));
  OAI21_X1  g524(.A(G71gat), .B1(new_n716_), .B2(new_n431_), .ZN(new_n726_));
  XNOR2_X1  g525(.A(new_n726_), .B(KEYINPUT49), .ZN(new_n727_));
  OR2_X1    g526(.A1(new_n431_), .A2(G71gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n723_), .B2(new_n728_), .ZN(G1334gat));
  OAI21_X1  g528(.A(G78gat), .B1(new_n716_), .B2(new_n432_), .ZN(new_n730_));
  XOR2_X1   g529(.A(new_n730_), .B(KEYINPUT50), .Z(new_n731_));
  NOR3_X1   g530(.A1(new_n723_), .A2(G78gat), .A3(new_n432_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT111), .ZN(G1335gat));
  INV_X1    g533(.A(KEYINPUT112), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n735_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n736_));
  NOR3_X1   g535(.A1(new_n569_), .A2(new_n625_), .A3(new_n477_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n663_), .A2(KEYINPUT112), .A3(new_n665_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n736_), .A2(new_n737_), .A3(new_n738_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT113), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND4_X1  g540(.A1(new_n736_), .A2(new_n738_), .A3(KEYINPUT113), .A4(new_n737_), .ZN(new_n742_));
  AND4_X1   g541(.A1(G85gat), .A2(new_n741_), .A3(new_n240_), .A4(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n715_), .A2(new_n679_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(G85gat), .B1(new_n745_), .B2(new_n621_), .ZN(new_n746_));
  NOR2_X1   g545(.A1(new_n743_), .A2(new_n746_), .ZN(G1336gat));
  NAND4_X1  g546(.A1(new_n741_), .A2(G92gat), .A3(new_n632_), .A4(new_n742_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n372_), .B1(new_n744_), .B2(new_n633_), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n748_), .A2(new_n749_), .ZN(G1337gat));
  OR3_X1    g549(.A1(new_n744_), .A2(new_n486_), .A3(new_n431_), .ZN(new_n751_));
  NAND3_X1  g550(.A1(new_n741_), .A2(new_n706_), .A3(new_n742_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT114), .ZN(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(new_n753_), .A3(G99gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G99gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n757_), .A2(KEYINPUT115), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  OAI221_X1 g558(.A(new_n751_), .B1(KEYINPUT115), .B2(new_n757_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n759_), .A2(new_n760_), .ZN(G1338gat));
  NAND3_X1  g560(.A1(new_n745_), .A2(new_n532_), .A3(new_n712_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n712_), .B(new_n737_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n763_), .A2(new_n764_), .A3(G106gat), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n764_), .B1(new_n763_), .B2(G106gat), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n762_), .B1(new_n765_), .B2(new_n766_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n767_), .A2(KEYINPUT116), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(KEYINPUT116), .ZN(new_n769_));
  AND3_X1   g568(.A1(new_n768_), .A2(KEYINPUT53), .A3(new_n769_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT53), .B1(new_n768_), .B2(new_n769_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1339gat));
  INV_X1    g571(.A(KEYINPUT56), .ZN(new_n773_));
  NAND4_X1  g572(.A1(new_n547_), .A2(KEYINPUT55), .A3(new_n548_), .A4(new_n553_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT119), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT68), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n512_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n526_), .B1(new_n777_), .B2(new_n528_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT69), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n779_), .B1(new_n521_), .B2(new_n541_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n548_), .B(new_n523_), .C1(new_n778_), .C2(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(KEYINPUT118), .ZN(new_n782_));
  INV_X1    g581(.A(new_n483_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT118), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n547_), .A2(new_n784_), .A3(new_n548_), .A4(new_n523_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n782_), .A2(new_n783_), .A3(new_n785_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n548_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n553_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n787_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  INV_X1    g589(.A(KEYINPUT117), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n554_), .A2(KEYINPUT117), .A3(new_n787_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n775_), .A2(new_n786_), .A3(new_n792_), .A4(new_n793_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n773_), .B1(new_n794_), .B2(new_n560_), .ZN(new_n795_));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n774_), .A2(new_n796_), .ZN(new_n797_));
  INV_X1    g596(.A(new_n788_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n798_), .A2(KEYINPUT119), .A3(KEYINPUT55), .A4(new_n553_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n786_), .A2(new_n797_), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n792_), .A2(new_n793_), .ZN(new_n801_));
  OAI211_X1 g600(.A(new_n773_), .B(new_n560_), .C1(new_n800_), .C2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n795_), .A2(new_n803_), .ZN(new_n804_));
  NAND4_X1  g603(.A1(new_n804_), .A2(KEYINPUT120), .A3(new_n477_), .A4(new_n561_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n457_), .A2(new_n465_), .A3(new_n460_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n464_), .A2(new_n458_), .A3(new_n468_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n806_), .A2(new_n807_), .A3(new_n473_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n476_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n563_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n560_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(KEYINPUT56), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n812_), .A2(new_n477_), .A3(new_n561_), .A4(new_n802_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT120), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n805_), .A2(new_n810_), .A3(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n597_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT57), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND4_X1  g618(.A1(new_n812_), .A2(new_n809_), .A3(new_n561_), .A4(new_n802_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT58), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n602_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT121), .ZN(new_n824_));
  OR2_X1    g623(.A1(new_n820_), .A2(new_n821_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT121), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n822_), .A2(new_n826_), .A3(new_n602_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n824_), .A2(new_n825_), .A3(new_n827_), .ZN(new_n828_));
  NAND3_X1  g627(.A1(new_n816_), .A2(KEYINPUT57), .A3(new_n597_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n819_), .A2(new_n828_), .A3(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n830_), .A2(new_n617_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n477_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n618_), .A2(new_n832_), .A3(new_n569_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT54), .ZN(new_n834_));
  XNOR2_X1  g633(.A(new_n833_), .B(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n831_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n338_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n675_), .A2(new_n632_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(new_n840_), .ZN(new_n841_));
  AOI21_X1  g640(.A(G113gat), .B1(new_n841_), .B2(new_n477_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT122), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT59), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n840_), .A2(new_n843_), .A3(new_n844_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n839_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n846_), .B1(new_n831_), .B2(new_n836_), .ZN(new_n847_));
  XOR2_X1   g646(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n848_));
  NAND3_X1  g647(.A1(new_n847_), .A2(new_n838_), .A3(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n832_), .B1(new_n845_), .B2(new_n849_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n842_), .B1(new_n850_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g650(.A(G120gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n852_), .B1(new_n569_), .B2(KEYINPUT60), .ZN(new_n853_));
  OAI211_X1 g652(.A(new_n841_), .B(new_n853_), .C1(KEYINPUT60), .C2(new_n852_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n569_), .B1(new_n845_), .B2(new_n849_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(new_n852_), .ZN(G1341gat));
  NAND2_X1  g655(.A1(new_n843_), .A2(new_n844_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n857_), .B1(new_n847_), .B2(new_n838_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n835_), .B1(new_n830_), .B2(new_n617_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n848_), .ZN(new_n860_));
  NOR4_X1   g659(.A1(new_n859_), .A2(new_n338_), .A3(new_n846_), .A4(new_n860_), .ZN(new_n861_));
  OAI211_X1 g660(.A(G127gat), .B(new_n625_), .C1(new_n858_), .C2(new_n861_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT123), .ZN(new_n863_));
  INV_X1    g662(.A(G127gat), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n863_), .B(new_n864_), .C1(new_n840_), .C2(new_n617_), .ZN(new_n865_));
  NOR4_X1   g664(.A1(new_n859_), .A2(new_n617_), .A3(new_n338_), .A4(new_n846_), .ZN(new_n866_));
  OAI21_X1  g665(.A(KEYINPUT123), .B1(new_n866_), .B2(G127gat), .ZN(new_n867_));
  AND3_X1   g666(.A1(new_n862_), .A2(new_n865_), .A3(new_n867_), .ZN(G1342gat));
  INV_X1    g667(.A(new_n597_), .ZN(new_n869_));
  AOI21_X1  g668(.A(G134gat), .B1(new_n841_), .B2(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n602_), .ZN(new_n871_));
  AOI21_X1  g670(.A(new_n871_), .B1(new_n845_), .B2(new_n849_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n870_), .B1(new_n872_), .B2(G134gat), .ZN(G1343gat));
  NOR3_X1   g672(.A1(new_n859_), .A2(new_n345_), .A3(new_n846_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n477_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n568_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g677(.A1(new_n874_), .A2(new_n625_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(KEYINPUT61), .B(G155gat), .ZN(new_n880_));
  XNOR2_X1  g679(.A(new_n879_), .B(new_n880_), .ZN(G1346gat));
  AOI21_X1  g680(.A(G162gat), .B1(new_n874_), .B2(new_n869_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n871_), .A2(new_n588_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n882_), .B1(new_n874_), .B2(new_n883_), .ZN(G1347gat));
  INV_X1    g683(.A(KEYINPUT62), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n859_), .A2(new_n338_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n633_), .A2(new_n621_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n886_), .A2(new_n477_), .A3(new_n887_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n885_), .B1(new_n888_), .B2(new_n307_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n358_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n886_), .A2(new_n887_), .ZN(new_n891_));
  OAI211_X1 g690(.A(KEYINPUT62), .B(G169gat), .C1(new_n891_), .C2(new_n832_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n889_), .A2(new_n890_), .A3(new_n892_), .ZN(G1348gat));
  NAND3_X1  g692(.A1(new_n886_), .A2(new_n568_), .A3(new_n887_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G176gat), .ZN(G1349gat));
  NOR2_X1   g694(.A1(new_n891_), .A2(new_n617_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n896_), .A2(new_n351_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n897_), .B1(new_n896_), .B2(new_n291_), .ZN(G1350gat));
  OAI21_X1  g697(.A(G190gat), .B1(new_n891_), .B2(new_n871_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n886_), .A2(new_n352_), .A3(new_n887_), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n597_), .B2(new_n900_), .ZN(G1351gat));
  NOR3_X1   g700(.A1(new_n633_), .A2(new_n240_), .A3(new_n345_), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n837_), .A2(new_n902_), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n903_), .A2(new_n832_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(new_n247_), .ZN(G1352gat));
  OAI22_X1  g704(.A1(new_n903_), .A2(new_n569_), .B1(KEYINPUT124), .B2(G204gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n907_));
  XOR2_X1   g706(.A(new_n907_), .B(KEYINPUT125), .Z(new_n908_));
  XNOR2_X1  g707(.A(new_n906_), .B(new_n908_), .ZN(G1353gat));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n617_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT126), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n903_), .A2(new_n912_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n914_));
  INV_X1    g713(.A(new_n914_), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n910_), .B1(new_n913_), .B2(new_n915_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n913_), .A2(new_n915_), .ZN(new_n917_));
  OAI211_X1 g716(.A(KEYINPUT127), .B(new_n914_), .C1(new_n903_), .C2(new_n912_), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n916_), .A2(new_n917_), .A3(new_n918_), .ZN(G1354gat));
  AND2_X1   g718(.A1(new_n837_), .A2(new_n902_), .ZN(new_n920_));
  AND3_X1   g719(.A1(new_n920_), .A2(G218gat), .A3(new_n602_), .ZN(new_n921_));
  AOI21_X1  g720(.A(G218gat), .B1(new_n920_), .B2(new_n869_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1355gat));
endmodule


