//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 0 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n575_,
    new_n576_, new_n577_, new_n578_, new_n579_, new_n580_, new_n581_,
    new_n583_, new_n584_, new_n585_, new_n586_, new_n587_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n814_, new_n815_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n842_, new_n843_, new_n845_, new_n846_,
    new_n847_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G85gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G57gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  XOR2_X1   g005(.A(G127gat), .B(G134gat), .Z(new_n207_));
  XOR2_X1   g006(.A(G113gat), .B(G120gat), .Z(new_n208_));
  XOR2_X1   g007(.A(new_n207_), .B(new_n208_), .Z(new_n209_));
  OR3_X1    g008(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT2), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  NAND3_X1  g012(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n210_), .A2(new_n213_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217_));
  OR2_X1    g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n217_), .A3(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(G141gat), .B(G148gat), .Z(new_n220_));
  OAI21_X1  g019(.A(KEYINPUT80), .B1(new_n217_), .B2(KEYINPUT1), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n217_), .A2(KEYINPUT1), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n221_), .A2(new_n222_), .A3(new_n218_), .ZN(new_n223_));
  NOR3_X1   g022(.A1(new_n217_), .A2(KEYINPUT80), .A3(KEYINPUT1), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n220_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n219_), .A2(new_n225_), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT92), .B1(new_n209_), .B2(new_n226_), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n207_), .B(new_n208_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n228_), .B1(new_n225_), .B2(new_n219_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n227_), .B(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT4), .ZN(new_n231_));
  NAND2_X1  g030(.A1(G225gat), .A2(G233gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  XOR2_X1   g032(.A(KEYINPUT93), .B(KEYINPUT4), .Z(new_n234_));
  NAND2_X1  g033(.A1(new_n229_), .A2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n231_), .A2(new_n233_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT94), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT94), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n231_), .A2(new_n238_), .A3(new_n233_), .A4(new_n235_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n230_), .A2(new_n232_), .ZN(new_n241_));
  XNOR2_X1  g040(.A(new_n241_), .B(KEYINPUT95), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n206_), .B1(new_n240_), .B2(new_n242_), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n242_), .A2(new_n239_), .A3(new_n237_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n206_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n244_), .A2(new_n245_), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n243_), .A2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G183gat), .A2(G190gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT23), .ZN(new_n249_));
  NOR2_X1   g048(.A1(G169gat), .A2(G176gat), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT24), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  AND2_X1   g051(.A1(new_n249_), .A2(new_n252_), .ZN(new_n253_));
  OR2_X1    g052(.A1(new_n253_), .A2(KEYINPUT78), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(KEYINPUT78), .ZN(new_n255_));
  INV_X1    g054(.A(G169gat), .ZN(new_n256_));
  INV_X1    g055(.A(G176gat), .ZN(new_n257_));
  OAI21_X1  g056(.A(KEYINPUT24), .B1(new_n256_), .B2(new_n257_), .ZN(new_n258_));
  NOR2_X1   g057(.A1(new_n258_), .A2(new_n250_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(KEYINPUT26), .B(G190gat), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT77), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT25), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n262_), .B1(new_n263_), .B2(G183gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT25), .B(G183gat), .ZN(new_n265_));
  OAI211_X1 g064(.A(new_n261_), .B(new_n264_), .C1(new_n265_), .C2(new_n262_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n254_), .A2(new_n255_), .A3(new_n260_), .A4(new_n266_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n249_), .B1(G183gat), .B2(G190gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n269_));
  XNOR2_X1  g068(.A(new_n269_), .B(new_n256_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n268_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n267_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G227gat), .A2(G233gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n274_), .B(G15gat), .Z(new_n275_));
  XNOR2_X1  g074(.A(new_n273_), .B(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(new_n276_), .B(KEYINPUT31), .Z(new_n277_));
  XNOR2_X1  g076(.A(G71gat), .B(G99gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n278_), .B(G43gat), .ZN(new_n279_));
  XNOR2_X1  g078(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n279_), .B(new_n280_), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n281_), .B(new_n228_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(new_n277_), .B(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n247_), .A2(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G78gat), .B(G106gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n285_), .B(KEYINPUT88), .Z(new_n286_));
  NAND2_X1  g085(.A1(G228gat), .A2(G233gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(G197gat), .ZN(new_n289_));
  INV_X1    g088(.A(G204gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(KEYINPUT84), .B(G197gat), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n291_), .B1(new_n292_), .B2(new_n290_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G211gat), .B(G218gat), .Z(new_n295_));
  NAND3_X1  g094(.A1(new_n294_), .A2(KEYINPUT21), .A3(new_n295_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n295_), .ZN(new_n297_));
  AND2_X1   g096(.A1(new_n292_), .A2(new_n290_), .ZN(new_n298_));
  OAI21_X1  g097(.A(KEYINPUT21), .B1(new_n289_), .B2(new_n290_), .ZN(new_n299_));
  XOR2_X1   g098(.A(KEYINPUT85), .B(KEYINPUT21), .Z(new_n300_));
  OAI221_X1 g099(.A(new_n297_), .B1(new_n298_), .B2(new_n299_), .C1(new_n294_), .C2(new_n300_), .ZN(new_n301_));
  AND2_X1   g100(.A1(new_n301_), .A2(KEYINPUT86), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(KEYINPUT86), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n296_), .B1(new_n302_), .B2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n226_), .A2(KEYINPUT29), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OAI21_X1  g105(.A(new_n288_), .B1(new_n306_), .B2(KEYINPUT87), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT83), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n304_), .A2(new_n308_), .A3(new_n305_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n307_), .B1(KEYINPUT87), .B2(new_n309_), .ZN(new_n310_));
  OAI211_X1 g109(.A(KEYINPUT87), .B(new_n287_), .C1(new_n306_), .C2(KEYINPUT83), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n286_), .B1(new_n310_), .B2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT89), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n313_), .A2(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n309_), .A2(KEYINPUT87), .ZN(new_n316_));
  OAI211_X1 g115(.A(new_n316_), .B(new_n288_), .C1(KEYINPUT87), .C2(new_n306_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n286_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(new_n318_), .A3(new_n311_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT90), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n318_), .B1(new_n317_), .B2(new_n311_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT89), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n317_), .A2(KEYINPUT90), .A3(new_n318_), .A4(new_n311_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n315_), .A2(new_n321_), .A3(new_n323_), .A4(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n226_), .A2(KEYINPUT29), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G22gat), .B(G50gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT82), .ZN(new_n328_));
  XNOR2_X1  g127(.A(new_n326_), .B(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT81), .B(KEYINPUT28), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n329_), .B(new_n330_), .Z(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n325_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n313_), .A2(new_n331_), .A3(new_n319_), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT27), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT19), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  OR2_X1    g137(.A1(new_n304_), .A2(new_n273_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT20), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT91), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n270_), .B1(new_n268_), .B2(new_n341_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n342_), .B1(new_n341_), .B2(new_n268_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n259_), .B1(new_n265_), .B2(new_n261_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n253_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n340_), .B1(new_n304_), .B2(new_n346_), .ZN(new_n347_));
  AOI21_X1  g146(.A(new_n338_), .B1(new_n339_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G8gat), .B(G36gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(KEYINPUT18), .ZN(new_n351_));
  XNOR2_X1  g150(.A(G64gat), .B(G92gat), .ZN(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  NAND2_X1  g152(.A1(new_n304_), .A2(new_n273_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n346_), .ZN(new_n355_));
  OAI211_X1 g154(.A(new_n355_), .B(new_n296_), .C1(new_n302_), .C2(new_n303_), .ZN(new_n356_));
  NAND4_X1  g155(.A1(new_n354_), .A2(new_n356_), .A3(KEYINPUT20), .A4(new_n338_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n349_), .A2(new_n353_), .A3(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n353_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n357_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n359_), .B1(new_n360_), .B2(new_n348_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n358_), .A2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n360_), .A2(new_n348_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n335_), .B1(new_n363_), .B2(new_n353_), .ZN(new_n364_));
  XOR2_X1   g163(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n365_));
  NAND3_X1  g164(.A1(new_n354_), .A2(new_n356_), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n337_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n339_), .A2(new_n347_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n367_), .B1(new_n368_), .B2(new_n337_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n359_), .ZN(new_n370_));
  AOI22_X1  g169(.A1(new_n335_), .A2(new_n362_), .B1(new_n364_), .B2(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n333_), .A2(new_n334_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT98), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT98), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n333_), .A2(new_n374_), .A3(new_n334_), .A4(new_n371_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n284_), .B1(new_n373_), .B2(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n322_), .A2(KEYINPUT89), .ZN(new_n377_));
  AOI211_X1 g176(.A(new_n314_), .B(new_n318_), .C1(new_n317_), .C2(new_n311_), .ZN(new_n378_));
  NOR2_X1   g177(.A1(new_n377_), .A2(new_n378_), .ZN(new_n379_));
  AND2_X1   g178(.A1(new_n321_), .A2(new_n324_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n331_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n334_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n247_), .B(new_n371_), .C1(new_n381_), .C2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n362_), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n240_), .A2(KEYINPUT33), .A3(new_n206_), .A4(new_n242_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n231_), .A2(new_n232_), .A3(new_n235_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT96), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n206_), .B1(new_n230_), .B2(new_n233_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n384_), .A2(new_n385_), .A3(new_n389_), .ZN(new_n390_));
  NOR2_X1   g189(.A1(new_n246_), .A2(KEYINPUT33), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n353_), .A2(KEYINPUT32), .ZN(new_n392_));
  MUX2_X1   g191(.A(new_n369_), .B(new_n363_), .S(new_n392_), .Z(new_n393_));
  OAI22_X1  g192(.A1(new_n390_), .A2(new_n391_), .B1(new_n247_), .B2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n394_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n283_), .B1(new_n383_), .B2(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(new_n376_), .A2(new_n396_), .ZN(new_n397_));
  AND2_X1   g196(.A1(G85gat), .A2(G92gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(KEYINPUT65), .B2(KEYINPUT9), .ZN(new_n399_));
  OAI211_X1 g198(.A(KEYINPUT65), .B(KEYINPUT9), .C1(G85gat), .C2(G92gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n399_), .B(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(G99gat), .A2(G106gat), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT6), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT6), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(G99gat), .A3(G106gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(KEYINPUT10), .B(G99gat), .ZN(new_n407_));
  OAI211_X1 g206(.A(new_n401_), .B(new_n406_), .C1(G106gat), .C2(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(G85gat), .A2(G92gat), .ZN(new_n409_));
  NOR3_X1   g208(.A1(new_n398_), .A2(new_n409_), .A3(KEYINPUT8), .ZN(new_n410_));
  AND2_X1   g209(.A1(new_n403_), .A2(new_n405_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT7), .ZN(new_n412_));
  INV_X1    g211(.A(G99gat), .ZN(new_n413_));
  INV_X1    g212(.A(G106gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n412_), .A2(new_n413_), .A3(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n410_), .B1(new_n411_), .B2(new_n417_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT66), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT66), .ZN(new_n420_));
  OAI211_X1 g219(.A(new_n420_), .B(new_n410_), .C1(new_n411_), .C2(new_n417_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT8), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n406_), .A2(KEYINPUT67), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT67), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n403_), .A2(new_n405_), .A3(new_n425_), .ZN(new_n426_));
  AND2_X1   g225(.A1(new_n415_), .A2(new_n416_), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n424_), .A2(new_n426_), .A3(new_n427_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n398_), .A2(new_n409_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n423_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n408_), .B1(new_n422_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G29gat), .B(G36gat), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G43gat), .B(G50gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT35), .ZN(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT70), .B(KEYINPUT34), .ZN(new_n437_));
  NAND2_X1  g236(.A1(G232gat), .A2(G233gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n432_), .A2(new_n435_), .B1(new_n436_), .B2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT68), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n431_), .A2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n429_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n417_), .B1(KEYINPUT67), .B2(new_n406_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n443_), .B1(new_n444_), .B2(new_n426_), .ZN(new_n445_));
  OAI211_X1 g244(.A(new_n419_), .B(new_n421_), .C1(new_n445_), .C2(new_n423_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n446_), .A2(KEYINPUT68), .A3(new_n408_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n435_), .B(KEYINPUT15), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n442_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n439_), .A2(new_n436_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  AND3_X1   g250(.A1(new_n440_), .A2(new_n449_), .A3(new_n451_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n451_), .B1(new_n440_), .B2(new_n449_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G190gat), .B(G218gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(G134gat), .B(G162gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  OR4_X1    g255(.A1(KEYINPUT36), .A2(new_n452_), .A3(new_n453_), .A4(new_n456_), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(KEYINPUT36), .Z(new_n458_));
  OAI21_X1  g257(.A(new_n458_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n457_), .A2(new_n459_), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n397_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G57gat), .B(G64gat), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n462_), .A2(KEYINPUT11), .ZN(new_n463_));
  XOR2_X1   g262(.A(G71gat), .B(G78gat), .Z(new_n464_));
  NOR2_X1   g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  AND2_X1   g264(.A1(new_n463_), .A2(new_n464_), .ZN(new_n466_));
  OR2_X1    g265(.A1(new_n462_), .A2(KEYINPUT11), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n465_), .B1(new_n466_), .B2(new_n467_), .ZN(new_n468_));
  NAND4_X1  g267(.A1(new_n442_), .A2(new_n447_), .A3(KEYINPUT12), .A4(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G230gat), .A2(G233gat), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n470_), .B(KEYINPUT64), .Z(new_n471_));
  INV_X1    g270(.A(new_n468_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n471_), .B1(new_n432_), .B2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT69), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n431_), .A2(new_n468_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT12), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  AOI211_X1 g276(.A(KEYINPUT69), .B(KEYINPUT12), .C1(new_n431_), .C2(new_n468_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n469_), .B(new_n473_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n432_), .A2(new_n472_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n472_), .B1(new_n446_), .B2(new_n408_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n471_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n479_), .A2(new_n483_), .ZN(new_n484_));
  XOR2_X1   g283(.A(G120gat), .B(G148gat), .Z(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT5), .ZN(new_n486_));
  XNOR2_X1  g285(.A(G176gat), .B(G204gat), .ZN(new_n487_));
  XNOR2_X1  g286(.A(new_n486_), .B(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n484_), .B(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT13), .ZN(new_n490_));
  OR2_X1    g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n489_), .A2(new_n490_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G15gat), .B(G22gat), .ZN(new_n494_));
  INV_X1    g293(.A(G8gat), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(G1gat), .B(G8gat), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n498_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(new_n435_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT75), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G229gat), .A2(G233gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n501_), .A2(new_n435_), .ZN(new_n505_));
  OR3_X1    g304(.A1(new_n503_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n504_), .ZN(new_n507_));
  INV_X1    g306(.A(new_n501_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n503_), .B1(new_n508_), .B2(new_n448_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n506_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G113gat), .B(G141gat), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G169gat), .B(G197gat), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n511_), .B(new_n512_), .Z(new_n513_));
  OR2_X1    g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(KEYINPUT76), .A3(new_n513_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n515_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT76), .B1(new_n510_), .B2(new_n513_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n514_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n518_), .ZN(new_n519_));
  NOR2_X1   g318(.A1(new_n493_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(G231gat), .A2(G233gat), .ZN(new_n521_));
  XNOR2_X1  g320(.A(new_n501_), .B(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(new_n468_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G127gat), .B(G155gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT73), .B(KEYINPUT16), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n524_), .B(new_n525_), .ZN(new_n526_));
  XOR2_X1   g325(.A(G183gat), .B(G211gat), .Z(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n529_));
  NOR3_X1   g328(.A1(new_n528_), .A2(KEYINPUT72), .A3(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n528_), .A2(new_n529_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n523_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  OAI21_X1  g331(.A(new_n532_), .B1(new_n530_), .B2(new_n523_), .ZN(new_n533_));
  XOR2_X1   g332(.A(new_n533_), .B(KEYINPUT74), .Z(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n520_), .A2(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT99), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n461_), .A2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(new_n247_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n202_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n397_), .A2(new_n518_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT71), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n457_), .A2(new_n543_), .A3(new_n459_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(KEYINPUT37), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(new_n535_), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(new_n493_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n542_), .A2(new_n547_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n548_), .A2(G1gat), .A3(new_n247_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n541_), .B1(KEYINPUT38), .B2(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n542_), .A2(new_n547_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n551_), .A2(new_n202_), .A3(new_n540_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT100), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT38), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n553_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n550_), .B1(new_n556_), .B2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(KEYINPUT101), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT101), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n550_), .B(new_n560_), .C1(new_n556_), .C2(new_n557_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n559_), .A2(new_n561_), .ZN(G1324gat));
  INV_X1    g361(.A(new_n371_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n551_), .A2(new_n495_), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n495_), .B1(new_n539_), .B2(new_n563_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT39), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n565_), .A2(new_n566_), .ZN(new_n569_));
  OAI21_X1  g368(.A(new_n564_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT40), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  OAI211_X1 g371(.A(KEYINPUT40), .B(new_n564_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n572_), .A2(new_n573_), .ZN(G1325gat));
  INV_X1    g373(.A(new_n283_), .ZN(new_n575_));
  OAI21_X1  g374(.A(G15gat), .B1(new_n538_), .B2(new_n575_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT102), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT41), .ZN(new_n578_));
  OR2_X1    g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n578_), .ZN(new_n580_));
  OR3_X1    g379(.A1(new_n548_), .A2(G15gat), .A3(new_n575_), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .ZN(G1326gat));
  NAND2_X1  g381(.A1(new_n333_), .A2(new_n334_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  OAI21_X1  g383(.A(G22gat), .B1(new_n538_), .B2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT42), .ZN(new_n586_));
  OR2_X1    g385(.A1(new_n584_), .A2(G22gat), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n586_), .B1(new_n548_), .B2(new_n587_), .ZN(G1327gat));
  INV_X1    g387(.A(new_n545_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n376_), .B2(new_n396_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT43), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n590_), .A2(new_n591_), .ZN(new_n592_));
  OAI211_X1 g391(.A(KEYINPUT43), .B(new_n589_), .C1(new_n376_), .C2(new_n396_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n592_), .A2(new_n534_), .A3(new_n520_), .A4(new_n593_), .ZN(new_n594_));
  XOR2_X1   g393(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n535_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT44), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n597_), .A2(new_n598_), .A3(new_n520_), .A4(new_n593_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n247_), .B1(new_n596_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(G29gat), .ZN(new_n601_));
  INV_X1    g400(.A(new_n460_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n534_), .A2(new_n602_), .ZN(new_n603_));
  XOR2_X1   g402(.A(new_n603_), .B(KEYINPUT104), .Z(new_n604_));
  NOR2_X1   g403(.A1(new_n604_), .A2(new_n493_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n397_), .A2(new_n518_), .A3(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n540_), .A2(new_n601_), .ZN(new_n607_));
  OAI22_X1  g406(.A1(new_n600_), .A2(new_n601_), .B1(new_n606_), .B2(new_n607_), .ZN(G1328gat));
  NOR2_X1   g407(.A1(new_n371_), .A2(G36gat), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  OR3_X1    g409(.A1(new_n606_), .A2(KEYINPUT106), .A3(new_n610_), .ZN(new_n611_));
  OAI21_X1  g410(.A(KEYINPUT106), .B1(new_n606_), .B2(new_n610_), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n611_), .A2(KEYINPUT45), .A3(new_n612_), .ZN(new_n613_));
  AOI21_X1  g412(.A(KEYINPUT45), .B1(new_n611_), .B2(new_n612_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n596_), .A2(new_n599_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT105), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(new_n617_), .A3(new_n563_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(G36gat), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n617_), .B1(new_n616_), .B2(new_n563_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n615_), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT108), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  OAI211_X1 g424(.A(new_n623_), .B(new_n615_), .C1(new_n619_), .C2(new_n620_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(G1329gat));
  AOI21_X1  g426(.A(new_n575_), .B1(new_n596_), .B2(new_n599_), .ZN(new_n628_));
  INV_X1    g427(.A(G43gat), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n283_), .A2(new_n629_), .ZN(new_n630_));
  OAI22_X1  g429(.A1(new_n628_), .A2(new_n629_), .B1(new_n606_), .B2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT47), .Z(G1330gat));
  AOI21_X1  g431(.A(new_n584_), .B1(new_n596_), .B2(new_n599_), .ZN(new_n633_));
  INV_X1    g432(.A(G50gat), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n583_), .A2(new_n634_), .ZN(new_n635_));
  XOR2_X1   g434(.A(new_n635_), .B(KEYINPUT109), .Z(new_n636_));
  OAI22_X1  g435(.A1(new_n633_), .A2(new_n634_), .B1(new_n606_), .B2(new_n636_), .ZN(G1331gat));
  NAND4_X1  g436(.A1(new_n461_), .A2(new_n519_), .A3(new_n493_), .A4(new_n535_), .ZN(new_n638_));
  INV_X1    g437(.A(G57gat), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n247_), .ZN(new_n640_));
  AND3_X1   g439(.A1(new_n397_), .A2(KEYINPUT110), .A3(new_n519_), .ZN(new_n641_));
  AOI21_X1  g440(.A(KEYINPUT110), .B1(new_n397_), .B2(new_n519_), .ZN(new_n642_));
  NOR2_X1   g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  INV_X1    g442(.A(new_n493_), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n643_), .A2(new_n644_), .A3(new_n546_), .ZN(new_n645_));
  AOI21_X1  g444(.A(G57gat), .B1(new_n645_), .B2(new_n540_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n646_), .A2(KEYINPUT111), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(KEYINPUT111), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n640_), .B1(new_n647_), .B2(new_n648_), .ZN(G1332gat));
  OAI21_X1  g448(.A(G64gat), .B1(new_n638_), .B2(new_n371_), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n650_), .B(KEYINPUT48), .ZN(new_n651_));
  INV_X1    g450(.A(G64gat), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n645_), .A2(new_n652_), .A3(new_n563_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(G1333gat));
  OAI21_X1  g453(.A(G71gat), .B1(new_n638_), .B2(new_n575_), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n655_), .B(KEYINPUT49), .ZN(new_n656_));
  INV_X1    g455(.A(G71gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n645_), .A2(new_n657_), .A3(new_n283_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n656_), .A2(new_n658_), .ZN(G1334gat));
  OAI21_X1  g458(.A(G78gat), .B1(new_n638_), .B2(new_n584_), .ZN(new_n660_));
  OR2_X1    g459(.A1(new_n660_), .A2(KEYINPUT112), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n660_), .A2(KEYINPUT112), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT50), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n661_), .A2(KEYINPUT50), .A3(new_n662_), .ZN(new_n666_));
  INV_X1    g465(.A(G78gat), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n645_), .A2(new_n667_), .A3(new_n583_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n665_), .A2(new_n666_), .A3(new_n668_), .ZN(G1335gat));
  NOR2_X1   g468(.A1(new_n644_), .A2(new_n518_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n597_), .A2(new_n593_), .A3(new_n670_), .ZN(new_n671_));
  OAI21_X1  g470(.A(G85gat), .B1(new_n671_), .B2(new_n247_), .ZN(new_n672_));
  OR3_X1    g471(.A1(new_n643_), .A2(new_n644_), .A3(new_n604_), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n247_), .A2(G85gat), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n672_), .B1(new_n673_), .B2(new_n674_), .ZN(G1336gat));
  OAI21_X1  g474(.A(G92gat), .B1(new_n671_), .B2(new_n371_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n371_), .A2(G92gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n673_), .B2(new_n677_), .ZN(G1337gat));
  OAI21_X1  g477(.A(G99gat), .B1(new_n671_), .B2(new_n575_), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n575_), .A2(new_n407_), .ZN(new_n680_));
  OAI21_X1  g479(.A(new_n679_), .B1(new_n673_), .B2(new_n680_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI21_X1  g481(.A(G106gat), .B1(new_n671_), .B2(new_n584_), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n683_), .A2(KEYINPUT113), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT52), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n683_), .B2(KEYINPUT113), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n683_), .A2(KEYINPUT113), .A3(new_n685_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n583_), .A2(new_n414_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n689_), .B1(new_n673_), .B2(new_n690_), .ZN(new_n691_));
  OAI21_X1  g490(.A(KEYINPUT53), .B1(new_n688_), .B2(new_n691_), .ZN(new_n692_));
  OR2_X1    g491(.A1(new_n673_), .A2(new_n690_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT53), .ZN(new_n694_));
  NAND4_X1  g493(.A1(new_n693_), .A2(new_n687_), .A3(new_n694_), .A4(new_n689_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n692_), .A2(new_n695_), .ZN(G1339gat));
  OR2_X1    g495(.A1(new_n484_), .A2(new_n488_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n518_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n479_), .A2(KEYINPUT55), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT69), .B1(new_n482_), .B2(KEYINPUT12), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n475_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT55), .ZN(new_n704_));
  NAND4_X1  g503(.A1(new_n703_), .A2(new_n704_), .A3(new_n469_), .A4(new_n473_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n700_), .A2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(new_n480_), .B(new_n469_), .C1(new_n477_), .C2(new_n478_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n471_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n706_), .A2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT115), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n706_), .A2(KEYINPUT115), .A3(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(new_n713_));
  AOI21_X1  g512(.A(KEYINPUT56), .B1(new_n713_), .B2(new_n488_), .ZN(new_n714_));
  AOI221_X4 g513(.A(new_n710_), .B1(new_n707_), .B2(new_n471_), .C1(new_n700_), .C2(new_n705_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT115), .B1(new_n706_), .B2(new_n708_), .ZN(new_n716_));
  OAI211_X1 g515(.A(KEYINPUT56), .B(new_n488_), .C1(new_n715_), .C2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  OAI21_X1  g517(.A(new_n699_), .B1(new_n714_), .B2(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT116), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n488_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT56), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n698_), .B1(new_n723_), .B2(new_n717_), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT116), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n510_), .A2(new_n513_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT76), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  OR2_X1    g528(.A1(new_n503_), .A2(new_n505_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n513_), .B1(new_n730_), .B2(new_n504_), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT117), .ZN(new_n732_));
  OR2_X1    g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  AOI22_X1  g532(.A1(new_n731_), .A2(new_n732_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n734_));
  AOI22_X1  g533(.A1(new_n729_), .A2(new_n515_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n735_), .A2(new_n489_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT118), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n735_), .A2(new_n489_), .A3(KEYINPUT118), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n720_), .A2(new_n726_), .A3(new_n740_), .ZN(new_n741_));
  AOI21_X1  g540(.A(KEYINPUT57), .B1(new_n741_), .B2(new_n460_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT57), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n602_), .A2(new_n743_), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n740_), .B1(new_n724_), .B2(new_n725_), .ZN(new_n745_));
  AOI211_X1 g544(.A(KEYINPUT116), .B(new_n698_), .C1(new_n723_), .C2(new_n717_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n744_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n735_), .A2(new_n697_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n723_), .B2(new_n717_), .ZN(new_n749_));
  OR2_X1    g548(.A1(new_n749_), .A2(KEYINPUT58), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n545_), .B1(new_n749_), .B2(KEYINPUT58), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n747_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n534_), .B1(new_n742_), .B2(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n535_), .A2(new_n519_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT114), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n756_), .A2(new_n644_), .A3(new_n545_), .ZN(new_n757_));
  XNOR2_X1  g556(.A(new_n757_), .B(KEYINPUT54), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n754_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT59), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n373_), .A2(new_n375_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(new_n540_), .A3(new_n283_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n759_), .A2(new_n760_), .A3(new_n763_), .ZN(new_n764_));
  INV_X1    g563(.A(G113gat), .ZN(new_n765_));
  NOR2_X1   g564(.A1(new_n519_), .A2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT119), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n767_), .B1(new_n742_), .B2(new_n753_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n460_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n743_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n770_), .A2(KEYINPUT119), .A3(new_n747_), .A4(new_n752_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n768_), .A2(new_n534_), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n762_), .B1(new_n772_), .B2(new_n758_), .ZN(new_n773_));
  OAI211_X1 g572(.A(new_n764_), .B(new_n766_), .C1(new_n773_), .C2(new_n760_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT120), .ZN(new_n775_));
  AOI211_X1 g574(.A(new_n775_), .B(G113gat), .C1(new_n773_), .C2(new_n518_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n772_), .A2(new_n758_), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n777_), .A2(new_n518_), .A3(new_n763_), .ZN(new_n778_));
  AOI21_X1  g577(.A(KEYINPUT120), .B1(new_n778_), .B2(new_n765_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n774_), .B1(new_n776_), .B2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT121), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  OAI211_X1 g581(.A(KEYINPUT121), .B(new_n774_), .C1(new_n776_), .C2(new_n779_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1340gat));
  XNOR2_X1  g583(.A(KEYINPUT122), .B(G120gat), .ZN(new_n785_));
  INV_X1    g584(.A(new_n773_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n786_), .A2(KEYINPUT59), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n787_), .A2(new_n764_), .ZN(new_n788_));
  OAI21_X1  g587(.A(new_n785_), .B1(new_n788_), .B2(new_n644_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT60), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n785_), .B1(new_n493_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT123), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT123), .B1(new_n785_), .B2(new_n790_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n791_), .B2(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n789_), .B1(new_n786_), .B2(new_n795_), .ZN(G1341gat));
  OAI21_X1  g595(.A(G127gat), .B1(new_n788_), .B2(new_n534_), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n534_), .A2(G127gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n797_), .B1(new_n786_), .B2(new_n798_), .ZN(G1342gat));
  INV_X1    g598(.A(G134gat), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n800_), .B1(new_n786_), .B2(new_n460_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT124), .ZN(new_n802_));
  OR2_X1    g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n802_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n788_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n545_), .A2(new_n800_), .ZN(new_n806_));
  AOI22_X1  g605(.A1(new_n803_), .A2(new_n804_), .B1(new_n805_), .B2(new_n806_), .ZN(G1343gat));
  AOI21_X1  g606(.A(new_n283_), .B1(new_n772_), .B2(new_n758_), .ZN(new_n808_));
  NAND4_X1  g607(.A1(new_n808_), .A2(new_n540_), .A3(new_n583_), .A4(new_n371_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(new_n519_), .ZN(new_n810_));
  XOR2_X1   g609(.A(new_n810_), .B(G141gat), .Z(G1344gat));
  NOR2_X1   g610(.A1(new_n809_), .A2(new_n644_), .ZN(new_n812_));
  XOR2_X1   g611(.A(new_n812_), .B(G148gat), .Z(G1345gat));
  NOR2_X1   g612(.A1(new_n809_), .A2(new_n534_), .ZN(new_n814_));
  XOR2_X1   g613(.A(KEYINPUT61), .B(G155gat), .Z(new_n815_));
  XNOR2_X1  g614(.A(new_n814_), .B(new_n815_), .ZN(G1346gat));
  OAI21_X1  g615(.A(G162gat), .B1(new_n809_), .B2(new_n545_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n460_), .A2(G162gat), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n817_), .B1(new_n809_), .B2(new_n818_), .ZN(G1347gat));
  NOR3_X1   g618(.A1(new_n583_), .A2(new_n371_), .A3(new_n284_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n759_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT125), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n759_), .A2(KEYINPUT125), .A3(new_n820_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  XOR2_X1   g624(.A(KEYINPUT22), .B(G169gat), .Z(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n825_), .A2(new_n518_), .A3(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT62), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n759_), .A2(new_n518_), .A3(new_n820_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(G169gat), .ZN(new_n831_));
  AND3_X1   g630(.A1(new_n830_), .A2(new_n829_), .A3(G169gat), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n828_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n833_), .A2(KEYINPUT126), .ZN(new_n834_));
  INV_X1    g633(.A(KEYINPUT126), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n828_), .B(new_n835_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(G1348gat));
  AOI21_X1  g636(.A(G176gat), .B1(new_n825_), .B2(new_n493_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n777_), .A2(new_n820_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n644_), .A2(new_n257_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n838_), .B1(new_n839_), .B2(new_n840_), .ZN(G1349gat));
  AOI21_X1  g640(.A(G183gat), .B1(new_n839_), .B2(new_n535_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n534_), .A2(new_n265_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n825_), .B2(new_n843_), .ZN(G1350gat));
  NAND3_X1  g643(.A1(new_n825_), .A2(new_n261_), .A3(new_n602_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n545_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n846_));
  INV_X1    g645(.A(G190gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n845_), .B1(new_n846_), .B2(new_n847_), .ZN(G1351gat));
  NOR3_X1   g647(.A1(new_n584_), .A2(new_n540_), .A3(new_n371_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n808_), .A2(new_n849_), .ZN(new_n850_));
  OR4_X1    g649(.A1(KEYINPUT127), .A2(new_n850_), .A3(new_n289_), .A4(new_n519_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n289_), .B1(new_n850_), .B2(new_n519_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n808_), .A2(new_n849_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n853_), .A2(G197gat), .A3(new_n518_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT127), .ZN(new_n855_));
  AND3_X1   g654(.A1(new_n851_), .A2(new_n852_), .A3(new_n855_), .ZN(G1352gat));
  NOR2_X1   g655(.A1(new_n850_), .A2(new_n644_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(new_n290_), .ZN(G1353gat));
  AOI21_X1  g657(.A(new_n534_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n853_), .A2(new_n859_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n861_));
  XOR2_X1   g660(.A(new_n860_), .B(new_n861_), .Z(G1354gat));
  OAI21_X1  g661(.A(G218gat), .B1(new_n850_), .B2(new_n545_), .ZN(new_n863_));
  OR2_X1    g662(.A1(new_n460_), .A2(G218gat), .ZN(new_n864_));
  OAI21_X1  g663(.A(new_n863_), .B1(new_n850_), .B2(new_n864_), .ZN(G1355gat));
endmodule


