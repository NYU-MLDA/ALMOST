//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:55 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n594_, new_n595_, new_n596_, new_n597_, new_n598_, new_n599_,
    new_n600_, new_n601_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n711_, new_n712_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n849_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n889_, new_n890_, new_n891_, new_n893_, new_n894_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n905_, new_n906_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT13), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT69), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT67), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  NOR3_X1   g006(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n205_), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT7), .ZN(new_n212_));
  INV_X1    g011(.A(G99gat), .ZN(new_n213_));
  INV_X1    g012(.A(G106gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(KEYINPUT67), .A3(new_n206_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n209_), .A2(new_n211_), .A3(new_n216_), .ZN(new_n217_));
  XOR2_X1   g016(.A(G85gat), .B(G92gat), .Z(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(KEYINPUT68), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT8), .ZN(new_n220_));
  AOI21_X1  g019(.A(KEYINPUT68), .B1(new_n217_), .B2(new_n218_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n204_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n217_), .A2(new_n218_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n225_), .A2(KEYINPUT69), .A3(KEYINPUT8), .A4(new_n219_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n211_), .A2(new_n215_), .A3(new_n206_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT8), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n227_), .A2(new_n228_), .A3(new_n218_), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n222_), .A2(new_n226_), .A3(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(new_n231_), .B(KEYINPUT65), .ZN(new_n232_));
  INV_X1    g031(.A(G85gat), .ZN(new_n233_));
  INV_X1    g032(.A(G92gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NOR2_X1   g034(.A1(new_n233_), .A2(new_n234_), .ZN(new_n236_));
  XOR2_X1   g035(.A(KEYINPUT64), .B(KEYINPUT9), .Z(new_n237_));
  OAI211_X1 g036(.A(new_n232_), .B(new_n235_), .C1(new_n236_), .C2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n239_));
  XNOR2_X1  g038(.A(new_n238_), .B(new_n239_), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT10), .B(G99gat), .Z(new_n241_));
  INV_X1    g040(.A(new_n241_), .ZN(new_n242_));
  OAI211_X1 g041(.A(new_n240_), .B(new_n211_), .C1(G106gat), .C2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n230_), .A2(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G57gat), .B(G64gat), .ZN(new_n245_));
  OR2_X1    g044(.A1(new_n245_), .A2(KEYINPUT11), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n245_), .A2(KEYINPUT11), .ZN(new_n247_));
  XOR2_X1   g046(.A(G71gat), .B(G78gat), .Z(new_n248_));
  NAND3_X1  g047(.A1(new_n246_), .A2(new_n247_), .A3(new_n248_), .ZN(new_n249_));
  OR2_X1    g048(.A1(new_n247_), .A2(new_n248_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n244_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(KEYINPUT12), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT12), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n244_), .A2(new_n255_), .A3(new_n252_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n254_), .A2(new_n256_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n230_), .A2(new_n243_), .A3(new_n251_), .ZN(new_n258_));
  INV_X1    g057(.A(G230gat), .ZN(new_n259_));
  INV_X1    g058(.A(G233gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(KEYINPUT71), .B1(new_n258_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n258_), .A2(KEYINPUT71), .A3(new_n262_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n257_), .A2(new_n264_), .A3(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n258_), .A2(KEYINPUT70), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n268_));
  NAND4_X1  g067(.A1(new_n230_), .A2(new_n268_), .A3(new_n243_), .A4(new_n251_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n267_), .A2(new_n253_), .A3(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n261_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G120gat), .B(G148gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT5), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G176gat), .B(G204gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n266_), .A2(new_n271_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n276_), .B1(new_n266_), .B2(new_n271_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n203_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n266_), .A2(new_n271_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n281_), .A2(new_n275_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n282_), .A2(KEYINPUT13), .A3(new_n277_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT72), .B1(new_n280_), .B2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n280_), .A2(KEYINPUT72), .A3(new_n283_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G15gat), .B(G22gat), .ZN(new_n288_));
  INV_X1    g087(.A(G8gat), .ZN(new_n289_));
  OAI21_X1  g088(.A(KEYINPUT14), .B1(new_n202_), .B2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n288_), .A2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G1gat), .B(G8gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(G29gat), .B(G36gat), .Z(new_n295_));
  XOR2_X1   g094(.A(G43gat), .B(G50gat), .Z(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n294_), .A2(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n297_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n299_), .A2(new_n293_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n301_), .B(KEYINPUT78), .Z(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(G229gat), .A3(G233gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n297_), .B(KEYINPUT15), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(new_n293_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G229gat), .A2(G233gat), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n306_), .B(KEYINPUT79), .Z(new_n307_));
  NAND3_X1  g106(.A1(new_n305_), .A2(new_n298_), .A3(new_n307_), .ZN(new_n308_));
  AND2_X1   g107(.A1(new_n303_), .A2(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(G113gat), .B(G141gat), .Z(new_n310_));
  XNOR2_X1  g109(.A(G169gat), .B(G197gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n309_), .B(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n287_), .A2(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n251_), .B(new_n293_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(G231gat), .A2(G233gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G127gat), .B(G155gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n319_), .B(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G183gat), .B(G211gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n321_), .B(new_n322_), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n323_), .A2(KEYINPUT17), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n323_), .A2(KEYINPUT17), .ZN(new_n325_));
  OAI21_X1  g124(.A(new_n318_), .B1(new_n324_), .B2(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n326_), .B1(new_n324_), .B2(new_n318_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT77), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n330_));
  XOR2_X1   g129(.A(new_n330_), .B(KEYINPUT86), .Z(new_n331_));
  NOR2_X1   g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT3), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G141gat), .A2(G148gat), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT2), .ZN(new_n335_));
  AOI22_X1  g134(.A1(new_n332_), .A2(new_n333_), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  OAI21_X1  g135(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  OAI21_X1  g137(.A(KEYINPUT87), .B1(new_n331_), .B2(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n330_), .B(KEYINPUT86), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT87), .ZN(new_n341_));
  NAND4_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(new_n337_), .A4(new_n336_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G155gat), .B(G162gat), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT88), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n343_), .B(new_n344_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n339_), .A2(new_n342_), .A3(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT29), .ZN(new_n347_));
  INV_X1    g146(.A(new_n334_), .ZN(new_n348_));
  NOR2_X1   g147(.A1(new_n348_), .A2(new_n332_), .ZN(new_n349_));
  NAND3_X1  g148(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n350_));
  OAI211_X1 g149(.A(new_n349_), .B(new_n350_), .C1(new_n343_), .C2(KEYINPUT1), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n346_), .A2(new_n347_), .A3(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(KEYINPUT28), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G22gat), .B(G50gat), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  OR2_X1    g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  XOR2_X1   g155(.A(G197gat), .B(G204gat), .Z(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT21), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G211gat), .B(G218gat), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G197gat), .B(G204gat), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT21), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n358_), .A2(KEYINPUT89), .A3(new_n359_), .A4(new_n362_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n358_), .A2(new_n359_), .A3(new_n362_), .ZN(new_n364_));
  INV_X1    g163(.A(KEYINPUT89), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n365_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n363_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n342_), .A2(new_n345_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n338_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n341_), .B1(new_n369_), .B2(new_n340_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n351_), .B1(new_n368_), .B2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n367_), .B1(new_n371_), .B2(KEYINPUT29), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G228gat), .A2(G233gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n373_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n347_), .B1(new_n346_), .B2(new_n351_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n375_), .B1(new_n376_), .B2(new_n367_), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G78gat), .B(G106gat), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n353_), .A2(new_n355_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n356_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n372_), .A2(new_n373_), .ZN(new_n383_));
  NOR3_X1   g182(.A1(new_n376_), .A2(new_n367_), .A3(new_n375_), .ZN(new_n384_));
  NOR3_X1   g183(.A1(new_n383_), .A2(new_n384_), .A3(KEYINPUT90), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT90), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n386_), .B1(new_n374_), .B2(new_n377_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n378_), .B1(new_n385_), .B2(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(KEYINPUT91), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT90), .B1(new_n383_), .B2(new_n384_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n374_), .A2(new_n377_), .A3(new_n386_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT91), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n393_), .A3(new_n378_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n382_), .B1(new_n389_), .B2(new_n394_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n356_), .A2(new_n381_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n378_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(new_n380_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n395_), .A2(new_n400_), .ZN(new_n401_));
  XOR2_X1   g200(.A(G127gat), .B(G134gat), .Z(new_n402_));
  XOR2_X1   g201(.A(G113gat), .B(G120gat), .Z(new_n403_));
  XOR2_X1   g202(.A(new_n402_), .B(new_n403_), .Z(new_n404_));
  NAND2_X1  g203(.A1(new_n371_), .A2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(new_n404_), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n346_), .A2(new_n406_), .A3(new_n351_), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n405_), .A2(KEYINPUT4), .A3(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409_));
  XOR2_X1   g208(.A(new_n409_), .B(KEYINPUT94), .Z(new_n410_));
  XOR2_X1   g209(.A(new_n410_), .B(KEYINPUT95), .Z(new_n411_));
  OAI211_X1 g210(.A(new_n408_), .B(new_n411_), .C1(KEYINPUT4), .C2(new_n405_), .ZN(new_n412_));
  AND2_X1   g211(.A1(new_n405_), .A2(new_n407_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(new_n410_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(new_n233_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT0), .B(G57gat), .ZN(new_n417_));
  XNOR2_X1  g216(.A(new_n416_), .B(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n412_), .A2(new_n414_), .A3(new_n418_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n418_), .B1(new_n412_), .B2(new_n414_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G226gat), .A2(G233gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT19), .ZN(new_n424_));
  NAND2_X1  g223(.A1(G183gat), .A2(G190gat), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT23), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(G183gat), .A2(G190gat), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT93), .ZN(new_n430_));
  XNOR2_X1  g229(.A(KEYINPUT22), .B(G169gat), .ZN(new_n431_));
  INV_X1    g230(.A(G176gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(G169gat), .A2(G176gat), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n429_), .B1(new_n430_), .B2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n433_), .A2(KEYINPUT93), .A3(new_n434_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n425_), .A2(KEYINPUT23), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n426_), .A2(G183gat), .A3(G190gat), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT24), .ZN(new_n440_));
  NOR2_X1   g239(.A1(G169gat), .A2(G176gat), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n438_), .A2(new_n439_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT92), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(KEYINPUT26), .B(G190gat), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT25), .B(G183gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n441_), .A2(KEYINPUT81), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT81), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n449_), .B1(G169gat), .B2(G176gat), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n448_), .A2(new_n450_), .A3(KEYINPUT24), .A4(new_n434_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n447_), .A2(new_n451_), .ZN(new_n452_));
  AOI22_X1  g251(.A1(new_n436_), .A2(new_n437_), .B1(new_n444_), .B2(new_n452_), .ZN(new_n453_));
  OAI21_X1  g252(.A(KEYINPUT20), .B1(new_n453_), .B2(new_n367_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n429_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT83), .ZN(new_n456_));
  NOR2_X1   g255(.A1(new_n431_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT22), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n456_), .B1(new_n458_), .B2(G169gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(new_n432_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n455_), .B(new_n434_), .C1(new_n457_), .C2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT80), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT25), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n462_), .A2(new_n463_), .A3(G183gat), .ZN(new_n464_));
  INV_X1    g263(.A(G183gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT25), .B1(new_n465_), .B2(KEYINPUT80), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n445_), .A2(new_n464_), .A3(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n467_), .A2(new_n451_), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT82), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n467_), .A2(new_n451_), .A3(KEYINPUT82), .ZN(new_n471_));
  AOI21_X1  g270(.A(KEYINPUT24), .B1(new_n448_), .B2(new_n450_), .ZN(new_n472_));
  NOR2_X1   g271(.A1(new_n472_), .A2(new_n427_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(new_n471_), .A3(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n367_), .A2(new_n461_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n424_), .B1(new_n454_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT20), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n478_), .B1(new_n453_), .B2(new_n367_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n424_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n461_), .A2(new_n474_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n367_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n479_), .A2(new_n480_), .A3(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n477_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G8gat), .B(G36gat), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n486_), .B(KEYINPUT18), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G64gat), .B(G92gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n487_), .B(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n489_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n477_), .A2(new_n491_), .A3(new_n484_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n490_), .A2(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n492_), .A2(KEYINPUT27), .ZN(new_n494_));
  NOR3_X1   g293(.A1(new_n454_), .A2(new_n476_), .A3(new_n424_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n480_), .B1(new_n479_), .B2(new_n483_), .ZN(new_n496_));
  OAI21_X1  g295(.A(new_n489_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n497_));
  AOI22_X1  g296(.A1(new_n422_), .A2(new_n493_), .B1(new_n494_), .B2(new_n497_), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT30), .ZN(new_n499_));
  XNOR2_X1  g298(.A(new_n481_), .B(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(KEYINPUT85), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G227gat), .A2(G233gat), .ZN(new_n503_));
  INV_X1    g302(.A(G71gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(new_n505_), .B(G99gat), .ZN(new_n506_));
  XOR2_X1   g305(.A(G15gat), .B(G43gat), .Z(new_n507_));
  XNOR2_X1  g306(.A(new_n507_), .B(KEYINPUT84), .ZN(new_n508_));
  XOR2_X1   g307(.A(new_n506_), .B(new_n508_), .Z(new_n509_));
  NAND2_X1  g308(.A1(new_n502_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(new_n404_), .B(KEYINPUT31), .ZN(new_n511_));
  OR2_X1    g310(.A1(new_n500_), .A2(new_n501_), .ZN(new_n512_));
  AND2_X1   g311(.A1(new_n512_), .A2(new_n502_), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n510_), .B(new_n511_), .C1(new_n513_), .C2(new_n509_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n511_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n509_), .B1(new_n512_), .B2(new_n502_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n510_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n515_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n514_), .A2(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n401_), .A2(new_n421_), .A3(new_n498_), .A4(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n493_), .A2(new_n422_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n494_), .A2(new_n497_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n396_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n393_), .B1(new_n392_), .B2(new_n378_), .ZN(new_n525_));
  AOI211_X1 g324(.A(KEYINPUT91), .B(new_n379_), .C1(new_n390_), .C2(new_n391_), .ZN(new_n526_));
  OAI211_X1 g325(.A(new_n380_), .B(new_n524_), .C1(new_n525_), .C2(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n523_), .B1(new_n527_), .B2(new_n399_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n412_), .A2(new_n414_), .A3(new_n418_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT33), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n418_), .B1(new_n413_), .B2(new_n411_), .ZN(new_n532_));
  OAI211_X1 g331(.A(new_n408_), .B(new_n410_), .C1(KEYINPUT4), .C2(new_n405_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND4_X1  g333(.A1(new_n531_), .A2(new_n534_), .A3(new_n492_), .A4(new_n490_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n529_), .A2(new_n530_), .ZN(new_n536_));
  AND2_X1   g335(.A1(new_n491_), .A2(KEYINPUT32), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n537_), .B1(new_n495_), .B2(new_n496_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n485_), .B2(new_n537_), .ZN(new_n539_));
  OAI22_X1  g338(.A1(new_n535_), .A2(new_n536_), .B1(new_n421_), .B2(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n528_), .A2(new_n421_), .B1(new_n401_), .B2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(new_n520_), .B1(new_n541_), .B2(new_n519_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n304_), .B1(new_n230_), .B2(new_n243_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n230_), .A2(new_n299_), .A3(new_n243_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G232gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT34), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n547_), .A2(KEYINPUT35), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n544_), .A2(new_n545_), .A3(new_n548_), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n547_), .A2(KEYINPUT35), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n545_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n551_), .B1(new_n552_), .B2(new_n543_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT74), .ZN(new_n554_));
  OAI21_X1  g353(.A(new_n549_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT36), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G190gat), .B(G218gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT73), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G134gat), .B(G162gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n559_), .B(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n553_), .A2(new_n554_), .ZN(new_n562_));
  NAND4_X1  g361(.A1(new_n556_), .A2(new_n557_), .A3(new_n561_), .A4(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n557_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n561_), .A2(new_n557_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n562_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n564_), .B(new_n565_), .C1(new_n566_), .C2(new_n555_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n563_), .A2(new_n567_), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n542_), .A2(new_n568_), .ZN(new_n569_));
  AND3_X1   g368(.A1(new_n315_), .A2(new_n329_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n421_), .ZN(new_n571_));
  AOI21_X1  g370(.A(new_n202_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(KEYINPUT75), .B(KEYINPUT37), .Z(new_n573_));
  AND3_X1   g372(.A1(new_n563_), .A2(new_n573_), .A3(new_n567_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n563_), .B2(new_n567_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n577_), .A2(new_n328_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n315_), .A2(new_n578_), .A3(new_n542_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n579_), .A2(G1gat), .A3(new_n421_), .ZN(new_n580_));
  AOI21_X1  g379(.A(new_n572_), .B1(KEYINPUT38), .B2(new_n580_), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(KEYINPUT38), .ZN(new_n582_));
  AND2_X1   g381(.A1(new_n582_), .A2(KEYINPUT96), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(KEYINPUT96), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n581_), .B1(new_n583_), .B2(new_n584_), .ZN(G1324gat));
  AOI21_X1  g384(.A(new_n289_), .B1(new_n570_), .B2(new_n523_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(KEYINPUT97), .B(KEYINPUT39), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n586_), .B(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n579_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n289_), .A3(new_n523_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n588_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT40), .ZN(new_n592_));
  XNOR2_X1  g391(.A(new_n591_), .B(new_n592_), .ZN(G1325gat));
  AND2_X1   g392(.A1(new_n570_), .A2(new_n519_), .ZN(new_n594_));
  INV_X1    g393(.A(G15gat), .ZN(new_n595_));
  OR3_X1    g394(.A1(new_n594_), .A2(KEYINPUT98), .A3(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(KEYINPUT98), .B1(new_n594_), .B2(new_n595_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n596_), .A2(KEYINPUT41), .A3(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n589_), .A2(new_n595_), .A3(new_n519_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AOI21_X1  g399(.A(KEYINPUT41), .B1(new_n596_), .B2(new_n597_), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n600_), .A2(new_n601_), .ZN(G1326gat));
  INV_X1    g401(.A(G22gat), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n527_), .A2(new_n399_), .ZN(new_n604_));
  AOI21_X1  g403(.A(new_n603_), .B1(new_n570_), .B2(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(KEYINPUT99), .B(KEYINPUT42), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n589_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n607_), .A2(new_n608_), .ZN(G1327gat));
  NOR2_X1   g408(.A1(new_n568_), .A2(new_n329_), .ZN(new_n610_));
  AND3_X1   g409(.A1(new_n315_), .A2(new_n542_), .A3(new_n610_), .ZN(new_n611_));
  AOI21_X1  g410(.A(G29gat), .B1(new_n611_), .B2(new_n571_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT100), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT43), .ZN(new_n614_));
  OAI211_X1 g413(.A(new_n542_), .B(new_n577_), .C1(new_n613_), .C2(new_n614_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n531_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n490_), .A2(new_n534_), .A3(new_n492_), .ZN(new_n617_));
  NOR3_X1   g416(.A1(new_n616_), .A2(new_n617_), .A3(new_n536_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n421_), .A2(new_n539_), .ZN(new_n619_));
  OAI211_X1 g418(.A(new_n399_), .B(new_n527_), .C1(new_n618_), .C2(new_n619_), .ZN(new_n620_));
  OAI211_X1 g419(.A(new_n421_), .B(new_n498_), .C1(new_n395_), .C2(new_n400_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n519_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n519_), .A2(new_n421_), .ZN(new_n623_));
  NOR3_X1   g422(.A1(new_n623_), .A2(new_n604_), .A3(new_n523_), .ZN(new_n624_));
  OAI22_X1  g423(.A1(new_n622_), .A2(new_n624_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n625_));
  OAI21_X1  g424(.A(new_n613_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n625_), .A2(KEYINPUT43), .A3(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n615_), .A2(new_n627_), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n285_), .A2(new_n328_), .A3(new_n286_), .A4(new_n313_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT44), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n631_), .A2(KEYINPUT101), .A3(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT101), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n629_), .B1(new_n615_), .B2(new_n627_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n634_), .B1(new_n635_), .B2(KEYINPUT44), .ZN(new_n636_));
  AOI22_X1  g435(.A1(new_n633_), .A2(new_n636_), .B1(KEYINPUT44), .B2(new_n635_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n571_), .A2(G29gat), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n612_), .B1(new_n637_), .B2(new_n638_), .ZN(G1328gat));
  INV_X1    g438(.A(G36gat), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n611_), .A2(new_n640_), .A3(new_n523_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT45), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n633_), .A2(new_n636_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n498_), .B1(new_n635_), .B2(KEYINPUT44), .ZN(new_n644_));
  AOI211_X1 g443(.A(KEYINPUT102), .B(new_n640_), .C1(new_n643_), .C2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n646_));
  AOI21_X1  g445(.A(KEYINPUT101), .B1(new_n631_), .B2(new_n632_), .ZN(new_n647_));
  NOR3_X1   g446(.A1(new_n635_), .A2(new_n634_), .A3(KEYINPUT44), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n644_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n646_), .B1(new_n649_), .B2(G36gat), .ZN(new_n650_));
  OAI21_X1  g449(.A(new_n642_), .B1(new_n645_), .B2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT46), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  OAI211_X1 g452(.A(KEYINPUT46), .B(new_n642_), .C1(new_n645_), .C2(new_n650_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(G1329gat));
  AND3_X1   g454(.A1(new_n637_), .A2(G43gat), .A3(new_n519_), .ZN(new_n656_));
  AOI21_X1  g455(.A(G43gat), .B1(new_n611_), .B2(new_n519_), .ZN(new_n657_));
  OR3_X1    g456(.A1(new_n656_), .A2(KEYINPUT47), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(KEYINPUT47), .B1(new_n656_), .B2(new_n657_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(G1330gat));
  INV_X1    g459(.A(G50gat), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n611_), .A2(new_n661_), .A3(new_n604_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n637_), .A2(new_n604_), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n662_), .B1(new_n663_), .B2(new_n661_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(KEYINPUT103), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT103), .ZN(new_n666_));
  OAI211_X1 g465(.A(new_n666_), .B(new_n662_), .C1(new_n663_), .C2(new_n661_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1331gat));
  AND2_X1   g467(.A1(new_n542_), .A2(new_n314_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n578_), .A2(new_n287_), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n669_), .B1(new_n670_), .B2(KEYINPUT104), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n671_), .B1(KEYINPUT104), .B2(new_n670_), .ZN(new_n672_));
  INV_X1    g471(.A(G57gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n672_), .A2(new_n673_), .A3(new_n571_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n313_), .A2(new_n328_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n569_), .A2(new_n287_), .A3(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT105), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(new_n571_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n674_), .B1(new_n673_), .B2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT106), .ZN(G1332gat));
  INV_X1    g479(.A(G64gat), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n672_), .A2(new_n681_), .A3(new_n523_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n677_), .A2(new_n523_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n683_), .A2(G64gat), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n683_), .B2(G64gat), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n682_), .B1(new_n685_), .B2(new_n686_), .ZN(G1333gat));
  NAND2_X1  g486(.A1(new_n519_), .A2(new_n504_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT108), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n672_), .A2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n677_), .A2(new_n519_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G71gat), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n692_), .A2(KEYINPUT49), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n692_), .A2(KEYINPUT49), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n690_), .B1(new_n693_), .B2(new_n694_), .ZN(G1334gat));
  INV_X1    g494(.A(G78gat), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n672_), .A2(new_n696_), .A3(new_n604_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n677_), .A2(new_n604_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G78gat), .ZN(new_n699_));
  AND2_X1   g498(.A1(new_n699_), .A2(KEYINPUT50), .ZN(new_n700_));
  NOR2_X1   g499(.A1(new_n699_), .A2(KEYINPUT50), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n697_), .B1(new_n700_), .B2(new_n701_), .ZN(G1335gat));
  NAND3_X1  g501(.A1(new_n669_), .A2(new_n287_), .A3(new_n610_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(G85gat), .B1(new_n704_), .B2(new_n571_), .ZN(new_n705_));
  AOI211_X1 g504(.A(new_n329_), .B(new_n313_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n628_), .A2(new_n706_), .ZN(new_n707_));
  XOR2_X1   g506(.A(new_n707_), .B(KEYINPUT109), .Z(new_n708_));
  NOR2_X1   g507(.A1(new_n421_), .A2(new_n233_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n705_), .B1(new_n708_), .B2(new_n709_), .ZN(G1336gat));
  AOI21_X1  g509(.A(G92gat), .B1(new_n704_), .B2(new_n523_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n498_), .A2(new_n234_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n711_), .B1(new_n708_), .B2(new_n712_), .ZN(G1337gat));
  AOI21_X1  g512(.A(new_n213_), .B1(new_n707_), .B2(new_n519_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n519_), .ZN(new_n715_));
  NOR3_X1   g514(.A1(new_n703_), .A2(new_n242_), .A3(new_n715_), .ZN(new_n716_));
  OR3_X1    g515(.A1(new_n714_), .A2(KEYINPUT111), .A3(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(KEYINPUT111), .B1(new_n714_), .B2(new_n716_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT51), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n720_), .A2(KEYINPUT110), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n719_), .B(new_n721_), .ZN(G1338gat));
  NAND4_X1  g521(.A1(new_n628_), .A2(KEYINPUT112), .A3(new_n604_), .A4(new_n706_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(G106gat), .ZN(new_n724_));
  INV_X1    g523(.A(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT52), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n707_), .A2(new_n604_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n725_), .B(new_n726_), .C1(new_n727_), .C2(KEYINPUT112), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT112), .B1(new_n707_), .B2(new_n604_), .ZN(new_n729_));
  OAI21_X1  g528(.A(KEYINPUT52), .B1(new_n729_), .B2(new_n724_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n728_), .A2(new_n730_), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n704_), .A2(new_n214_), .A3(new_n604_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n731_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n733_), .A2(KEYINPUT53), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT53), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n731_), .A2(new_n735_), .A3(new_n732_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n734_), .A2(new_n736_), .ZN(G1339gat));
  NAND3_X1  g536(.A1(new_n280_), .A2(new_n675_), .A3(new_n283_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT113), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  NAND4_X1  g539(.A1(new_n280_), .A2(new_n675_), .A3(new_n283_), .A4(KEYINPUT113), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT54), .ZN(new_n743_));
  AND3_X1   g542(.A1(new_n742_), .A2(new_n743_), .A3(new_n576_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n742_), .B2(new_n576_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n744_), .A2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT116), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n302_), .A2(new_n307_), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n307_), .B1(new_n294_), .B2(new_n297_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n312_), .B1(new_n305_), .B2(new_n749_), .ZN(new_n750_));
  AOI22_X1  g549(.A1(new_n309_), .A2(new_n312_), .B1(new_n748_), .B2(new_n750_), .ZN(new_n751_));
  AND2_X1   g550(.A1(new_n277_), .A2(new_n751_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT115), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n753_), .A2(KEYINPUT58), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n255_), .B1(new_n244_), .B2(new_n252_), .ZN(new_n756_));
  AOI211_X1 g555(.A(KEYINPUT12), .B(new_n251_), .C1(new_n230_), .C2(new_n243_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n267_), .A2(new_n269_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n261_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(KEYINPUT114), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT55), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n265_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(new_n263_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n257_), .A2(new_n264_), .A3(KEYINPUT55), .A4(new_n265_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT114), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n766_), .B(new_n261_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n767_));
  NAND4_X1  g566(.A1(new_n761_), .A2(new_n764_), .A3(new_n765_), .A4(new_n767_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n768_), .A2(KEYINPUT56), .A3(new_n275_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT56), .B1(new_n768_), .B2(new_n275_), .ZN(new_n770_));
  OAI211_X1 g569(.A(new_n752_), .B(new_n755_), .C1(new_n769_), .C2(new_n770_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n771_), .A2(new_n577_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n768_), .A2(new_n275_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT56), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n768_), .A2(KEYINPUT56), .A3(new_n275_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n755_), .B1(new_n777_), .B2(new_n752_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n747_), .B1(new_n772_), .B2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n313_), .A2(new_n277_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n282_), .A2(new_n277_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n751_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n783_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n568_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT57), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n752_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(new_n754_), .ZN(new_n789_));
  NAND4_X1  g588(.A1(new_n789_), .A2(KEYINPUT116), .A3(new_n577_), .A4(new_n771_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n780_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n783_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n793_), .A2(KEYINPUT57), .A3(new_n568_), .ZN(new_n794_));
  NAND4_X1  g593(.A1(new_n779_), .A2(new_n787_), .A3(new_n790_), .A4(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n746_), .B1(new_n795_), .B2(new_n328_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n715_), .A2(new_n421_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n604_), .A2(new_n523_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(KEYINPUT59), .B1(new_n796_), .B2(new_n799_), .ZN(new_n800_));
  NOR2_X1   g599(.A1(new_n799_), .A2(KEYINPUT59), .ZN(new_n801_));
  AOI21_X1  g600(.A(KEYINPUT57), .B1(new_n793_), .B2(new_n568_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n568_), .ZN(new_n803_));
  AOI211_X1 g602(.A(new_n786_), .B(new_n803_), .C1(new_n792_), .C2(new_n783_), .ZN(new_n804_));
  NOR2_X1   g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n789_), .A2(new_n577_), .A3(new_n771_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n329_), .B1(new_n805_), .B2(new_n806_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n801_), .B1(new_n807_), .B2(new_n746_), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n800_), .A2(new_n313_), .A3(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(G113gat), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n795_), .A2(new_n328_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n746_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n799_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  OAI21_X1  g614(.A(KEYINPUT117), .B1(new_n796_), .B2(new_n799_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  OR2_X1    g616(.A1(new_n314_), .A2(G113gat), .ZN(new_n818_));
  OAI21_X1  g617(.A(new_n810_), .B1(new_n817_), .B2(new_n818_), .ZN(G1340gat));
  INV_X1    g618(.A(KEYINPUT59), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n287_), .B(new_n808_), .C1(new_n813_), .C2(new_n820_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n821_), .A2(KEYINPUT119), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT119), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n800_), .A2(new_n823_), .A3(new_n287_), .A4(new_n808_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(G120gat), .A3(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT60), .ZN(new_n826_));
  AOI21_X1  g625(.A(G120gat), .B1(new_n287_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n826_), .A2(G120gat), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n827_), .B1(KEYINPUT118), .B2(new_n828_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n829_), .B1(KEYINPUT118), .B2(new_n827_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n815_), .A2(new_n816_), .A3(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n825_), .A2(new_n831_), .ZN(G1341gat));
  NAND3_X1  g631(.A1(new_n815_), .A2(new_n329_), .A3(new_n816_), .ZN(new_n833_));
  INV_X1    g632(.A(G127gat), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n800_), .A2(new_n808_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n328_), .A2(KEYINPUT120), .ZN(new_n836_));
  MUX2_X1   g635(.A(KEYINPUT120), .B(new_n836_), .S(G127gat), .Z(new_n837_));
  AOI22_X1  g636(.A1(new_n833_), .A2(new_n834_), .B1(new_n835_), .B2(new_n837_), .ZN(G1342gat));
  NAND3_X1  g637(.A1(new_n800_), .A2(new_n577_), .A3(new_n808_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(G134gat), .ZN(new_n840_));
  OR2_X1    g639(.A1(new_n568_), .A2(G134gat), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n840_), .B1(new_n817_), .B2(new_n841_), .ZN(G1343gat));
  NOR2_X1   g641(.A1(new_n796_), .A2(new_n519_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n528_), .A2(new_n571_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n843_), .A2(new_n313_), .A3(new_n845_), .ZN(new_n846_));
  XOR2_X1   g645(.A(KEYINPUT121), .B(G141gat), .Z(new_n847_));
  XNOR2_X1  g646(.A(new_n846_), .B(new_n847_), .ZN(G1344gat));
  NAND3_X1  g647(.A1(new_n843_), .A2(new_n287_), .A3(new_n845_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G148gat), .ZN(G1345gat));
  NAND3_X1  g649(.A1(new_n843_), .A2(new_n329_), .A3(new_n845_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT61), .B(G155gat), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1346gat));
  NOR2_X1   g652(.A1(new_n568_), .A2(G162gat), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n843_), .A2(new_n845_), .A3(new_n854_), .ZN(new_n855_));
  NOR4_X1   g654(.A1(new_n796_), .A2(new_n576_), .A3(new_n519_), .A4(new_n844_), .ZN(new_n856_));
  INV_X1    g655(.A(G162gat), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  OAI211_X1 g659(.A(new_n855_), .B(KEYINPUT122), .C1(new_n857_), .C2(new_n856_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n860_), .A2(new_n861_), .ZN(G1347gat));
  INV_X1    g661(.A(KEYINPUT124), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n498_), .A2(new_n571_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n519_), .ZN(new_n865_));
  NOR2_X1   g664(.A1(new_n865_), .A2(new_n604_), .ZN(new_n866_));
  OAI211_X1 g665(.A(new_n313_), .B(new_n866_), .C1(new_n807_), .C2(new_n746_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n863_), .B1(new_n867_), .B2(G169gat), .ZN(new_n868_));
  XOR2_X1   g667(.A(KEYINPUT123), .B(KEYINPUT62), .Z(new_n869_));
  INV_X1    g668(.A(new_n867_), .ZN(new_n870_));
  AOI22_X1  g669(.A1(new_n868_), .A2(new_n869_), .B1(new_n870_), .B2(new_n431_), .ZN(new_n871_));
  OR2_X1    g670(.A1(new_n868_), .A2(new_n869_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n867_), .A2(new_n863_), .A3(G169gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n872_), .B2(new_n873_), .ZN(G1348gat));
  OAI21_X1  g673(.A(new_n866_), .B1(new_n807_), .B2(new_n746_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(G176gat), .B1(new_n876_), .B2(new_n287_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n796_), .A2(new_n604_), .ZN(new_n878_));
  AOI211_X1 g677(.A(new_n432_), .B(new_n865_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n877_), .B1(new_n878_), .B2(new_n879_), .ZN(G1349gat));
  NOR2_X1   g679(.A1(new_n865_), .A2(new_n328_), .ZN(new_n881_));
  AOI21_X1  g680(.A(G183gat), .B1(new_n878_), .B2(new_n881_), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n875_), .A2(new_n328_), .A3(new_n446_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n882_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT125), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT125), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n886_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(G1350gat));
  OAI21_X1  g687(.A(G190gat), .B1(new_n875_), .B2(new_n576_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n803_), .A2(new_n445_), .ZN(new_n890_));
  XOR2_X1   g689(.A(new_n890_), .B(KEYINPUT126), .Z(new_n891_));
  OAI21_X1  g690(.A(new_n889_), .B1(new_n875_), .B2(new_n891_), .ZN(G1351gat));
  AND2_X1   g691(.A1(new_n604_), .A2(new_n864_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n843_), .A2(new_n313_), .A3(new_n893_), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n894_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g694(.A1(new_n843_), .A2(new_n287_), .A3(new_n893_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g696(.A1(new_n843_), .A2(new_n893_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  XOR2_X1   g698(.A(KEYINPUT63), .B(G211gat), .Z(new_n900_));
  NAND3_X1  g699(.A1(new_n899_), .A2(new_n329_), .A3(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n902_), .B1(new_n898_), .B2(new_n328_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n901_), .A2(new_n903_), .ZN(G1354gat));
  OR3_X1    g703(.A1(new_n898_), .A2(G218gat), .A3(new_n568_), .ZN(new_n905_));
  OAI21_X1  g704(.A(G218gat), .B1(new_n898_), .B2(new_n576_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1355gat));
endmodule


