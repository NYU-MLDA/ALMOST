//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n630_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n828_, new_n829_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n839_, new_n841_,
    new_n842_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n856_,
    new_n858_, new_n860_, new_n861_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n890_, new_n891_, new_n892_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G134gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT83), .B(G127gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT84), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT1), .ZN(new_n213_));
  AND2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n212_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n213_), .A2(G155gat), .A3(G162gat), .ZN(new_n216_));
  XOR2_X1   g015(.A(new_n216_), .B(KEYINPUT85), .Z(new_n217_));
  OAI211_X1 g016(.A(new_n207_), .B(new_n209_), .C1(new_n215_), .C2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(new_n214_), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT88), .ZN(new_n220_));
  AOI22_X1  g019(.A1(new_n220_), .A2(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(KEYINPUT2), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n221_), .B(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT87), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT86), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n224_), .B1(new_n208_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT86), .B1(new_n227_), .B2(KEYINPUT87), .ZN(new_n228_));
  AOI22_X1  g027(.A1(new_n226_), .A2(new_n227_), .B1(new_n208_), .B2(new_n228_), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n219_), .B(new_n212_), .C1(new_n223_), .C2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n218_), .A2(new_n230_), .ZN(new_n231_));
  OAI211_X1 g030(.A(KEYINPUT97), .B(new_n206_), .C1(new_n231_), .C2(KEYINPUT98), .ZN(new_n232_));
  INV_X1    g031(.A(new_n205_), .ZN(new_n233_));
  OR2_X1    g032(.A1(new_n204_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n204_), .A2(new_n233_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n234_), .A2(new_n235_), .A3(KEYINPUT97), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT98), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n236_), .A2(new_n237_), .A3(new_n218_), .A4(new_n230_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n232_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n231_), .A2(new_n206_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT97), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n239_), .A2(KEYINPUT99), .A3(KEYINPUT4), .A4(new_n242_), .ZN(new_n243_));
  INV_X1    g042(.A(KEYINPUT99), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n242_), .A2(new_n238_), .A3(new_n232_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT4), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n243_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G225gat), .A2(G233gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n231_), .A2(new_n246_), .A3(new_n206_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n248_), .A2(new_n250_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n245_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n253_), .A2(new_n249_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(G1gat), .B(G29gat), .ZN(new_n255_));
  INV_X1    g054(.A(G85gat), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n255_), .B(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT0), .B(G57gat), .ZN(new_n258_));
  XOR2_X1   g057(.A(new_n257_), .B(new_n258_), .Z(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n252_), .A2(new_n254_), .A3(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT102), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n252_), .A2(new_n254_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n263_), .A2(new_n259_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT102), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n252_), .A2(new_n265_), .A3(new_n254_), .A4(new_n260_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n262_), .A2(new_n264_), .A3(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(G226gat), .A2(G233gat), .ZN(new_n268_));
  XNOR2_X1  g067(.A(new_n268_), .B(KEYINPUT19), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT20), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT21), .ZN(new_n272_));
  INV_X1    g071(.A(G197gat), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(G204gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT91), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n272_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(G197gat), .B(G204gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n276_), .B(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G211gat), .B(G218gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(new_n280_), .B(KEYINPUT92), .ZN(new_n281_));
  OR3_X1    g080(.A1(new_n279_), .A2(new_n277_), .A3(new_n272_), .ZN(new_n282_));
  XOR2_X1   g081(.A(new_n282_), .B(KEYINPUT93), .Z(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n281_), .A2(new_n284_), .ZN(new_n285_));
  NAND2_X1  g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(KEYINPUT23), .ZN(new_n287_));
  OR2_X1    g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288_));
  AOI22_X1  g087(.A1(new_n287_), .A2(new_n288_), .B1(G169gat), .B2(G176gat), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT22), .B(G169gat), .ZN(new_n290_));
  INV_X1    g089(.A(G176gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n289_), .A2(new_n292_), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT25), .B(G183gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT26), .B(G190gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT24), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G169gat), .A2(G176gat), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n297_), .A2(KEYINPUT24), .A3(new_n299_), .ZN(new_n300_));
  NAND4_X1  g099(.A1(new_n296_), .A2(new_n287_), .A3(new_n298_), .A4(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n293_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n271_), .B1(new_n285_), .B2(new_n302_), .ZN(new_n303_));
  OR2_X1    g102(.A1(new_n280_), .A2(KEYINPUT92), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n280_), .A2(KEYINPUT92), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n283_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n290_), .B(KEYINPUT96), .Z(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n289_), .B1(new_n308_), .B2(G176gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n306_), .A2(new_n301_), .A3(new_n309_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n270_), .B1(new_n303_), .B2(new_n310_), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n301_), .B(KEYINPUT95), .Z(new_n312_));
  NAND2_X1  g111(.A1(new_n312_), .A2(new_n309_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n285_), .A2(new_n313_), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n281_), .A2(new_n293_), .A3(new_n301_), .A4(new_n284_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n314_), .A2(KEYINPUT20), .A3(new_n315_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n316_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n311_), .B1(new_n270_), .B2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(G8gat), .B(G36gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(G92gat), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT18), .B(G64gat), .ZN(new_n321_));
  XOR2_X1   g120(.A(new_n320_), .B(new_n321_), .Z(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT32), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n318_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n316_), .A2(new_n269_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n303_), .B(new_n270_), .C1(new_n285_), .C2(new_n313_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n325_), .A2(new_n326_), .A3(new_n323_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n267_), .A2(new_n324_), .A3(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT33), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n261_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n325_), .A2(new_n326_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n322_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n325_), .A2(new_n326_), .A3(new_n322_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n259_), .B1(new_n245_), .B2(new_n249_), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT100), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n248_), .A2(new_n249_), .A3(new_n251_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND4_X1  g138(.A1(new_n252_), .A2(KEYINPUT33), .A3(new_n254_), .A4(new_n260_), .ZN(new_n340_));
  NAND4_X1  g139(.A1(new_n330_), .A2(new_n335_), .A3(new_n339_), .A4(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT101), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n333_), .A2(new_n334_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n344_), .B1(new_n329_), .B2(new_n261_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n345_), .A2(KEYINPUT101), .A3(new_n339_), .A4(new_n340_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n328_), .A2(new_n343_), .A3(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n231_), .A2(KEYINPUT29), .ZN(new_n348_));
  XOR2_X1   g147(.A(G78gat), .B(G106gat), .Z(new_n349_));
  XNOR2_X1  g148(.A(new_n349_), .B(KEYINPUT90), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G228gat), .A2(G233gat), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n350_), .B(new_n351_), .ZN(new_n352_));
  OR3_X1    g151(.A1(new_n306_), .A2(new_n348_), .A3(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n352_), .B1(new_n306_), .B2(new_n348_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n353_), .A2(new_n354_), .A3(KEYINPUT89), .ZN(new_n355_));
  XNOR2_X1  g154(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n356_));
  OR2_X1    g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  OR2_X1    g156(.A1(new_n231_), .A2(KEYINPUT29), .ZN(new_n358_));
  XNOR2_X1  g157(.A(G22gat), .B(G50gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(new_n356_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n357_), .A2(new_n360_), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n360_), .B1(new_n357_), .B2(new_n361_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  OR2_X1    g164(.A1(new_n302_), .A2(KEYINPUT30), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n302_), .A2(KEYINPUT30), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n366_), .A2(KEYINPUT82), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G227gat), .A2(G233gat), .ZN(new_n369_));
  INV_X1    g168(.A(G71gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(new_n371_), .B(G99gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G15gat), .B(G43gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n372_), .B(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n368_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT31), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT31), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n368_), .A2(new_n377_), .A3(new_n374_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n379_), .A2(new_n206_), .ZN(new_n380_));
  INV_X1    g179(.A(new_n206_), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n376_), .A2(new_n378_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n366_), .A2(new_n367_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT82), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n383_), .A2(new_n386_), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n380_), .A2(new_n385_), .A3(new_n384_), .A4(new_n382_), .ZN(new_n388_));
  AND2_X1   g187(.A1(new_n387_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(new_n365_), .A2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(new_n267_), .ZN(new_n391_));
  OAI211_X1 g190(.A(KEYINPUT27), .B(new_n334_), .C1(new_n318_), .C2(new_n322_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n392_), .B1(new_n335_), .B2(KEYINPUT27), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n389_), .B1(new_n363_), .B2(new_n364_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n364_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n387_), .A2(new_n388_), .ZN(new_n396_));
  NAND3_X1  g195(.A1(new_n395_), .A2(new_n396_), .A3(new_n362_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n393_), .B1(new_n394_), .B2(new_n397_), .ZN(new_n398_));
  AOI22_X1  g197(.A1(new_n347_), .A2(new_n390_), .B1(new_n391_), .B2(new_n398_), .ZN(new_n399_));
  XOR2_X1   g198(.A(G71gat), .B(G78gat), .Z(new_n400_));
  AND2_X1   g199(.A1(G57gat), .A2(G64gat), .ZN(new_n401_));
  NOR2_X1   g200(.A1(G57gat), .A2(G64gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT11), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(G57gat), .ZN(new_n404_));
  INV_X1    g203(.A(G64gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT11), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G57gat), .A2(G64gat), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n400_), .A2(new_n403_), .A3(new_n409_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(G71gat), .B(G78gat), .ZN(new_n411_));
  OAI211_X1 g210(.A(new_n411_), .B(KEYINPUT11), .C1(new_n402_), .C2(new_n401_), .ZN(new_n412_));
  AND3_X1   g211(.A1(new_n410_), .A2(new_n412_), .A3(KEYINPUT68), .ZN(new_n413_));
  AOI21_X1  g212(.A(KEYINPUT68), .B1(new_n410_), .B2(new_n412_), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  XOR2_X1   g214(.A(G85gat), .B(G92gat), .Z(new_n416_));
  XOR2_X1   g215(.A(KEYINPUT10), .B(G99gat), .Z(new_n417_));
  INV_X1    g216(.A(G106gat), .ZN(new_n418_));
  AOI22_X1  g217(.A1(KEYINPUT9), .A2(new_n416_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(KEYINPUT9), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(G85gat), .A3(G92gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT65), .ZN(new_n422_));
  AND3_X1   g221(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G99gat), .A2(G106gat), .ZN(new_n426_));
  INV_X1    g225(.A(KEYINPUT6), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n426_), .A2(new_n427_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n428_), .A2(KEYINPUT65), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n425_), .A2(new_n430_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n419_), .A2(new_n421_), .A3(new_n431_), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT8), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT67), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n428_), .A2(KEYINPUT67), .A3(new_n429_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(G99gat), .A2(G106gat), .ZN(new_n437_));
  AND2_X1   g236(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n438_));
  NOR2_X1   g237(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n437_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  OAI22_X1  g239(.A1(KEYINPUT66), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n435_), .A2(new_n436_), .A3(new_n440_), .A4(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n433_), .B1(new_n442_), .B2(new_n416_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n416_), .A2(new_n433_), .ZN(new_n444_));
  AND2_X1   g243(.A1(new_n440_), .A2(new_n441_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n444_), .B1(new_n445_), .B2(new_n431_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n432_), .B1(new_n443_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n415_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT12), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G230gat), .A2(G233gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT64), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n442_), .A2(new_n416_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(KEYINPUT8), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n445_), .A2(new_n431_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n444_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n413_), .A2(new_n414_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n432_), .A3(new_n459_), .ZN(new_n460_));
  NAND4_X1  g259(.A1(new_n447_), .A2(KEYINPUT12), .A3(new_n412_), .A4(new_n410_), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n450_), .A2(new_n452_), .A3(new_n460_), .A4(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(new_n452_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n459_), .B1(new_n458_), .B2(new_n432_), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n415_), .A2(new_n447_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G120gat), .B(G148gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(G204gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(KEYINPUT5), .B(G176gat), .ZN(new_n469_));
  XOR2_X1   g268(.A(new_n468_), .B(new_n469_), .Z(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n462_), .A2(new_n466_), .A3(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT69), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n471_), .B1(new_n462_), .B2(new_n466_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  AOI211_X1 g275(.A(new_n473_), .B(new_n471_), .C1(new_n462_), .C2(new_n466_), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT13), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT13), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n480_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n479_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G113gat), .B(G141gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G169gat), .B(G197gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT79), .ZN(new_n488_));
  AND2_X1   g287(.A1(G29gat), .A2(G36gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(G29gat), .A2(G36gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(G50gat), .B1(new_n489_), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(G29gat), .ZN(new_n492_));
  INV_X1    g291(.A(G36gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G50gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(G29gat), .A2(G36gat), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT70), .B(G43gat), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n491_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n498_), .B1(new_n491_), .B2(new_n497_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n488_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(new_n498_), .ZN(new_n502_));
  NOR3_X1   g301(.A1(new_n489_), .A2(new_n490_), .A3(G50gat), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n495_), .B1(new_n494_), .B2(new_n496_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n502_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n491_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n505_), .A2(KEYINPUT79), .A3(new_n506_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G15gat), .B(G22gat), .ZN(new_n508_));
  NAND2_X1  g307(.A1(G1gat), .A2(G8gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT14), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(G8gat), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n202_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n509_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n511_), .A2(new_n514_), .ZN(new_n515_));
  AOI22_X1  g314(.A1(new_n508_), .A2(new_n510_), .B1(new_n509_), .B2(new_n513_), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n515_), .A2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n501_), .A2(new_n507_), .A3(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT80), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n501_), .A2(new_n507_), .A3(new_n517_), .A4(KEYINPUT80), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n501_), .A2(new_n507_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n511_), .B(new_n514_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n523_), .A2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n522_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(G229gat), .A2(G233gat), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT15), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n530_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n505_), .A2(KEYINPUT15), .A3(new_n506_), .ZN(new_n532_));
  AND3_X1   g331(.A1(new_n531_), .A2(new_n532_), .A3(new_n524_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n522_), .A2(new_n527_), .A3(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n487_), .B1(new_n529_), .B2(new_n535_), .ZN(new_n536_));
  AOI22_X1  g335(.A1(new_n520_), .A2(new_n521_), .B1(new_n524_), .B2(new_n523_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n535_), .B(new_n487_), .C1(new_n527_), .C2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT81), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT81), .ZN(new_n540_));
  NAND4_X1  g339(.A1(new_n529_), .A2(new_n540_), .A3(new_n535_), .A4(new_n487_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n536_), .B1(new_n539_), .B2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n483_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n399_), .A2(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(G231gat), .A2(G233gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n524_), .B(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n410_), .A2(new_n412_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n547_), .B(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT68), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G127gat), .B(G155gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(G211gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT16), .B(G183gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n550_), .B1(new_n554_), .B2(KEYINPUT17), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  OR2_X1    g355(.A1(new_n549_), .A2(new_n556_), .ZN(new_n557_));
  OR2_X1    g356(.A1(new_n554_), .A2(KEYINPUT17), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n549_), .A2(new_n556_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n557_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n545_), .A2(new_n560_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n531_), .A2(new_n532_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n447_), .ZN(new_n563_));
  OAI221_X1 g362(.A(new_n432_), .B1(new_n499_), .B2(new_n500_), .C1(new_n443_), .C2(new_n446_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(G232gat), .A2(G233gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT34), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT35), .ZN(new_n568_));
  INV_X1    g367(.A(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n565_), .A2(new_n569_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n567_), .A2(KEYINPUT35), .ZN(new_n571_));
  XOR2_X1   g370(.A(new_n568_), .B(KEYINPUT73), .Z(new_n572_));
  NAND4_X1  g371(.A1(new_n563_), .A2(new_n571_), .A3(new_n564_), .A4(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT74), .ZN(new_n574_));
  AND2_X1   g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n573_), .A2(new_n574_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n570_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(G190gat), .B(G218gat), .Z(new_n578_));
  XNOR2_X1  g377(.A(G134gat), .B(G162gat), .ZN(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  XOR2_X1   g379(.A(new_n580_), .B(KEYINPUT36), .Z(new_n581_));
  INV_X1    g380(.A(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n577_), .A2(new_n582_), .ZN(new_n583_));
  XNOR2_X1  g382(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n585_), .B(KEYINPUT72), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n570_), .B(new_n586_), .C1(new_n575_), .C2(new_n576_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n583_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n561_), .A2(new_n589_), .ZN(new_n590_));
  AOI21_X1  g389(.A(new_n202_), .B1(new_n590_), .B2(new_n267_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT103), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT76), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n573_), .A2(new_n574_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n573_), .A2(new_n574_), .ZN(new_n595_));
  AOI22_X1  g394(.A1(new_n594_), .A2(new_n595_), .B1(new_n565_), .B2(new_n569_), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n581_), .B(KEYINPUT75), .Z(new_n597_));
  OAI21_X1  g396(.A(new_n587_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n593_), .B1(new_n598_), .B2(KEYINPUT37), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n593_), .A3(KEYINPUT37), .ZN(new_n601_));
  XNOR2_X1  g400(.A(KEYINPUT77), .B(KEYINPUT37), .ZN(new_n602_));
  OAI211_X1 g401(.A(new_n587_), .B(new_n602_), .C1(new_n596_), .C2(new_n581_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT78), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT78), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n583_), .A2(new_n605_), .A3(new_n587_), .A4(new_n602_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n600_), .A2(new_n601_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n561_), .A2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(new_n202_), .A3(new_n267_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT38), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n592_), .A2(new_n610_), .ZN(G1324gat));
  NAND3_X1  g410(.A1(new_n608_), .A2(new_n512_), .A3(new_n393_), .ZN(new_n612_));
  NAND4_X1  g411(.A1(new_n545_), .A2(new_n588_), .A3(new_n560_), .A4(new_n393_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT39), .ZN(new_n614_));
  AND3_X1   g413(.A1(new_n613_), .A2(new_n614_), .A3(G8gat), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n614_), .B1(new_n613_), .B2(G8gat), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n612_), .B1(new_n615_), .B2(new_n616_), .ZN(new_n617_));
  XOR2_X1   g416(.A(new_n617_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g417(.A1(new_n590_), .A2(new_n389_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(G15gat), .ZN(new_n620_));
  XOR2_X1   g419(.A(new_n620_), .B(KEYINPUT41), .Z(new_n621_));
  NOR4_X1   g420(.A1(new_n561_), .A2(G15gat), .A3(new_n396_), .A4(new_n607_), .ZN(new_n622_));
  XOR2_X1   g421(.A(new_n622_), .B(KEYINPUT104), .Z(new_n623_));
  NAND2_X1  g422(.A1(new_n621_), .A2(new_n623_), .ZN(G1326gat));
  INV_X1    g423(.A(G22gat), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n625_), .B1(new_n590_), .B2(new_n365_), .ZN(new_n626_));
  XOR2_X1   g425(.A(new_n626_), .B(KEYINPUT42), .Z(new_n627_));
  NAND2_X1  g426(.A1(new_n365_), .A2(new_n625_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT105), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n608_), .A2(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n627_), .A2(new_n630_), .ZN(G1327gat));
  INV_X1    g430(.A(new_n560_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n543_), .A2(new_n632_), .ZN(new_n633_));
  NOR3_X1   g432(.A1(new_n399_), .A2(new_n588_), .A3(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(G29gat), .B1(new_n634_), .B2(new_n267_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n347_), .A2(new_n390_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n398_), .A2(new_n391_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT43), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n607_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n604_), .A2(new_n606_), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n598_), .A2(new_n593_), .A3(KEYINPUT37), .ZN(new_n642_));
  OAI21_X1  g441(.A(new_n641_), .B1(new_n599_), .B2(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT43), .B1(new_n399_), .B2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n640_), .A2(new_n644_), .ZN(new_n645_));
  INV_X1    g444(.A(new_n633_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT106), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT44), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n647_), .A2(new_n648_), .A3(new_n649_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n633_), .B1(new_n640_), .B2(new_n644_), .ZN(new_n651_));
  OAI21_X1  g450(.A(KEYINPUT106), .B1(new_n651_), .B2(KEYINPUT44), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n650_), .A2(new_n652_), .ZN(new_n653_));
  AOI211_X1 g452(.A(new_n492_), .B(new_n391_), .C1(new_n651_), .C2(KEYINPUT44), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n635_), .B1(new_n653_), .B2(new_n654_), .ZN(G1328gat));
  INV_X1    g454(.A(KEYINPUT46), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n645_), .A2(KEYINPUT44), .A3(new_n646_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n657_), .A2(new_n393_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n493_), .B1(new_n653_), .B2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n634_), .A2(new_n493_), .A3(new_n393_), .ZN(new_n661_));
  XOR2_X1   g460(.A(KEYINPUT107), .B(KEYINPUT45), .Z(new_n662_));
  XNOR2_X1  g461(.A(new_n661_), .B(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n663_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n656_), .B1(new_n660_), .B2(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n658_), .B1(new_n650_), .B2(new_n652_), .ZN(new_n666_));
  OAI211_X1 g465(.A(KEYINPUT46), .B(new_n663_), .C1(new_n666_), .C2(new_n493_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n665_), .A2(new_n667_), .ZN(G1329gat));
  INV_X1    g467(.A(G43gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n669_), .B1(new_n651_), .B2(KEYINPUT44), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n648_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n671_));
  NOR3_X1   g470(.A1(new_n651_), .A2(KEYINPUT106), .A3(KEYINPUT44), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n389_), .B(new_n670_), .C1(new_n671_), .C2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n634_), .A2(new_n389_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(new_n669_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n673_), .A2(new_n675_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT47), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT47), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n673_), .A2(new_n678_), .A3(new_n675_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n677_), .A2(new_n679_), .ZN(G1330gat));
  NAND3_X1  g479(.A1(new_n634_), .A2(new_n495_), .A3(new_n365_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n365_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n682_), .B1(new_n651_), .B2(KEYINPUT44), .ZN(new_n683_));
  AOI211_X1 g482(.A(KEYINPUT108), .B(new_n495_), .C1(new_n653_), .C2(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n683_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n686_));
  AOI21_X1  g485(.A(new_n685_), .B1(new_n686_), .B2(G50gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n681_), .B1(new_n684_), .B2(new_n687_), .ZN(G1331gat));
  NOR2_X1   g487(.A1(new_n399_), .A2(new_n482_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n536_), .ZN(new_n690_));
  AOI211_X1 g489(.A(new_n528_), .B(new_n533_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n527_), .B1(new_n522_), .B2(new_n525_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n540_), .B1(new_n693_), .B2(new_n487_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n538_), .A2(KEYINPUT81), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n690_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n696_), .A2(new_n632_), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n689_), .A2(new_n643_), .A3(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(G57gat), .B1(new_n698_), .B2(new_n267_), .ZN(new_n699_));
  NAND3_X1  g498(.A1(new_n689_), .A2(new_n588_), .A3(new_n697_), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT109), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(KEYINPUT109), .ZN(new_n702_));
  AND2_X1   g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n391_), .A2(new_n404_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n699_), .B1(new_n703_), .B2(new_n704_), .ZN(G1332gat));
  NAND3_X1  g504(.A1(new_n698_), .A2(new_n405_), .A3(new_n393_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n701_), .A2(new_n393_), .A3(new_n702_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT48), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n707_), .A2(new_n708_), .A3(G64gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n708_), .B1(new_n707_), .B2(G64gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n706_), .B1(new_n709_), .B2(new_n710_), .ZN(G1333gat));
  NAND3_X1  g510(.A1(new_n698_), .A2(new_n370_), .A3(new_n389_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n701_), .A2(new_n389_), .A3(new_n702_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT49), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n713_), .A2(new_n714_), .A3(G71gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n713_), .B2(G71gat), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n712_), .B1(new_n715_), .B2(new_n716_), .ZN(G1334gat));
  INV_X1    g516(.A(G78gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n698_), .A2(new_n718_), .A3(new_n365_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n701_), .A2(new_n365_), .A3(new_n702_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n721_));
  AND3_X1   g520(.A1(new_n720_), .A2(new_n721_), .A3(G78gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n720_), .B2(G78gat), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n719_), .B1(new_n722_), .B2(new_n723_), .ZN(G1335gat));
  NOR3_X1   g523(.A1(new_n482_), .A2(new_n560_), .A3(new_n696_), .ZN(new_n725_));
  AND3_X1   g524(.A1(new_n638_), .A2(new_n589_), .A3(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(G85gat), .B1(new_n726_), .B2(new_n267_), .ZN(new_n727_));
  AND2_X1   g526(.A1(new_n645_), .A2(new_n725_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n391_), .A2(new_n256_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n727_), .B1(new_n728_), .B2(new_n729_), .ZN(G1336gat));
  AOI21_X1  g529(.A(G92gat), .B1(new_n726_), .B2(new_n393_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n393_), .A2(G92gat), .ZN(new_n732_));
  XOR2_X1   g531(.A(new_n732_), .B(KEYINPUT110), .Z(new_n733_));
  AOI21_X1  g532(.A(new_n731_), .B1(new_n728_), .B2(new_n733_), .ZN(G1337gat));
  AND2_X1   g533(.A1(new_n389_), .A2(new_n417_), .ZN(new_n735_));
  AOI21_X1  g534(.A(KEYINPUT111), .B1(new_n726_), .B2(new_n735_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n728_), .A2(new_n389_), .ZN(new_n737_));
  INV_X1    g536(.A(G99gat), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n736_), .B1(new_n737_), .B2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(KEYINPUT112), .B(KEYINPUT51), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  XNOR2_X1  g540(.A(new_n739_), .B(new_n741_), .ZN(G1338gat));
  NAND3_X1  g541(.A1(new_n726_), .A2(new_n418_), .A3(new_n365_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n645_), .A2(new_n365_), .A3(new_n725_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT52), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n744_), .A2(new_n745_), .A3(G106gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n744_), .B2(G106gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g548(.A1(new_n642_), .A2(new_n599_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n604_), .A2(new_n606_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n482_), .B(new_n697_), .C1(new_n750_), .C2(new_n751_), .ZN(new_n752_));
  XOR2_X1   g551(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n752_), .A2(new_n754_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n643_), .A2(new_n482_), .A3(new_n697_), .A4(new_n753_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n696_), .A2(new_n758_), .A3(new_n472_), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n460_), .B(new_n461_), .C1(new_n464_), .C2(KEYINPUT12), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n760_), .A2(new_n463_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n761_), .A2(KEYINPUT55), .A3(new_n462_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n465_), .B1(new_n449_), .B2(new_n448_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT55), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n763_), .A2(new_n764_), .A3(new_n452_), .A4(new_n461_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n762_), .A2(new_n470_), .A3(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n762_), .A2(KEYINPUT56), .A3(new_n470_), .A4(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n472_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT114), .B1(new_n542_), .B2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n759_), .A2(new_n770_), .A3(new_n772_), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n527_), .B(new_n533_), .C1(new_n520_), .C2(new_n521_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n774_), .B1(new_n527_), .B2(new_n526_), .ZN(new_n775_));
  AOI22_X1  g574(.A1(new_n539_), .A2(new_n541_), .B1(new_n486_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n478_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n773_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n778_), .A2(new_n588_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT57), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n770_), .A2(new_n472_), .A3(new_n776_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT58), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n783_), .A2(new_n784_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n770_), .A2(new_n472_), .A3(new_n786_), .A4(new_n776_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n607_), .A2(new_n785_), .A3(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n778_), .A2(KEYINPUT57), .A3(new_n588_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n781_), .A2(new_n788_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n757_), .B1(new_n790_), .B2(new_n632_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n391_), .A2(new_n393_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NOR3_X1   g592(.A1(new_n791_), .A2(new_n394_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT116), .ZN(new_n795_));
  XNOR2_X1  g594(.A(new_n794_), .B(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(G113gat), .B1(new_n796_), .B2(new_n696_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n798_));
  XNOR2_X1  g597(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n790_), .A2(new_n632_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n757_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n394_), .B1(new_n800_), .B2(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n799_), .B1(new_n802_), .B2(new_n792_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(KEYINPUT117), .A2(KEYINPUT59), .ZN(new_n804_));
  NOR4_X1   g603(.A1(new_n791_), .A2(new_n394_), .A3(new_n793_), .A4(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n798_), .B1(new_n803_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n800_), .A2(new_n801_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n394_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n804_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n807_), .A2(new_n808_), .A3(new_n792_), .A4(new_n809_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n810_), .B(KEYINPUT118), .C1(new_n794_), .C2(new_n799_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n542_), .B1(new_n806_), .B2(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n797_), .B1(new_n812_), .B2(G113gat), .ZN(G1340gat));
  INV_X1    g612(.A(G120gat), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n814_), .B1(new_n482_), .B2(KEYINPUT60), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n796_), .B(new_n815_), .C1(KEYINPUT60), .C2(new_n814_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n803_), .A2(new_n805_), .ZN(new_n817_));
  OAI21_X1  g616(.A(G120gat), .B1(new_n817_), .B2(new_n482_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n816_), .A2(new_n818_), .ZN(G1341gat));
  INV_X1    g618(.A(G127gat), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n796_), .A2(new_n820_), .A3(new_n560_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n632_), .B1(new_n806_), .B2(new_n811_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n821_), .B1(new_n822_), .B2(new_n820_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(KEYINPUT119), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT119), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n821_), .B(new_n825_), .C1(new_n822_), .C2(new_n820_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n824_), .A2(new_n826_), .ZN(G1342gat));
  AOI21_X1  g626(.A(G134gat), .B1(new_n796_), .B2(new_n589_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n806_), .A2(new_n811_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n607_), .A2(G134gat), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n830_), .B(KEYINPUT120), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n828_), .B1(new_n829_), .B2(new_n831_), .ZN(G1343gat));
  INV_X1    g631(.A(new_n397_), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n792_), .A2(new_n833_), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT121), .Z(new_n835_));
  NOR2_X1   g634(.A1(new_n835_), .A2(new_n791_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n696_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n483_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g639(.A1(new_n836_), .A2(new_n560_), .ZN(new_n841_));
  XNOR2_X1  g640(.A(KEYINPUT61), .B(G155gat), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n841_), .B(new_n842_), .ZN(G1346gat));
  AOI21_X1  g642(.A(G162gat), .B1(new_n836_), .B2(new_n589_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n607_), .A2(G162gat), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n836_), .B2(new_n845_), .ZN(G1347gat));
  NAND4_X1  g645(.A1(new_n807_), .A2(new_n391_), .A3(new_n808_), .A4(new_n393_), .ZN(new_n847_));
  OR3_X1    g646(.A1(new_n847_), .A2(KEYINPUT122), .A3(new_n542_), .ZN(new_n848_));
  OAI21_X1  g647(.A(KEYINPUT122), .B1(new_n847_), .B2(new_n542_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(G169gat), .A3(new_n849_), .ZN(new_n850_));
  AND2_X1   g649(.A1(new_n850_), .A2(KEYINPUT62), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n850_), .A2(KEYINPUT62), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n542_), .A2(new_n308_), .ZN(new_n853_));
  XNOR2_X1  g652(.A(new_n853_), .B(KEYINPUT123), .ZN(new_n854_));
  OAI22_X1  g653(.A1(new_n851_), .A2(new_n852_), .B1(new_n847_), .B2(new_n854_), .ZN(G1348gat));
  NOR2_X1   g654(.A1(new_n847_), .A2(new_n482_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(new_n291_), .ZN(G1349gat));
  NOR2_X1   g656(.A1(new_n847_), .A2(new_n632_), .ZN(new_n858_));
  MUX2_X1   g657(.A(G183gat), .B(new_n294_), .S(new_n858_), .Z(G1350gat));
  OAI21_X1  g658(.A(G190gat), .B1(new_n847_), .B2(new_n643_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n589_), .A2(new_n295_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n860_), .B1(new_n847_), .B2(new_n861_), .ZN(G1351gat));
  NAND4_X1  g661(.A1(new_n807_), .A2(new_n391_), .A3(new_n833_), .A4(new_n393_), .ZN(new_n863_));
  INV_X1    g662(.A(new_n863_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n864_), .A2(new_n696_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n865_), .A2(new_n866_), .A3(new_n273_), .ZN(new_n867_));
  INV_X1    g666(.A(new_n867_), .ZN(new_n868_));
  NOR2_X1   g667(.A1(new_n865_), .A2(new_n273_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n866_), .B1(new_n865_), .B2(new_n273_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n868_), .A2(new_n869_), .A3(new_n870_), .ZN(G1352gat));
  NAND2_X1  g670(.A1(new_n864_), .A2(new_n483_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT125), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(G204gat), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT125), .B(G204gat), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n872_), .B2(new_n875_), .ZN(G1353gat));
  XOR2_X1   g675(.A(KEYINPUT63), .B(G211gat), .Z(new_n877_));
  NAND3_X1  g676(.A1(new_n864_), .A2(new_n560_), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT126), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n864_), .A2(new_n560_), .ZN(new_n880_));
  NOR2_X1   g679(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(new_n882_));
  OAI211_X1 g681(.A(new_n879_), .B(new_n881_), .C1(new_n863_), .C2(new_n632_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n878_), .B1(new_n882_), .B2(new_n884_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT127), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n878_), .B(KEYINPUT127), .C1(new_n882_), .C2(new_n884_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(G1354gat));
  INV_X1    g688(.A(G218gat), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n863_), .A2(new_n890_), .A3(new_n643_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n864_), .A2(new_n589_), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n891_), .B1(new_n890_), .B2(new_n892_), .ZN(G1355gat));
endmodule


