//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n682_, new_n683_,
    new_n684_, new_n686_, new_n687_, new_n688_, new_n689_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n763_, new_n764_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n773_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n800_, new_n801_, new_n802_,
    new_n804_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n905_, new_n906_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n936_, new_n937_, new_n939_, new_n940_, new_n942_, new_n943_,
    new_n944_, new_n946_, new_n947_, new_n948_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_;
  INV_X1    g000(.A(KEYINPUT13), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT69), .ZN(new_n203_));
  XOR2_X1   g002(.A(G120gat), .B(G148gat), .Z(new_n204_));
  XNOR2_X1  g003(.A(G176gat), .B(G204gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT68), .B(KEYINPUT5), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n206_), .B(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G230gat), .A2(G233gat), .ZN(new_n209_));
  INV_X1    g008(.A(new_n209_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n215_), .A2(KEYINPUT64), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n212_), .A2(new_n214_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT64), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n221_), .A2(KEYINPUT9), .ZN(new_n222_));
  XOR2_X1   g021(.A(G85gat), .B(G92gat), .Z(new_n223_));
  AOI21_X1  g022(.A(new_n222_), .B1(new_n223_), .B2(KEYINPUT9), .ZN(new_n224_));
  XNOR2_X1  g023(.A(KEYINPUT10), .B(G99gat), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n224_), .B1(G106gat), .B2(new_n225_), .ZN(new_n226_));
  OR2_X1    g025(.A1(new_n220_), .A2(new_n226_), .ZN(new_n227_));
  NOR2_X1   g026(.A1(G99gat), .A2(G106gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT7), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n228_), .B(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n223_), .B1(new_n230_), .B2(new_n215_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT8), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n230_), .B1(new_n216_), .B2(new_n219_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n234_), .A2(KEYINPUT8), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(KEYINPUT8), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n223_), .A2(new_n235_), .A3(new_n236_), .ZN(new_n237_));
  OAI21_X1  g036(.A(new_n232_), .B1(new_n233_), .B2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n227_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(G57gat), .B(G64gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n242_));
  XOR2_X1   g041(.A(G71gat), .B(G78gat), .Z(new_n243_));
  OR2_X1    g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n241_), .A2(KEYINPUT11), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n242_), .A2(new_n243_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n244_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n240_), .A2(new_n247_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n248_), .A2(KEYINPUT66), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n240_), .A2(new_n247_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n250_), .B1(new_n248_), .B2(KEYINPUT66), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n210_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT67), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n247_), .B(new_n253_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n254_), .A2(KEYINPUT12), .A3(new_n239_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n250_), .A2(new_n255_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n247_), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT12), .B1(new_n239_), .B2(new_n257_), .ZN(new_n258_));
  NOR3_X1   g057(.A1(new_n256_), .A2(new_n258_), .A3(new_n210_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n259_), .ZN(new_n260_));
  AOI21_X1  g059(.A(new_n208_), .B1(new_n252_), .B2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(new_n261_), .ZN(new_n262_));
  NAND3_X1  g061(.A1(new_n252_), .A2(new_n260_), .A3(new_n208_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n203_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n263_), .ZN(new_n265_));
  NOR3_X1   g064(.A1(new_n265_), .A2(new_n261_), .A3(KEYINPUT69), .ZN(new_n266_));
  OAI21_X1  g065(.A(new_n202_), .B1(new_n264_), .B2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n262_), .A2(new_n203_), .A3(new_n263_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT69), .B1(new_n265_), .B2(new_n261_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(KEYINPUT13), .ZN(new_n270_));
  AND2_X1   g069(.A1(new_n267_), .A2(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G232gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT34), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G29gat), .B(G36gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G43gat), .B(G50gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n227_), .A2(new_n238_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT70), .B(KEYINPUT15), .ZN(new_n279_));
  XNOR2_X1  g078(.A(new_n276_), .B(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n280_), .B1(new_n227_), .B2(new_n238_), .ZN(new_n281_));
  OAI211_X1 g080(.A(KEYINPUT35), .B(new_n273_), .C1(new_n278_), .C2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n280_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n239_), .A2(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n273_), .A2(KEYINPUT35), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n273_), .A2(KEYINPUT35), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n284_), .A2(new_n285_), .A3(new_n286_), .A4(new_n277_), .ZN(new_n287_));
  XNOR2_X1  g086(.A(G190gat), .B(G218gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(G134gat), .B(G162gat), .ZN(new_n289_));
  XOR2_X1   g088(.A(new_n288_), .B(new_n289_), .Z(new_n290_));
  INV_X1    g089(.A(KEYINPUT36), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n290_), .A2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n292_), .B(KEYINPUT71), .Z(new_n293_));
  NAND3_X1  g092(.A1(new_n282_), .A2(new_n287_), .A3(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT72), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND4_X1  g095(.A1(new_n282_), .A2(new_n287_), .A3(KEYINPUT72), .A4(new_n293_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n290_), .B(KEYINPUT36), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  AOI21_X1  g099(.A(new_n300_), .B1(new_n282_), .B2(new_n287_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(KEYINPUT37), .B1(new_n298_), .B2(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT37), .ZN(new_n305_));
  AOI211_X1 g104(.A(new_n305_), .B(new_n301_), .C1(new_n296_), .C2(new_n297_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(KEYINPUT73), .B(G1gat), .Z(new_n309_));
  INV_X1    g108(.A(G8gat), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT14), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G15gat), .B(G22gat), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n311_), .A2(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G1gat), .B(G8gat), .ZN(new_n314_));
  INV_X1    g113(.A(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(G231gat), .A2(G233gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n321_), .A2(new_n254_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n254_), .ZN(new_n323_));
  XOR2_X1   g122(.A(G127gat), .B(G155gat), .Z(new_n324_));
  XNOR2_X1  g123(.A(G183gat), .B(G211gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n324_), .B(new_n325_), .ZN(new_n326_));
  XOR2_X1   g125(.A(KEYINPUT74), .B(KEYINPUT16), .Z(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  NAND4_X1  g127(.A1(new_n322_), .A2(KEYINPUT17), .A3(new_n323_), .A4(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n321_), .A2(new_n247_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n320_), .A2(new_n257_), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n328_), .B(KEYINPUT17), .Z(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n329_), .A2(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n308_), .A2(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n271_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(KEYINPUT79), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT79), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n339_), .A2(G169gat), .A3(G176gat), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n338_), .A2(new_n340_), .A3(KEYINPUT24), .ZN(new_n341_));
  INV_X1    g140(.A(G169gat), .ZN(new_n342_));
  INV_X1    g141(.A(G176gat), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n342_), .A2(new_n343_), .A3(KEYINPUT78), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT78), .ZN(new_n345_));
  OAI21_X1  g144(.A(new_n345_), .B1(G169gat), .B2(G176gat), .ZN(new_n346_));
  AND2_X1   g145(.A1(new_n344_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n341_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(new_n346_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT24), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT23), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(G183gat), .A3(G190gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(G183gat), .A2(G190gat), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(KEYINPUT23), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n349_), .A2(new_n350_), .B1(new_n352_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT26), .ZN(new_n356_));
  OAI21_X1  g155(.A(KEYINPUT76), .B1(new_n356_), .B2(G190gat), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT76), .ZN(new_n358_));
  INV_X1    g157(.A(G190gat), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n358_), .A2(new_n359_), .A3(KEYINPUT26), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n357_), .A2(new_n360_), .ZN(new_n361_));
  OR3_X1    g160(.A1(new_n359_), .A2(KEYINPUT77), .A3(KEYINPUT26), .ZN(new_n362_));
  XNOR2_X1  g161(.A(KEYINPUT25), .B(G183gat), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n356_), .A2(G190gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT77), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n361_), .A2(new_n362_), .A3(new_n363_), .A4(new_n365_), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n348_), .A2(new_n355_), .A3(new_n366_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(G183gat), .A2(G190gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n353_), .A2(KEYINPUT80), .A3(KEYINPUT23), .ZN(new_n369_));
  INV_X1    g168(.A(new_n369_), .ZN(new_n370_));
  AOI21_X1  g169(.A(KEYINPUT80), .B1(new_n353_), .B2(KEYINPUT23), .ZN(new_n371_));
  NOR2_X1   g170(.A1(new_n370_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT81), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n373_), .B1(new_n353_), .B2(KEYINPUT23), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n351_), .A2(KEYINPUT81), .A3(G183gat), .A4(G190gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  AOI21_X1  g175(.A(new_n368_), .B1(new_n372_), .B2(new_n376_), .ZN(new_n377_));
  AND2_X1   g176(.A1(new_n338_), .A2(new_n340_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n342_), .A2(KEYINPUT22), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT22), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n380_), .A2(G169gat), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n381_), .A3(new_n343_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n367_), .B1(new_n377_), .B2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(G71gat), .B(G99gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(new_n385_), .B(G43gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n384_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G113gat), .B(G120gat), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  INV_X1    g188(.A(G134gat), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n390_), .A2(G127gat), .ZN(new_n391_));
  INV_X1    g190(.A(G127gat), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n392_), .A2(G134gat), .ZN(new_n393_));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n391_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n394_), .B1(new_n391_), .B2(new_n393_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n389_), .B1(new_n395_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n391_), .A2(new_n393_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(KEYINPUT82), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n391_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n399_), .A2(new_n400_), .A3(new_n388_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(new_n387_), .B(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(G227gat), .A2(G233gat), .ZN(new_n404_));
  INV_X1    g203(.A(G15gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(KEYINPUT30), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT31), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n403_), .A2(new_n409_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n403_), .A2(new_n409_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G155gat), .ZN(new_n413_));
  INV_X1    g212(.A(G162gat), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n413_), .A2(new_n414_), .A3(KEYINPUT83), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT83), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(G155gat), .B2(G162gat), .ZN(new_n417_));
  NAND2_X1  g216(.A1(G155gat), .A2(G162gat), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n415_), .A2(new_n417_), .A3(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT84), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT84), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n415_), .A2(new_n417_), .A3(new_n421_), .A4(new_n418_), .ZN(new_n422_));
  OR3_X1    g221(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G141gat), .A2(G148gat), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT2), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n424_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n428_));
  NAND4_X1  g227(.A1(new_n423_), .A2(new_n426_), .A3(new_n427_), .A4(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n420_), .A2(new_n422_), .A3(new_n429_), .ZN(new_n430_));
  OR2_X1    g229(.A1(G141gat), .A2(G148gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(new_n418_), .B(KEYINPUT1), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n415_), .A2(new_n417_), .ZN(new_n433_));
  OAI211_X1 g232(.A(new_n431_), .B(new_n424_), .C1(new_n432_), .C2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n430_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n402_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n430_), .A2(new_n401_), .A3(new_n434_), .A4(new_n397_), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n436_), .A2(KEYINPUT4), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT93), .ZN(new_n440_));
  AOI22_X1  g239(.A1(new_n430_), .A2(new_n434_), .B1(new_n401_), .B2(new_n397_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT4), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n440_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n438_), .A2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n436_), .A2(new_n437_), .A3(new_n439_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G1gat), .B(G29gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(KEYINPUT94), .B(KEYINPUT0), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n447_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G57gat), .B(G85gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n449_), .B(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n445_), .A2(new_n451_), .ZN(new_n453_));
  AOI22_X1  g252(.A1(new_n446_), .A2(new_n452_), .B1(new_n453_), .B2(new_n444_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n412_), .A2(new_n454_), .ZN(new_n455_));
  XOR2_X1   g254(.A(G22gat), .B(G50gat), .Z(new_n456_));
  INV_X1    g255(.A(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT29), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n430_), .A2(new_n458_), .A3(new_n434_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT28), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT28), .ZN(new_n462_));
  NAND4_X1  g261(.A1(new_n430_), .A2(new_n462_), .A3(new_n434_), .A4(new_n458_), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n460_), .A2(new_n461_), .A3(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n464_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n461_), .B1(new_n460_), .B2(new_n463_), .ZN(new_n466_));
  OAI21_X1  g265(.A(new_n457_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n460_), .A2(new_n463_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n468_), .A2(KEYINPUT85), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(new_n456_), .A3(new_n464_), .ZN(new_n470_));
  XOR2_X1   g269(.A(G78gat), .B(G106gat), .Z(new_n471_));
  XNOR2_X1  g270(.A(new_n471_), .B(KEYINPUT88), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT89), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n435_), .A2(KEYINPUT29), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n476_));
  INV_X1    g275(.A(G197gat), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n476_), .B1(new_n477_), .B2(G204gat), .ZN(new_n478_));
  INV_X1    g277(.A(G204gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n479_), .A2(KEYINPUT87), .A3(G197gat), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n477_), .A2(G204gat), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n478_), .A2(new_n480_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT21), .ZN(new_n483_));
  INV_X1    g282(.A(G218gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n484_), .A2(G211gat), .ZN(new_n485_));
  INV_X1    g284(.A(G211gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(G218gat), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n483_), .B1(new_n485_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n482_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G197gat), .B(G204gat), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n485_), .B(new_n487_), .C1(new_n490_), .C2(new_n483_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n478_), .A2(new_n480_), .A3(new_n483_), .A4(new_n481_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  OAI21_X1  g292(.A(new_n489_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(G233gat), .ZN(new_n495_));
  NOR2_X1   g294(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(KEYINPUT86), .A2(G228gat), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n495_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n475_), .A2(new_n494_), .A3(new_n500_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n458_), .B1(new_n430_), .B2(new_n434_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n485_), .A2(new_n487_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n479_), .A2(G197gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(new_n481_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n503_), .B1(KEYINPUT21), .B2(new_n505_), .ZN(new_n506_));
  AOI22_X1  g305(.A1(new_n506_), .A2(new_n492_), .B1(new_n482_), .B2(new_n488_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n499_), .B1(new_n502_), .B2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n474_), .A2(new_n501_), .A3(new_n508_), .ZN(new_n509_));
  AND3_X1   g308(.A1(new_n467_), .A2(new_n470_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n501_), .A2(new_n508_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(new_n472_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n512_), .A2(KEYINPUT91), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT91), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n511_), .A2(new_n514_), .A3(new_n472_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n513_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n510_), .A2(new_n516_), .ZN(new_n517_));
  AOI21_X1  g316(.A(new_n500_), .B1(new_n475_), .B2(new_n494_), .ZN(new_n518_));
  NOR3_X1   g317(.A1(new_n502_), .A2(new_n507_), .A3(new_n499_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n473_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n520_), .A2(KEYINPUT90), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT90), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n511_), .A2(new_n522_), .A3(new_n473_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n523_), .A3(new_n509_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n467_), .A2(new_n470_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n517_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT27), .ZN(new_n528_));
  NAND2_X1  g327(.A1(G226gat), .A2(G233gat), .ZN(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT19), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n354_), .A2(new_n352_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n368_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(new_n382_), .A3(new_n378_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT80), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n354_), .A2(new_n536_), .ZN(new_n537_));
  AND3_X1   g336(.A1(new_n376_), .A2(new_n537_), .A3(new_n369_), .ZN(new_n538_));
  NAND4_X1  g337(.A1(new_n344_), .A2(new_n346_), .A3(KEYINPUT24), .A4(new_n337_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n359_), .A2(KEYINPUT26), .ZN(new_n540_));
  INV_X1    g339(.A(G183gat), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n541_), .A2(KEYINPUT25), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT25), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(G183gat), .ZN(new_n544_));
  NAND4_X1  g343(.A1(new_n540_), .A2(new_n364_), .A3(new_n542_), .A4(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(G169gat), .A2(G176gat), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(new_n350_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n539_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n535_), .B1(new_n538_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n531_), .B1(new_n549_), .B2(new_n494_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n374_), .A2(new_n375_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n537_), .A2(new_n369_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n533_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(new_n378_), .A2(new_n382_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n507_), .B1(new_n555_), .B2(new_n367_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT20), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n550_), .A2(new_n556_), .A3(new_n557_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n557_), .B1(new_n549_), .B2(new_n494_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n555_), .A2(new_n367_), .A3(new_n507_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n531_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  XOR2_X1   g360(.A(G8gat), .B(G36gat), .Z(new_n562_));
  XNOR2_X1  g361(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  XNOR2_X1  g363(.A(G64gat), .B(G92gat), .ZN(new_n565_));
  XNOR2_X1  g364(.A(new_n564_), .B(new_n565_), .ZN(new_n566_));
  NOR3_X1   g365(.A1(new_n558_), .A2(new_n561_), .A3(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n566_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n539_), .A2(new_n545_), .A3(new_n547_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n376_), .A2(new_n537_), .A3(new_n369_), .ZN(new_n570_));
  AOI22_X1  g369(.A1(new_n569_), .A2(new_n570_), .B1(new_n554_), .B2(new_n534_), .ZN(new_n571_));
  OAI21_X1  g370(.A(KEYINPUT20), .B1(new_n571_), .B2(new_n507_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n348_), .A2(new_n355_), .A3(new_n366_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n383_), .B1(new_n570_), .B2(new_n533_), .ZN(new_n574_));
  NOR3_X1   g373(.A1(new_n573_), .A2(new_n574_), .A3(new_n494_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n530_), .B1(new_n572_), .B2(new_n575_), .ZN(new_n576_));
  INV_X1    g375(.A(new_n550_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n557_), .B1(new_n384_), .B2(new_n494_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n568_), .B1(new_n576_), .B2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n528_), .B1(new_n567_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT96), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n549_), .A2(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(KEYINPUT96), .B(new_n535_), .C1(new_n538_), .C2(new_n548_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n583_), .A2(new_n507_), .A3(new_n584_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n531_), .B1(new_n585_), .B2(new_n578_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n572_), .A2(new_n575_), .A3(new_n530_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n566_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n576_), .A2(new_n579_), .A3(new_n568_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(KEYINPUT27), .A3(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n581_), .A2(new_n590_), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT98), .B1(new_n527_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n591_), .ZN(new_n593_));
  AOI22_X1  g392(.A1(new_n510_), .A2(new_n516_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT98), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n455_), .B1(new_n592_), .B2(new_n596_), .ZN(new_n597_));
  AOI211_X1 g396(.A(KEYINPUT95), .B(KEYINPUT33), .C1(new_n453_), .C2(new_n444_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT95), .ZN(new_n599_));
  NAND3_X1  g398(.A1(new_n444_), .A2(new_n445_), .A3(new_n451_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT33), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n599_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n598_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n453_), .A2(KEYINPUT33), .A3(new_n444_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n566_), .B1(new_n558_), .B2(new_n561_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n441_), .A2(new_n442_), .ZN(new_n606_));
  NAND3_X1  g405(.A1(new_n438_), .A2(new_n606_), .A3(new_n439_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n440_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n436_), .A2(new_n437_), .A3(new_n608_), .ZN(new_n609_));
  NAND3_X1  g408(.A1(new_n607_), .A2(new_n452_), .A3(new_n609_), .ZN(new_n610_));
  AND4_X1   g409(.A1(new_n604_), .A2(new_n605_), .A3(new_n589_), .A4(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n568_), .A2(KEYINPUT32), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n612_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n568_), .A2(KEYINPUT32), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n576_), .A2(new_n579_), .A3(new_n614_), .ZN(new_n615_));
  AND2_X1   g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n446_), .A2(new_n452_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n600_), .ZN(new_n618_));
  AOI22_X1  g417(.A1(new_n603_), .A2(new_n611_), .B1(new_n616_), .B2(new_n618_), .ZN(new_n619_));
  OAI21_X1  g418(.A(KEYINPUT97), .B1(new_n619_), .B2(new_n527_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n618_), .A2(new_n613_), .A3(new_n615_), .ZN(new_n621_));
  AND2_X1   g420(.A1(new_n438_), .A2(new_n443_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n445_), .A2(new_n451_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n601_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n624_), .A2(KEYINPUT95), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n600_), .A2(new_n599_), .A3(new_n601_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n605_), .A2(new_n604_), .A3(new_n589_), .A4(new_n610_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n621_), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT97), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n630_), .A3(new_n594_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n581_), .A2(new_n590_), .A3(new_n454_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n594_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n620_), .A2(new_n631_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n412_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n597_), .B1(new_n635_), .B2(new_n636_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n318_), .A2(new_n276_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT75), .ZN(new_n639_));
  INV_X1    g438(.A(new_n318_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n276_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n639_), .B(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(G229gat), .A2(G233gat), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n643_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n283_), .A2(new_n640_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n647_), .A2(new_n644_), .A3(new_n638_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n646_), .A2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(G113gat), .B(G141gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(G169gat), .B(G197gat), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n650_), .B(new_n651_), .Z(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n649_), .A2(new_n653_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n646_), .A2(new_n648_), .A3(new_n652_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n637_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n336_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n660_), .A2(new_n309_), .A3(new_n618_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT38), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT99), .Z(new_n663_));
  INV_X1    g462(.A(new_n271_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n664_), .A2(new_n657_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n637_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n298_), .A2(new_n302_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n667_), .ZN(new_n668_));
  NOR2_X1   g467(.A1(new_n668_), .A2(new_n334_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n666_), .A2(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n665_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G1gat), .B1(new_n672_), .B2(new_n454_), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n663_), .B(new_n673_), .C1(KEYINPUT38), .C2(new_n661_), .ZN(G1324gat));
  NOR3_X1   g473(.A1(new_n659_), .A2(G8gat), .A3(new_n593_), .ZN(new_n675_));
  OAI21_X1  g474(.A(G8gat), .B1(new_n672_), .B2(new_n593_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n676_), .A2(KEYINPUT39), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(KEYINPUT39), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n675_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n679_), .B(new_n680_), .Z(G1325gat));
  OAI21_X1  g480(.A(G15gat), .B1(new_n672_), .B2(new_n636_), .ZN(new_n682_));
  XOR2_X1   g481(.A(new_n682_), .B(KEYINPUT41), .Z(new_n683_));
  NAND3_X1  g482(.A1(new_n660_), .A2(new_n405_), .A3(new_n412_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n683_), .A2(new_n684_), .ZN(G1326gat));
  OAI21_X1  g484(.A(G22gat), .B1(new_n672_), .B2(new_n594_), .ZN(new_n686_));
  XOR2_X1   g485(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  OR2_X1    g487(.A1(new_n594_), .A2(G22gat), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n688_), .B1(new_n659_), .B2(new_n689_), .ZN(G1327gat));
  INV_X1    g489(.A(new_n334_), .ZN(new_n691_));
  NOR3_X1   g490(.A1(new_n664_), .A2(new_n691_), .A3(new_n667_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n692_), .A2(new_n658_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  AOI21_X1  g493(.A(G29gat), .B1(new_n694_), .B2(new_n618_), .ZN(new_n695_));
  INV_X1    g494(.A(new_n308_), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n637_), .A2(KEYINPUT43), .A3(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT104), .B1(new_n304_), .B2(new_n307_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT104), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n303_), .A2(new_n306_), .A3(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n702_), .B1(new_n637_), .B2(KEYINPUT103), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n629_), .A2(new_n594_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n633_), .B1(new_n704_), .B2(KEYINPUT97), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n412_), .B1(new_n705_), .B2(new_n631_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n707_));
  NOR3_X1   g506(.A1(new_n706_), .A2(new_n707_), .A3(new_n597_), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT105), .B(KEYINPUT43), .C1(new_n703_), .C2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n707_), .B1(new_n706_), .B2(new_n597_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n635_), .A2(new_n636_), .ZN(new_n712_));
  INV_X1    g511(.A(new_n597_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n712_), .A2(KEYINPUT103), .A3(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n711_), .A2(new_n714_), .A3(new_n702_), .ZN(new_n715_));
  AOI21_X1  g514(.A(KEYINPUT105), .B1(new_n715_), .B2(KEYINPUT43), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n698_), .B1(new_n710_), .B2(new_n716_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n271_), .A2(new_n656_), .A3(new_n334_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT102), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n717_), .A2(KEYINPUT44), .A3(new_n720_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n721_), .A2(KEYINPUT106), .ZN(new_n722_));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n723_));
  NAND4_X1  g522(.A1(new_n717_), .A2(new_n723_), .A3(KEYINPUT44), .A4(new_n720_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n722_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726_));
  OAI21_X1  g525(.A(KEYINPUT43), .B1(new_n703_), .B2(new_n708_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT105), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n697_), .B1(new_n729_), .B2(new_n709_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n718_), .B(KEYINPUT102), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n726_), .B1(new_n730_), .B2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n725_), .A2(new_n732_), .ZN(new_n733_));
  INV_X1    g532(.A(new_n733_), .ZN(new_n734_));
  AND2_X1   g533(.A1(new_n618_), .A2(G29gat), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n695_), .B1(new_n734_), .B2(new_n735_), .ZN(G1328gat));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737_));
  INV_X1    g536(.A(G36gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(KEYINPUT44), .B1(new_n717_), .B2(new_n720_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n739_), .A2(new_n593_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n725_), .B2(new_n740_), .ZN(new_n741_));
  OR2_X1    g540(.A1(new_n591_), .A2(KEYINPUT107), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n591_), .A2(KEYINPUT107), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NOR3_X1   g544(.A1(new_n693_), .A2(G36gat), .A3(new_n745_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT45), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n737_), .B1(new_n741_), .B2(new_n747_), .ZN(new_n748_));
  INV_X1    g547(.A(new_n747_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n732_), .A2(new_n591_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n750_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n749_), .B(KEYINPUT46), .C1(new_n751_), .C2(new_n738_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n748_), .A2(new_n752_), .ZN(G1329gat));
  NAND2_X1  g552(.A1(new_n412_), .A2(G43gat), .ZN(new_n754_));
  AOI211_X1 g553(.A(new_n739_), .B(new_n754_), .C1(new_n722_), .C2(new_n724_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(KEYINPUT108), .B(G43gat), .ZN(new_n756_));
  OAI21_X1  g555(.A(new_n756_), .B1(new_n693_), .B2(new_n636_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(KEYINPUT47), .B1(new_n755_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT47), .ZN(new_n760_));
  OAI211_X1 g559(.A(new_n760_), .B(new_n757_), .C1(new_n733_), .C2(new_n754_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n759_), .A2(new_n761_), .ZN(G1330gat));
  AOI21_X1  g561(.A(G50gat), .B1(new_n694_), .B2(new_n527_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n527_), .A2(G50gat), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n763_), .B1(new_n734_), .B2(new_n764_), .ZN(G1331gat));
  NAND2_X1  g564(.A1(new_n666_), .A2(new_n657_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT109), .ZN(new_n767_));
  AND3_X1   g566(.A1(new_n767_), .A2(new_n335_), .A3(new_n664_), .ZN(new_n768_));
  AOI21_X1  g567(.A(G57gat), .B1(new_n768_), .B2(new_n618_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT110), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n664_), .A2(new_n657_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n771_), .A2(new_n670_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n618_), .A2(G57gat), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n770_), .B1(new_n772_), .B2(new_n773_), .ZN(G1332gat));
  INV_X1    g573(.A(G64gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n775_), .B1(new_n772_), .B2(new_n744_), .ZN(new_n776_));
  XOR2_X1   g575(.A(new_n776_), .B(KEYINPUT48), .Z(new_n777_));
  NAND3_X1  g576(.A1(new_n768_), .A2(new_n775_), .A3(new_n744_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(G1333gat));
  INV_X1    g578(.A(G71gat), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n780_), .B1(new_n772_), .B2(new_n412_), .ZN(new_n781_));
  XOR2_X1   g580(.A(new_n781_), .B(KEYINPUT49), .Z(new_n782_));
  NAND3_X1  g581(.A1(new_n768_), .A2(new_n780_), .A3(new_n412_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(G1334gat));
  INV_X1    g583(.A(G78gat), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n785_), .B1(new_n772_), .B2(new_n527_), .ZN(new_n786_));
  XOR2_X1   g585(.A(new_n786_), .B(KEYINPUT50), .Z(new_n787_));
  NAND3_X1  g586(.A1(new_n768_), .A2(new_n785_), .A3(new_n527_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1335gat));
  NOR3_X1   g588(.A1(new_n271_), .A2(new_n691_), .A3(new_n667_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n767_), .A2(new_n790_), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n791_), .A2(new_n454_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n792_), .A2(G85gat), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT111), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n771_), .A2(new_n691_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n730_), .A2(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n618_), .A2(G85gat), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(G1336gat));
  NOR3_X1   g598(.A1(new_n791_), .A2(G92gat), .A3(new_n593_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n744_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n800_), .B1(new_n801_), .B2(G92gat), .ZN(new_n802_));
  XNOR2_X1  g601(.A(new_n802_), .B(KEYINPUT112), .ZN(G1337gat));
  OR3_X1    g602(.A1(new_n791_), .A2(new_n636_), .A3(new_n225_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n717_), .A2(new_n412_), .A3(new_n795_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(G99gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n805_), .B2(G99gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n804_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(new_n809_), .B(KEYINPUT51), .ZN(G1338gat));
  NOR3_X1   g609(.A1(new_n730_), .A2(new_n796_), .A3(new_n594_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812_));
  INV_X1    g611(.A(G106gat), .ZN(new_n813_));
  OR3_X1    g612(.A1(new_n811_), .A2(new_n812_), .A3(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n812_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n767_), .A2(new_n813_), .A3(new_n527_), .A4(new_n790_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT114), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n814_), .A2(new_n815_), .A3(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT53), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n814_), .A2(new_n820_), .A3(new_n815_), .A4(new_n817_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1339gat));
  NAND4_X1  g621(.A1(new_n267_), .A2(new_n335_), .A3(new_n657_), .A4(new_n270_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT54), .ZN(new_n824_));
  XNOR2_X1  g623(.A(new_n823_), .B(new_n824_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT56), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(KEYINPUT116), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n210_), .B1(new_n256_), .B2(new_n258_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT55), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n260_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n256_), .A2(new_n258_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n831_), .A2(KEYINPUT55), .A3(new_n209_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n208_), .B1(new_n830_), .B2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT115), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n827_), .B1(new_n833_), .B2(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n208_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n259_), .B1(KEYINPUT55), .B2(new_n828_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n832_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n836_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n839_), .A2(KEYINPUT115), .A3(new_n826_), .ZN(new_n840_));
  OAI211_X1 g639(.A(KEYINPUT56), .B(new_n836_), .C1(new_n837_), .C2(new_n838_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(KEYINPUT116), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n835_), .A2(new_n840_), .A3(new_n842_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n657_), .A2(new_n265_), .ZN(new_n844_));
  AND2_X1   g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n643_), .A2(new_n644_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n653_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n847_), .A2(KEYINPUT117), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT117), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n846_), .A2(new_n849_), .A3(new_n653_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n647_), .A2(new_n645_), .A3(new_n638_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n848_), .A2(new_n850_), .A3(new_n851_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n852_), .A2(new_n655_), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n853_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT57), .B(new_n667_), .C1(new_n845_), .C2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n854_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n856_), .B1(new_n857_), .B2(new_n668_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n839_), .A2(new_n826_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n859_), .A2(new_n860_), .A3(new_n841_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n839_), .A2(KEYINPUT118), .A3(new_n826_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n853_), .A2(new_n265_), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n861_), .A2(new_n862_), .A3(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT58), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n861_), .A2(new_n863_), .A3(KEYINPUT58), .A4(new_n862_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n866_), .A2(new_n308_), .A3(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n855_), .A2(new_n858_), .A3(new_n868_), .ZN(new_n869_));
  AOI21_X1  g668(.A(new_n825_), .B1(new_n869_), .B2(new_n334_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n592_), .A2(new_n596_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n871_), .A2(new_n412_), .A3(new_n618_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n870_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(G113gat), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n873_), .A2(new_n874_), .A3(new_n656_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n870_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n872_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(KEYINPUT59), .A3(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n879_), .B1(new_n870_), .B2(new_n872_), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n657_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n875_), .B1(new_n881_), .B2(new_n874_), .ZN(G1340gat));
  INV_X1    g681(.A(G120gat), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n883_), .B1(new_n271_), .B2(KEYINPUT60), .ZN(new_n884_));
  OAI211_X1 g683(.A(new_n873_), .B(new_n884_), .C1(KEYINPUT60), .C2(new_n883_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n271_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n886_));
  OAI21_X1  g685(.A(new_n885_), .B1(new_n886_), .B2(new_n883_), .ZN(new_n887_));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI211_X1 g688(.A(KEYINPUT119), .B(new_n885_), .C1(new_n886_), .C2(new_n883_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1341gat));
  AOI21_X1  g690(.A(G127gat), .B1(new_n873_), .B2(new_n691_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n878_), .A2(new_n880_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n334_), .A2(KEYINPUT120), .ZN(new_n894_));
  MUX2_X1   g693(.A(KEYINPUT120), .B(new_n894_), .S(G127gat), .Z(new_n895_));
  AOI21_X1  g694(.A(new_n892_), .B1(new_n893_), .B2(new_n895_), .ZN(G1342gat));
  NAND3_X1  g695(.A1(new_n873_), .A2(new_n390_), .A3(new_n668_), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n696_), .B1(new_n878_), .B2(new_n880_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n897_), .B1(new_n898_), .B2(new_n390_), .ZN(G1343gat));
  NOR4_X1   g698(.A1(new_n744_), .A2(new_n412_), .A3(new_n594_), .A4(new_n454_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n876_), .A2(new_n900_), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n901_), .A2(new_n657_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(KEYINPUT121), .B(G141gat), .ZN(new_n903_));
  XNOR2_X1  g702(.A(new_n902_), .B(new_n903_), .ZN(G1344gat));
  INV_X1    g703(.A(new_n901_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n664_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G148gat), .ZN(G1345gat));
  OR3_X1    g706(.A1(new_n901_), .A2(KEYINPUT122), .A3(new_n334_), .ZN(new_n908_));
  OAI21_X1  g707(.A(KEYINPUT122), .B1(new_n901_), .B2(new_n334_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT61), .B(G155gat), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n908_), .A2(new_n909_), .A3(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n910_), .B1(new_n908_), .B2(new_n909_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n911_), .A2(new_n912_), .ZN(G1346gat));
  AOI21_X1  g712(.A(G162gat), .B1(new_n905_), .B2(new_n668_), .ZN(new_n914_));
  NOR3_X1   g713(.A1(new_n699_), .A2(new_n701_), .A3(new_n414_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n905_), .B2(new_n915_), .ZN(G1347gat));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917_));
  NOR2_X1   g716(.A1(new_n745_), .A2(new_n455_), .ZN(new_n918_));
  XOR2_X1   g717(.A(new_n918_), .B(KEYINPUT123), .Z(new_n919_));
  NOR2_X1   g718(.A1(new_n919_), .A2(new_n527_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n876_), .A2(new_n920_), .ZN(new_n921_));
  OAI21_X1  g720(.A(KEYINPUT124), .B1(new_n921_), .B2(new_n657_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(G169gat), .ZN(new_n923_));
  NOR3_X1   g722(.A1(new_n921_), .A2(KEYINPUT124), .A3(new_n657_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n917_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n921_), .ZN(new_n926_));
  NAND4_X1  g725(.A1(new_n926_), .A2(new_n656_), .A3(new_n379_), .A4(new_n381_), .ZN(new_n927_));
  OR3_X1    g726(.A1(new_n921_), .A2(KEYINPUT124), .A3(new_n657_), .ZN(new_n928_));
  NAND4_X1  g727(.A1(new_n928_), .A2(KEYINPUT62), .A3(new_n922_), .A4(G169gat), .ZN(new_n929_));
  NAND3_X1  g728(.A1(new_n925_), .A2(new_n927_), .A3(new_n929_), .ZN(G1348gat));
  NAND2_X1  g729(.A1(new_n926_), .A2(new_n664_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n931_), .B1(new_n932_), .B2(new_n343_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(KEYINPUT125), .B(G176gat), .ZN(new_n934_));
  AOI21_X1  g733(.A(new_n933_), .B1(new_n931_), .B2(new_n934_), .ZN(G1349gat));
  NAND2_X1  g734(.A1(new_n926_), .A2(new_n691_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n936_), .A2(new_n363_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n937_), .B1(new_n541_), .B2(new_n936_), .ZN(G1350gat));
  NAND4_X1  g737(.A1(new_n926_), .A2(new_n540_), .A3(new_n364_), .A4(new_n668_), .ZN(new_n939_));
  OAI21_X1  g738(.A(G190gat), .B1(new_n921_), .B2(new_n696_), .ZN(new_n940_));
  NAND2_X1  g739(.A1(new_n939_), .A2(new_n940_), .ZN(G1351gat));
  NAND3_X1  g740(.A1(new_n636_), .A2(new_n527_), .A3(new_n454_), .ZN(new_n942_));
  NOR3_X1   g741(.A1(new_n870_), .A2(new_n745_), .A3(new_n942_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n943_), .A2(new_n656_), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n944_), .B(G197gat), .ZN(G1352gat));
  AOI22_X1  g744(.A1(new_n943_), .A2(new_n664_), .B1(KEYINPUT126), .B2(new_n479_), .ZN(new_n946_));
  NOR2_X1   g745(.A1(new_n479_), .A2(KEYINPUT126), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(KEYINPUT127), .ZN(new_n948_));
  XNOR2_X1  g747(.A(new_n946_), .B(new_n948_), .ZN(G1353gat));
  NAND2_X1  g748(.A1(new_n943_), .A2(new_n691_), .ZN(new_n950_));
  NOR2_X1   g749(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n951_));
  AND2_X1   g750(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n950_), .A2(new_n951_), .A3(new_n952_), .ZN(new_n953_));
  AOI21_X1  g752(.A(new_n953_), .B1(new_n950_), .B2(new_n951_), .ZN(G1354gat));
  NAND3_X1  g753(.A1(new_n943_), .A2(new_n484_), .A3(new_n668_), .ZN(new_n955_));
  AND2_X1   g754(.A1(new_n943_), .A2(new_n308_), .ZN(new_n956_));
  OAI21_X1  g755(.A(new_n955_), .B1(new_n956_), .B2(new_n484_), .ZN(G1355gat));
endmodule


