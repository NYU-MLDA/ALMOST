//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n886_, new_n888_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n921_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n929_, new_n930_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n205_), .A3(KEYINPUT88), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT88), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n207_), .B1(new_n202_), .B2(new_n204_), .ZN(new_n208_));
  AND3_X1   g007(.A1(new_n202_), .A2(new_n204_), .A3(KEYINPUT87), .ZN(new_n209_));
  AOI21_X1  g008(.A(KEYINPUT87), .B1(new_n202_), .B2(new_n204_), .ZN(new_n210_));
  OAI211_X1 g009(.A(new_n206_), .B(new_n208_), .C1(new_n209_), .C2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  AOI21_X1  g013(.A(new_n213_), .B1(KEYINPUT1), .B2(new_n214_), .ZN(new_n215_));
  OR2_X1    g014(.A1(new_n214_), .A2(KEYINPUT1), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G141gat), .A2(G148gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  NOR2_X1   g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n217_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT3), .ZN(new_n223_));
  INV_X1    g022(.A(G141gat), .ZN(new_n224_));
  INV_X1    g023(.A(G148gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n223_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT2), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n218_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n229_));
  OAI21_X1  g028(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n230_));
  NAND4_X1  g029(.A1(new_n226_), .A2(new_n228_), .A3(new_n229_), .A4(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT90), .ZN(new_n232_));
  XOR2_X1   g031(.A(G155gat), .B(G162gat), .Z(new_n233_));
  AND3_X1   g032(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n232_), .B1(new_n231_), .B2(new_n233_), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n222_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n212_), .A2(new_n236_), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n202_), .B(new_n204_), .ZN(new_n238_));
  OAI211_X1 g037(.A(new_n222_), .B(new_n238_), .C1(new_n234_), .C2(new_n235_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G225gat), .A2(G233gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(KEYINPUT100), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n237_), .A2(new_n239_), .A3(new_n241_), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G1gat), .B(G29gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(G85gat), .ZN(new_n244_));
  XNOR2_X1  g043(.A(KEYINPUT0), .B(G57gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n244_), .B(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  AOI21_X1  g046(.A(KEYINPUT4), .B1(new_n212_), .B2(new_n236_), .ZN(new_n248_));
  AOI211_X1 g047(.A(new_n219_), .B(new_n220_), .C1(new_n215_), .C2(new_n216_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n231_), .A2(new_n233_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(KEYINPUT90), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n231_), .A2(new_n232_), .A3(new_n233_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n249_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n239_), .B1(new_n253_), .B2(new_n211_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n248_), .B1(KEYINPUT4), .B2(new_n254_), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n241_), .B(KEYINPUT101), .ZN(new_n256_));
  OAI211_X1 g055(.A(new_n242_), .B(new_n247_), .C1(new_n255_), .C2(new_n256_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n246_), .B1(new_n254_), .B2(new_n256_), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n254_), .A2(KEYINPUT4), .ZN(new_n259_));
  INV_X1    g058(.A(new_n248_), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n258_), .B1(new_n261_), .B2(new_n241_), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT33), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n257_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  XOR2_X1   g063(.A(G8gat), .B(G36gat), .Z(new_n265_));
  XNOR2_X1  g064(.A(new_n265_), .B(KEYINPUT18), .ZN(new_n266_));
  XNOR2_X1  g065(.A(G64gat), .B(G92gat), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT19), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT20), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT97), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(G197gat), .A2(G204gat), .ZN(new_n277_));
  INV_X1    g076(.A(G204gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(KEYINPUT93), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT93), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(G204gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n279_), .A2(new_n281_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n277_), .B1(new_n282_), .B2(G197gat), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n276_), .A2(KEYINPUT21), .A3(new_n283_), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n274_), .B(KEYINPUT97), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT96), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT95), .B(KEYINPUT21), .ZN(new_n287_));
  INV_X1    g086(.A(G197gat), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n288_), .B1(new_n279_), .B2(new_n281_), .ZN(new_n289_));
  OAI211_X1 g088(.A(new_n286_), .B(new_n287_), .C1(new_n289_), .C2(new_n277_), .ZN(new_n290_));
  INV_X1    g089(.A(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n277_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT93), .B(G204gat), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n292_), .B1(new_n293_), .B2(new_n288_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n286_), .B1(new_n294_), .B2(new_n287_), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n285_), .B1(new_n291_), .B2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n278_), .A2(G197gat), .ZN(new_n297_));
  AOI21_X1  g096(.A(G197gat), .B1(new_n279_), .B2(new_n281_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT94), .ZN(new_n299_));
  OAI21_X1  g098(.A(new_n297_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  NOR3_X1   g099(.A1(new_n293_), .A2(KEYINPUT94), .A3(G197gat), .ZN(new_n301_));
  OAI21_X1  g100(.A(KEYINPUT21), .B1(new_n300_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n284_), .B1(new_n296_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305_));
  OAI21_X1  g104(.A(KEYINPUT85), .B1(G169gat), .B2(G176gat), .ZN(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NOR3_X1   g106(.A1(KEYINPUT85), .A2(G169gat), .A3(G176gat), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n305_), .B1(new_n307_), .B2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT25), .B(G183gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT26), .B(G190gat), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(G183gat), .A2(G190gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(KEYINPUT23), .ZN(new_n314_));
  AND3_X1   g113(.A1(new_n309_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n305_), .B1(G169gat), .B2(G176gat), .ZN(new_n316_));
  INV_X1    g115(.A(KEYINPUT85), .ZN(new_n317_));
  INV_X1    g116(.A(G169gat), .ZN(new_n318_));
  INV_X1    g117(.A(G176gat), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(KEYINPUT86), .A3(new_n306_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  AOI21_X1  g121(.A(KEYINPUT86), .B1(new_n320_), .B2(new_n306_), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n316_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT23), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n313_), .A2(new_n325_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n327_));
  OAI211_X1 g126(.A(new_n326_), .B(new_n327_), .C1(G183gat), .C2(G190gat), .ZN(new_n328_));
  NAND2_X1  g127(.A1(G169gat), .A2(G176gat), .ZN(new_n329_));
  AND2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n318_), .A2(KEYINPUT22), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT22), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(G169gat), .ZN(new_n333_));
  INV_X1    g132(.A(KEYINPUT99), .ZN(new_n334_));
  AND3_X1   g133(.A1(new_n331_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n334_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n319_), .B1(new_n335_), .B2(new_n336_), .ZN(new_n337_));
  AOI22_X1  g136(.A1(new_n315_), .A2(new_n324_), .B1(new_n330_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  AOI21_X1  g138(.A(new_n273_), .B1(new_n304_), .B2(new_n339_), .ZN(new_n340_));
  AND3_X1   g139(.A1(new_n276_), .A2(KEYINPUT21), .A3(new_n283_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n287_), .ZN(new_n342_));
  OAI21_X1  g141(.A(KEYINPUT96), .B1(new_n283_), .B2(new_n342_), .ZN(new_n343_));
  AOI21_X1  g142(.A(new_n276_), .B1(new_n343_), .B2(new_n290_), .ZN(new_n344_));
  AOI21_X1  g143(.A(new_n341_), .B1(new_n344_), .B2(new_n302_), .ZN(new_n345_));
  OAI21_X1  g144(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n332_), .A2(new_n318_), .A3(new_n319_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n328_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT84), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n312_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n310_), .A2(new_n311_), .A3(KEYINPUT84), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n323_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n353_), .A2(new_n305_), .A3(new_n321_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n352_), .A2(new_n324_), .A3(new_n354_), .A4(new_n314_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n345_), .A2(new_n348_), .A3(new_n355_), .ZN(new_n356_));
  AOI21_X1  g155(.A(new_n272_), .B1(new_n340_), .B2(new_n356_), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n284_), .B(new_n338_), .C1(new_n296_), .C2(new_n303_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT20), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n302_), .B(new_n285_), .C1(new_n295_), .C2(new_n291_), .ZN(new_n360_));
  AOI22_X1  g159(.A1(new_n360_), .A2(new_n284_), .B1(new_n355_), .B2(new_n348_), .ZN(new_n361_));
  NOR3_X1   g160(.A1(new_n359_), .A2(new_n271_), .A3(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n269_), .B1(new_n357_), .B2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT20), .B1(new_n345_), .B2(new_n338_), .ZN(new_n364_));
  AND4_X1   g163(.A1(new_n360_), .A2(new_n284_), .A3(new_n348_), .A4(new_n355_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n271_), .B1(new_n364_), .B2(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n273_), .B1(new_n345_), .B2(new_n338_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n355_), .A2(new_n348_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n304_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n367_), .A2(new_n272_), .A3(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n366_), .A2(new_n268_), .A3(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(new_n256_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n261_), .A2(new_n372_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n373_), .A2(KEYINPUT33), .A3(new_n242_), .A4(new_n247_), .ZN(new_n374_));
  NAND4_X1  g173(.A1(new_n264_), .A2(new_n363_), .A3(new_n371_), .A4(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT102), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n268_), .A2(KEYINPUT32), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NOR3_X1   g177(.A1(new_n364_), .A2(new_n365_), .A3(new_n271_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n272_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n376_), .B(new_n378_), .C1(new_n379_), .C2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n256_), .B1(new_n259_), .B2(new_n260_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n242_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n246_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n384_), .A2(new_n257_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n366_), .A2(new_n377_), .A3(new_n370_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n381_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n340_), .A2(new_n272_), .A3(new_n356_), .ZN(new_n388_));
  OAI21_X1  g187(.A(new_n271_), .B1(new_n359_), .B2(new_n361_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n376_), .B1(new_n390_), .B2(new_n378_), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n375_), .B1(new_n387_), .B2(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n393_));
  XOR2_X1   g192(.A(G22gat), .B(G50gat), .Z(new_n394_));
  OAI21_X1  g193(.A(new_n394_), .B1(new_n236_), .B2(KEYINPUT29), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT29), .ZN(new_n396_));
  INV_X1    g195(.A(new_n394_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n253_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n393_), .B1(new_n395_), .B2(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT98), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n395_), .A2(new_n398_), .A3(new_n393_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n400_), .A2(new_n401_), .A3(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n402_), .ZN(new_n404_));
  OAI21_X1  g203(.A(KEYINPUT98), .B1(new_n404_), .B2(new_n399_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n403_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n253_), .A2(new_n396_), .ZN(new_n408_));
  OAI21_X1  g207(.A(G78gat), .B1(new_n345_), .B2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(G78gat), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n236_), .A2(KEYINPUT29), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n304_), .A2(new_n410_), .A3(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(G106gat), .ZN(new_n413_));
  AND3_X1   g212(.A1(new_n409_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n413_), .B1(new_n409_), .B2(new_n412_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G228gat), .A2(G233gat), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n416_), .B1(new_n345_), .B2(KEYINPUT92), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR3_X1   g217(.A1(new_n414_), .A2(new_n415_), .A3(new_n418_), .ZN(new_n419_));
  NOR3_X1   g218(.A1(new_n345_), .A2(new_n408_), .A3(G78gat), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n410_), .B1(new_n304_), .B2(new_n411_), .ZN(new_n421_));
  OAI21_X1  g220(.A(G106gat), .B1(new_n420_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n409_), .A2(new_n412_), .A3(new_n413_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n417_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n407_), .B1(new_n419_), .B2(new_n424_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n418_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n417_), .A3(new_n423_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n403_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n426_), .A2(new_n427_), .A3(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n425_), .A2(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n392_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(KEYINPUT103), .ZN(new_n432_));
  AND3_X1   g231(.A1(new_n426_), .A2(new_n428_), .A3(new_n427_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n406_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n434_));
  NOR2_X1   g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n371_), .A2(KEYINPUT27), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n268_), .B(KEYINPUT105), .Z(new_n437_));
  AOI21_X1  g236(.A(new_n437_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n436_), .A2(new_n438_), .ZN(new_n439_));
  AOI21_X1  g238(.A(KEYINPUT27), .B1(new_n363_), .B2(new_n371_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n385_), .B(KEYINPUT104), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n435_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT103), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n392_), .A2(new_n444_), .A3(new_n430_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n432_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G227gat), .A2(G233gat), .ZN(new_n447_));
  XOR2_X1   g246(.A(new_n447_), .B(G15gat), .Z(new_n448_));
  XNOR2_X1  g247(.A(new_n448_), .B(KEYINPUT30), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n368_), .B(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(new_n211_), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452_));
  INV_X1    g251(.A(G43gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT31), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n451_), .B(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT89), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n456_), .B(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n441_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(new_n435_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n442_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n461_), .A2(new_n456_), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n446_), .A2(new_n458_), .B1(new_n460_), .B2(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G29gat), .B(G36gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G43gat), .B(G50gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT75), .B(KEYINPUT15), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XOR2_X1   g267(.A(G15gat), .B(G22gat), .Z(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT78), .B(G1gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(G8gat), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n469_), .B1(new_n471_), .B2(KEYINPUT14), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n472_), .B(KEYINPUT79), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G1gat), .B(G8gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT79), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n472_), .B(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n474_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n468_), .B1(new_n475_), .B2(new_n479_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n480_), .A2(KEYINPUT83), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(KEYINPUT83), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n475_), .A2(new_n479_), .A3(new_n466_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G229gat), .A2(G233gat), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n483_), .A2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G113gat), .B(G141gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(G169gat), .B(G197gat), .ZN(new_n490_));
  XOR2_X1   g289(.A(new_n489_), .B(new_n490_), .Z(new_n491_));
  AOI21_X1  g290(.A(new_n466_), .B1(new_n475_), .B2(new_n479_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  AND2_X1   g292(.A1(new_n493_), .A2(new_n484_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n488_), .B(new_n491_), .C1(new_n494_), .C2(new_n485_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n491_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n494_), .A2(new_n485_), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n486_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n498_));
  OAI21_X1  g297(.A(new_n496_), .B1(new_n497_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n463_), .A2(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT12), .ZN(new_n503_));
  XOR2_X1   g302(.A(G85gat), .B(G92gat), .Z(new_n504_));
  INV_X1    g303(.A(KEYINPUT8), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT67), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT6), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n508_), .B1(G99gat), .B2(G106gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G99gat), .A2(G106gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n510_), .A2(KEYINPUT6), .ZN(new_n511_));
  OAI21_X1  g310(.A(new_n507_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  OR3_X1    g311(.A1(KEYINPUT68), .A2(G99gat), .A3(G106gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(KEYINPUT7), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n510_), .A2(KEYINPUT6), .ZN(new_n515_));
  NAND3_X1  g314(.A1(new_n508_), .A2(G99gat), .A3(G106gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n515_), .A2(new_n516_), .A3(KEYINPUT67), .ZN(new_n517_));
  NOR3_X1   g316(.A1(KEYINPUT68), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT7), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n512_), .A2(new_n514_), .A3(new_n517_), .A4(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT69), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n506_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  AND2_X1   g322(.A1(new_n514_), .A2(new_n520_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n524_), .A2(KEYINPUT69), .A3(new_n517_), .A4(new_n512_), .ZN(new_n525_));
  OAI21_X1  g324(.A(KEYINPUT70), .B1(new_n509_), .B2(new_n511_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT70), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n515_), .A2(new_n516_), .A3(new_n527_), .ZN(new_n528_));
  NAND4_X1  g327(.A1(new_n526_), .A2(new_n528_), .A3(new_n514_), .A4(new_n520_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(new_n504_), .ZN(new_n530_));
  AOI22_X1  g329(.A1(new_n523_), .A2(new_n525_), .B1(new_n530_), .B2(KEYINPUT8), .ZN(new_n531_));
  INV_X1    g330(.A(G85gat), .ZN(new_n532_));
  INV_X1    g331(.A(G92gat), .ZN(new_n533_));
  NOR3_X1   g332(.A1(new_n532_), .A2(new_n533_), .A3(KEYINPUT9), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n504_), .B2(KEYINPUT9), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT10), .B(G99gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(KEYINPUT66), .B(G106gat), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n512_), .A2(new_n517_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n531_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G57gat), .B(G64gat), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n544_));
  XOR2_X1   g343(.A(G71gat), .B(G78gat), .Z(new_n545_));
  OR2_X1    g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n545_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n543_), .A2(KEYINPUT11), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n546_), .B1(new_n547_), .B2(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n503_), .B1(new_n542_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n542_), .A2(new_n549_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G230gat), .A2(G233gat), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n552_), .B(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n523_), .A2(new_n525_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n530_), .A2(KEYINPUT8), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT71), .B1(new_n539_), .B2(new_n540_), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n512_), .A2(new_n517_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT71), .ZN(new_n560_));
  NAND4_X1  g359(.A1(new_n559_), .A2(new_n560_), .A3(new_n538_), .A4(new_n535_), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n558_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n557_), .A2(new_n562_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n549_), .A2(new_n503_), .ZN(new_n564_));
  INV_X1    g363(.A(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n563_), .A2(new_n565_), .ZN(new_n566_));
  NAND4_X1  g365(.A1(new_n550_), .A2(new_n551_), .A3(new_n554_), .A4(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n554_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n542_), .A2(new_n549_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n541_), .ZN(new_n570_));
  AND3_X1   g369(.A1(new_n557_), .A2(new_n549_), .A3(new_n570_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n568_), .B1(new_n569_), .B2(new_n571_), .ZN(new_n572_));
  XOR2_X1   g371(.A(G120gat), .B(G148gat), .Z(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n574_));
  XNOR2_X1  g373(.A(new_n573_), .B(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G176gat), .B(G204gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n567_), .A2(new_n572_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT73), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n567_), .A2(new_n572_), .A3(KEYINPUT73), .A4(new_n578_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  AOI21_X1  g382(.A(new_n578_), .B1(new_n567_), .B2(new_n572_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n586_), .A2(KEYINPUT74), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT74), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n583_), .A2(new_n588_), .A3(new_n585_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n587_), .A2(KEYINPUT13), .A3(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT13), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n588_), .B1(new_n583_), .B2(new_n585_), .ZN(new_n592_));
  AOI211_X1 g391(.A(KEYINPUT74), .B(new_n584_), .C1(new_n581_), .C2(new_n582_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n591_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n590_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n549_), .B(new_n596_), .Z(new_n597_));
  NAND2_X1  g396(.A1(new_n475_), .A2(new_n479_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n597_), .B(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(G127gat), .B(G155gat), .Z(new_n600_));
  XNOR2_X1  g399(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(G183gat), .B(G211gat), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n599_), .A2(KEYINPUT17), .A3(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(KEYINPUT81), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n604_), .B(KEYINPUT17), .ZN(new_n607_));
  XNOR2_X1  g406(.A(new_n607_), .B(KEYINPUT82), .ZN(new_n608_));
  OR2_X1    g407(.A1(new_n608_), .A2(new_n599_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n606_), .A2(new_n609_), .ZN(new_n610_));
  INV_X1    g409(.A(new_n610_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n557_), .A2(new_n466_), .A3(new_n570_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n468_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n558_), .A2(new_n561_), .ZN(new_n614_));
  OAI21_X1  g413(.A(new_n613_), .B1(new_n531_), .B2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n612_), .A2(new_n615_), .A3(KEYINPUT76), .ZN(new_n616_));
  XNOR2_X1  g415(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n617_));
  NAND2_X1  g416(.A1(G232gat), .A2(G233gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n616_), .A2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n612_), .A2(new_n615_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT35), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n612_), .A2(new_n615_), .A3(KEYINPUT76), .A4(new_n619_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n621_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  XNOR2_X1  g425(.A(G190gat), .B(G218gat), .ZN(new_n627_));
  XNOR2_X1  g426(.A(G134gat), .B(G162gat), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n627_), .B(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n629_), .A2(KEYINPUT36), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n626_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n629_), .A2(KEYINPUT36), .ZN(new_n632_));
  AND3_X1   g431(.A1(new_n626_), .A2(KEYINPUT77), .A3(new_n632_), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n632_), .B1(new_n626_), .B2(KEYINPUT77), .ZN(new_n634_));
  OAI21_X1  g433(.A(new_n631_), .B1(new_n633_), .B2(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT37), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT37), .ZN(new_n637_));
  OAI211_X1 g436(.A(new_n631_), .B(new_n637_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n611_), .A2(new_n636_), .A3(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n595_), .A2(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n502_), .A2(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n641_), .B(KEYINPUT106), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n442_), .B(KEYINPUT107), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n643_), .A2(new_n470_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n642_), .A2(new_n644_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n645_), .A2(KEYINPUT38), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n645_), .A2(KEYINPUT38), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n463_), .A2(new_n635_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n595_), .A2(new_n501_), .A3(new_n610_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  OAI21_X1  g450(.A(G1gat), .B1(new_n651_), .B2(new_n442_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n646_), .A2(new_n647_), .A3(new_n652_), .ZN(G1324gat));
  INV_X1    g452(.A(G8gat), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n642_), .A2(new_n654_), .A3(new_n459_), .ZN(new_n655_));
  OAI21_X1  g454(.A(G8gat), .B1(new_n651_), .B2(new_n441_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n656_), .A2(KEYINPUT39), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(KEYINPUT39), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n655_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT40), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(KEYINPUT40), .B(new_n655_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n661_), .A2(new_n662_), .ZN(G1325gat));
  OAI21_X1  g462(.A(G15gat), .B1(new_n651_), .B2(new_n458_), .ZN(new_n664_));
  OR2_X1    g463(.A1(new_n664_), .A2(KEYINPUT41), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n664_), .A2(KEYINPUT41), .ZN(new_n666_));
  NOR3_X1   g465(.A1(new_n641_), .A2(G15gat), .A3(new_n458_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT108), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n665_), .A2(new_n666_), .A3(new_n668_), .ZN(G1326gat));
  INV_X1    g468(.A(G22gat), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n670_), .B1(new_n650_), .B2(new_n435_), .ZN(new_n671_));
  XOR2_X1   g470(.A(new_n671_), .B(KEYINPUT42), .Z(new_n672_));
  NAND2_X1  g471(.A1(new_n435_), .A2(new_n670_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n672_), .B1(new_n641_), .B2(new_n673_), .ZN(G1327gat));
  NAND2_X1  g473(.A1(new_n610_), .A2(new_n635_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n595_), .A2(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n502_), .A2(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G29gat), .B1(new_n677_), .B2(new_n461_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n636_), .A2(new_n638_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n680_), .ZN(new_n681_));
  NOR3_X1   g480(.A1(new_n463_), .A2(KEYINPUT43), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n636_), .A2(KEYINPUT109), .A3(new_n638_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  OAI21_X1  g485(.A(KEYINPUT43), .B1(new_n463_), .B2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(KEYINPUT110), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n443_), .A2(new_n445_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n444_), .B1(new_n392_), .B2(new_n430_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n458_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n460_), .A2(new_n462_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AND3_X1   g492(.A1(new_n636_), .A2(KEYINPUT109), .A3(new_n638_), .ZN(new_n694_));
  AOI21_X1  g493(.A(KEYINPUT109), .B1(new_n636_), .B2(new_n638_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n693_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT110), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n697_), .A2(new_n698_), .A3(KEYINPUT43), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n682_), .B1(new_n688_), .B2(new_n699_), .ZN(new_n700_));
  AND2_X1   g499(.A1(new_n590_), .A2(new_n594_), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n701_), .A2(new_n500_), .A3(new_n610_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n679_), .B1(new_n700_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n682_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n698_), .B1(new_n697_), .B2(KEYINPUT43), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT43), .ZN(new_n706_));
  AOI211_X1 g505(.A(KEYINPUT110), .B(new_n706_), .C1(new_n693_), .C2(new_n696_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n704_), .B1(new_n705_), .B2(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(new_n702_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n708_), .A2(KEYINPUT44), .A3(new_n709_), .ZN(new_n710_));
  AND2_X1   g509(.A1(new_n703_), .A2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n643_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n712_), .A2(G29gat), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n678_), .B1(new_n711_), .B2(new_n713_), .ZN(G1328gat));
  XNOR2_X1  g513(.A(KEYINPUT111), .B(KEYINPUT46), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n703_), .A2(new_n710_), .A3(new_n459_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G36gat), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n441_), .A2(G36gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n502_), .A2(new_n676_), .A3(new_n718_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT45), .Z(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(new_n715_), .B1(new_n717_), .B2(new_n721_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n715_), .ZN(new_n723_));
  AOI211_X1 g522(.A(new_n720_), .B(new_n723_), .C1(new_n716_), .C2(G36gat), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n722_), .A2(new_n724_), .ZN(G1329gat));
  INV_X1    g524(.A(new_n456_), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n703_), .A2(new_n710_), .A3(G43gat), .A4(new_n726_), .ZN(new_n727_));
  INV_X1    g526(.A(new_n458_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n677_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(new_n453_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n727_), .A2(new_n730_), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g531(.A(G50gat), .B1(new_n677_), .B2(new_n435_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n435_), .A2(G50gat), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n711_), .B2(new_n734_), .ZN(G1331gat));
  NOR2_X1   g534(.A1(new_n463_), .A2(new_n500_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n701_), .A2(new_n639_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  OR2_X1    g538(.A1(new_n739_), .A2(KEYINPUT112), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(KEYINPUT112), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n740_), .A2(new_n712_), .A3(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(G57gat), .ZN(new_n743_));
  AND4_X1   g542(.A1(new_n501_), .A2(new_n648_), .A3(new_n595_), .A4(new_n611_), .ZN(new_n744_));
  NOR2_X1   g543(.A1(new_n442_), .A2(new_n743_), .ZN(new_n745_));
  AOI22_X1  g544(.A1(new_n742_), .A2(new_n743_), .B1(new_n744_), .B2(new_n745_), .ZN(G1332gat));
  INV_X1    g545(.A(G64gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n747_), .B1(new_n744_), .B2(new_n459_), .ZN(new_n748_));
  XOR2_X1   g547(.A(new_n748_), .B(KEYINPUT48), .Z(new_n749_));
  NAND3_X1  g548(.A1(new_n739_), .A2(new_n747_), .A3(new_n459_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(G1333gat));
  INV_X1    g550(.A(G71gat), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n744_), .B2(new_n728_), .ZN(new_n753_));
  XOR2_X1   g552(.A(new_n753_), .B(KEYINPUT49), .Z(new_n754_));
  NAND3_X1  g553(.A1(new_n739_), .A2(new_n752_), .A3(new_n728_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n754_), .A2(new_n755_), .ZN(G1334gat));
  AOI21_X1  g555(.A(new_n410_), .B1(new_n744_), .B2(new_n435_), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT50), .Z(new_n758_));
  NOR2_X1   g557(.A1(new_n430_), .A2(G78gat), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT113), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n758_), .B1(new_n738_), .B2(new_n760_), .ZN(G1335gat));
  NOR2_X1   g560(.A1(new_n701_), .A2(new_n675_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n736_), .A2(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n764_), .A2(new_n532_), .A3(new_n712_), .ZN(new_n765_));
  NAND3_X1  g564(.A1(new_n595_), .A2(new_n501_), .A3(new_n610_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT114), .ZN(new_n767_));
  INV_X1    g566(.A(new_n767_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n700_), .A2(new_n442_), .A3(new_n768_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n765_), .B1(new_n769_), .B2(new_n532_), .ZN(G1336gat));
  NAND3_X1  g569(.A1(new_n764_), .A2(new_n533_), .A3(new_n459_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n700_), .A2(new_n441_), .A3(new_n768_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(new_n533_), .ZN(G1337gat));
  NOR3_X1   g572(.A1(new_n763_), .A2(new_n456_), .A3(new_n536_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n700_), .A2(new_n768_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n775_), .A2(new_n728_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n774_), .B1(new_n776_), .B2(G99gat), .ZN(new_n777_));
  NAND2_X1  g576(.A1(KEYINPUT115), .A2(KEYINPUT51), .ZN(new_n778_));
  XNOR2_X1  g577(.A(new_n777_), .B(new_n778_), .ZN(G1338gat));
  OR3_X1    g578(.A1(new_n763_), .A2(new_n430_), .A3(new_n537_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n708_), .A2(new_n435_), .A3(new_n767_), .ZN(new_n781_));
  INV_X1    g580(.A(KEYINPUT52), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n781_), .A2(new_n782_), .A3(G106gat), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n782_), .B1(new_n781_), .B2(G106gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n780_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(KEYINPUT53), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT53), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n787_), .B(new_n780_), .C1(new_n783_), .C2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n786_), .A2(new_n788_), .ZN(G1339gat));
  NAND3_X1  g588(.A1(new_n712_), .A2(new_n726_), .A3(new_n460_), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT118), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n792_), .A2(KEYINPUT57), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n485_), .ZN(new_n795_));
  OAI211_X1 g594(.A(KEYINPUT117), .B(new_n496_), .C1(new_n494_), .C2(new_n795_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n483_), .A2(new_n484_), .A3(new_n795_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT117), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n795_), .B1(new_n493_), .B2(new_n484_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n491_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n796_), .A2(new_n797_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n495_), .ZN(new_n802_));
  INV_X1    g601(.A(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n803_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n804_));
  AOI22_X1  g603(.A1(new_n563_), .A2(new_n565_), .B1(new_n542_), .B2(new_n549_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(new_n550_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n568_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n567_), .A2(new_n808_), .ZN(new_n809_));
  NAND4_X1  g608(.A1(new_n805_), .A2(KEYINPUT55), .A3(new_n554_), .A4(new_n550_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n807_), .A2(new_n809_), .A3(new_n810_), .ZN(new_n811_));
  AND3_X1   g610(.A1(new_n811_), .A2(KEYINPUT56), .A3(new_n577_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT56), .B1(new_n811_), .B2(new_n577_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n500_), .B(new_n583_), .C1(new_n812_), .C2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n804_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n635_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n794_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  AOI211_X1 g616(.A(new_n635_), .B(new_n793_), .C1(new_n804_), .C2(new_n814_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n811_), .A2(KEYINPUT56), .A3(new_n577_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT119), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n811_), .A2(KEYINPUT119), .A3(KEYINPUT56), .A4(new_n577_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n811_), .A2(new_n577_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT56), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n822_), .A2(new_n823_), .A3(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n802_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT58), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n827_), .A2(new_n828_), .A3(KEYINPUT58), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n831_), .A2(new_n680_), .A3(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n611_), .B1(new_n819_), .B2(new_n833_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n639_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n701_), .A2(new_n501_), .A3(new_n835_), .ZN(new_n836_));
  XOR2_X1   g635(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n838_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n640_), .A2(new_n501_), .A3(new_n837_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n791_), .B1(new_n834_), .B2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(KEYINPUT120), .A2(KEYINPUT59), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  INV_X1    g645(.A(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n842_), .A2(new_n847_), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n791_), .B(new_n843_), .C1(new_n834_), .C2(new_n841_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n848_), .A2(new_n849_), .ZN(new_n850_));
  OAI21_X1  g649(.A(G113gat), .B1(new_n850_), .B2(new_n501_), .ZN(new_n851_));
  OR2_X1    g650(.A1(new_n501_), .A2(G113gat), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n851_), .B1(new_n842_), .B2(new_n852_), .ZN(G1340gat));
  NAND2_X1  g652(.A1(new_n815_), .A2(new_n816_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n793_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n815_), .A2(new_n816_), .A3(new_n794_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n855_), .A2(new_n833_), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n610_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n837_), .B1(new_n640_), .B2(new_n501_), .ZN(new_n859_));
  NOR4_X1   g658(.A1(new_n595_), .A2(new_n639_), .A3(new_n500_), .A4(new_n838_), .ZN(new_n860_));
  NOR2_X1   g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n790_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n849_), .B(new_n595_), .C1(new_n862_), .C2(new_n846_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT121), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n701_), .A2(G120gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n862_), .B1(KEYINPUT60), .B2(new_n865_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n848_), .A2(new_n867_), .A3(new_n595_), .A4(new_n849_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n864_), .A2(new_n866_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(G120gat), .ZN(new_n870_));
  OR2_X1    g669(.A1(new_n866_), .A2(KEYINPUT60), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(G1341gat));
  INV_X1    g671(.A(G127gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n873_), .B1(new_n842_), .B2(new_n610_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n874_), .A2(KEYINPUT122), .ZN(new_n875_));
  XOR2_X1   g674(.A(KEYINPUT123), .B(G127gat), .Z(new_n876_));
  NAND4_X1  g675(.A1(new_n848_), .A2(new_n611_), .A3(new_n849_), .A4(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n874_), .A2(KEYINPUT122), .ZN(new_n878_));
  AND3_X1   g677(.A1(new_n875_), .A2(new_n877_), .A3(new_n878_), .ZN(G1342gat));
  OAI21_X1  g678(.A(G134gat), .B1(new_n850_), .B2(new_n681_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n816_), .A2(G134gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n842_), .B2(new_n881_), .ZN(G1343gat));
  NAND2_X1  g681(.A1(new_n858_), .A2(new_n861_), .ZN(new_n883_));
  NOR4_X1   g682(.A1(new_n728_), .A2(new_n643_), .A3(new_n430_), .A4(new_n459_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n885_), .A2(new_n501_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(new_n224_), .ZN(G1344gat));
  NOR2_X1   g686(.A1(new_n885_), .A2(new_n701_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(new_n888_), .B(new_n225_), .ZN(G1345gat));
  NOR2_X1   g688(.A1(new_n885_), .A2(new_n610_), .ZN(new_n890_));
  XOR2_X1   g689(.A(KEYINPUT61), .B(G155gat), .Z(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1346gat));
  INV_X1    g691(.A(G162gat), .ZN(new_n893_));
  NOR3_X1   g692(.A1(new_n885_), .A2(new_n893_), .A3(new_n686_), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n883_), .A2(new_n635_), .A3(new_n884_), .ZN(new_n895_));
  AND2_X1   g694(.A1(new_n895_), .A2(new_n893_), .ZN(new_n896_));
  OR2_X1    g695(.A1(new_n896_), .A2(KEYINPUT124), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(KEYINPUT124), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n894_), .B1(new_n897_), .B2(new_n898_), .ZN(G1347gat));
  NOR3_X1   g698(.A1(new_n712_), .A2(new_n435_), .A3(new_n458_), .ZN(new_n900_));
  OAI211_X1 g699(.A(new_n459_), .B(new_n900_), .C1(new_n834_), .C2(new_n841_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT125), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n901_), .A2(new_n902_), .ZN(new_n903_));
  NAND4_X1  g702(.A1(new_n883_), .A2(KEYINPUT125), .A3(new_n459_), .A4(new_n900_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n905_), .B(new_n500_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n906_));
  INV_X1    g705(.A(new_n901_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(new_n500_), .ZN(new_n908_));
  INV_X1    g707(.A(KEYINPUT62), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n908_), .A2(new_n909_), .A3(G169gat), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n909_), .B1(new_n908_), .B2(G169gat), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n906_), .B1(new_n911_), .B2(new_n912_), .ZN(G1348gat));
  NAND3_X1  g712(.A1(new_n905_), .A2(new_n319_), .A3(new_n595_), .ZN(new_n914_));
  OAI21_X1  g713(.A(G176gat), .B1(new_n901_), .B2(new_n701_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(G1349gat));
  AOI21_X1  g715(.A(G183gat), .B1(new_n907_), .B2(new_n611_), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n610_), .A2(new_n310_), .ZN(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n917_), .B1(new_n905_), .B2(new_n919_), .ZN(G1350gat));
  NAND3_X1  g719(.A1(new_n905_), .A2(new_n311_), .A3(new_n635_), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n441_), .B1(new_n858_), .B2(new_n861_), .ZN(new_n922_));
  AOI21_X1  g721(.A(KEYINPUT125), .B1(new_n922_), .B2(new_n900_), .ZN(new_n923_));
  NOR2_X1   g722(.A1(new_n901_), .A2(new_n902_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n680_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(KEYINPUT126), .B1(new_n925_), .B2(G190gat), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n681_), .B1(new_n903_), .B2(new_n904_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT126), .ZN(new_n928_));
  INV_X1    g727(.A(G190gat), .ZN(new_n929_));
  NOR3_X1   g728(.A1(new_n927_), .A2(new_n928_), .A3(new_n929_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n921_), .B1(new_n926_), .B2(new_n930_), .ZN(G1351gat));
  NAND2_X1  g730(.A1(new_n883_), .A2(new_n459_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n458_), .A2(new_n435_), .A3(new_n442_), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n933_), .B(KEYINPUT127), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n932_), .A2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n500_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n595_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n293_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n939_), .B1(new_n278_), .B2(new_n938_), .ZN(G1353gat));
  AOI211_X1 g739(.A(KEYINPUT63), .B(G211gat), .C1(new_n935_), .C2(new_n611_), .ZN(new_n941_));
  INV_X1    g740(.A(new_n935_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n610_), .ZN(new_n943_));
  XOR2_X1   g742(.A(KEYINPUT63), .B(G211gat), .Z(new_n944_));
  AOI21_X1  g743(.A(new_n941_), .B1(new_n943_), .B2(new_n944_), .ZN(G1354gat));
  OAI21_X1  g744(.A(G218gat), .B1(new_n942_), .B2(new_n681_), .ZN(new_n946_));
  OR2_X1    g745(.A1(new_n816_), .A2(G218gat), .ZN(new_n947_));
  OAI21_X1  g746(.A(new_n946_), .B1(new_n942_), .B2(new_n947_), .ZN(G1355gat));
endmodule


