//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n695_,
    new_n696_, new_n697_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n822_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n900_, new_n901_, new_n902_, new_n903_, new_n905_,
    new_n906_, new_n907_, new_n908_, new_n909_, new_n910_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n953_, new_n954_, new_n955_,
    new_n957_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n968_, new_n969_, new_n970_;
  INV_X1    g000(.A(KEYINPUT29), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT3), .ZN(new_n203_));
  INV_X1    g002(.A(G141gat), .ZN(new_n204_));
  INV_X1    g003(.A(G148gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT2), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND3_X1  g008(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n206_), .A2(new_n209_), .A3(new_n210_), .A4(new_n211_), .ZN(new_n212_));
  OR2_X1    g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214_));
  AND2_X1   g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n212_), .A2(new_n215_), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT82), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT82), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(G141gat), .B2(G148gat), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n213_), .A2(new_n221_), .A3(new_n214_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n223_), .A2(new_n207_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n220_), .A2(new_n222_), .A3(new_n224_), .ZN(new_n225_));
  AND3_X1   g024(.A1(new_n216_), .A2(KEYINPUT83), .A3(new_n225_), .ZN(new_n226_));
  AOI21_X1  g025(.A(KEYINPUT83), .B1(new_n216_), .B2(new_n225_), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n202_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(KEYINPUT28), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT28), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n230_), .B(new_n202_), .C1(new_n226_), .C2(new_n227_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n229_), .A2(new_n231_), .ZN(new_n232_));
  XNOR2_X1  g031(.A(G22gat), .B(G50gat), .ZN(new_n233_));
  XOR2_X1   g032(.A(new_n233_), .B(KEYINPUT84), .Z(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n229_), .A2(new_n231_), .A3(new_n234_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT85), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n236_), .A2(KEYINPUT85), .A3(new_n237_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n216_), .A2(new_n225_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT83), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n242_), .A2(new_n243_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n216_), .A2(new_n225_), .A3(KEYINPUT83), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n244_), .A2(KEYINPUT29), .A3(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT90), .ZN(new_n247_));
  INV_X1    g046(.A(G211gat), .ZN(new_n248_));
  NOR2_X1   g047(.A1(new_n248_), .A2(G218gat), .ZN(new_n249_));
  INV_X1    g048(.A(G218gat), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n250_), .A2(G211gat), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n247_), .B1(new_n249_), .B2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(G197gat), .ZN(new_n253_));
  OAI21_X1  g052(.A(KEYINPUT87), .B1(new_n253_), .B2(G204gat), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT87), .ZN(new_n255_));
  INV_X1    g054(.A(G204gat), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(G197gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n253_), .A2(G204gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n254_), .A2(new_n257_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n250_), .A2(G211gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n248_), .A2(G218gat), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(KEYINPUT90), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n252_), .A2(new_n259_), .A3(KEYINPUT21), .A4(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n260_), .A2(new_n261_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n256_), .A2(G197gat), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n265_), .A2(new_n258_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n264_), .B1(KEYINPUT21), .B2(new_n266_), .ZN(new_n267_));
  AND2_X1   g066(.A1(KEYINPUT88), .A2(KEYINPUT21), .ZN(new_n268_));
  NOR2_X1   g067(.A1(KEYINPUT88), .A2(KEYINPUT21), .ZN(new_n269_));
  NOR2_X1   g068(.A1(new_n268_), .A2(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n270_), .A2(new_n254_), .A3(new_n258_), .A4(new_n257_), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n267_), .A2(KEYINPUT89), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT89), .B1(new_n267_), .B2(new_n271_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n263_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G228gat), .A2(G233gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(new_n275_), .B(KEYINPUT86), .Z(new_n276_));
  AND3_X1   g075(.A1(new_n246_), .A2(new_n274_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n277_), .ZN(new_n278_));
  XNOR2_X1  g077(.A(G78gat), .B(G106gat), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n279_), .B(KEYINPUT92), .Z(new_n280_));
  INV_X1    g079(.A(KEYINPUT91), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n242_), .A2(KEYINPUT29), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n274_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n276_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n281_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(new_n263_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT89), .ZN(new_n287_));
  XNOR2_X1  g086(.A(KEYINPUT88), .B(KEYINPUT21), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n259_), .A2(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(G197gat), .B(G204gat), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT21), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n260_), .B(new_n261_), .C1(new_n290_), .C2(new_n291_), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n287_), .B1(new_n289_), .B2(new_n292_), .ZN(new_n293_));
  NAND3_X1  g092(.A1(new_n267_), .A2(KEYINPUT89), .A3(new_n271_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n286_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n282_), .ZN(new_n296_));
  OAI211_X1 g095(.A(new_n281_), .B(new_n284_), .C1(new_n295_), .C2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(new_n278_), .B(new_n280_), .C1(new_n285_), .C2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n284_), .B1(new_n295_), .B2(new_n296_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n301_), .A2(KEYINPUT91), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(new_n297_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n280_), .B1(new_n303_), .B2(new_n278_), .ZN(new_n304_));
  OAI211_X1 g103(.A(new_n240_), .B(new_n241_), .C1(new_n300_), .C2(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n277_), .B1(new_n302_), .B2(new_n297_), .ZN(new_n306_));
  AOI22_X1  g105(.A1(new_n306_), .A2(new_n280_), .B1(new_n237_), .B2(new_n236_), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n278_), .B1(new_n285_), .B2(new_n298_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT93), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n308_), .A2(new_n309_), .A3(new_n279_), .ZN(new_n310_));
  INV_X1    g109(.A(new_n279_), .ZN(new_n311_));
  OAI21_X1  g110(.A(KEYINPUT93), .B1(new_n306_), .B2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n307_), .A2(new_n310_), .A3(new_n312_), .ZN(new_n313_));
  AND2_X1   g112(.A1(new_n305_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(G8gat), .B(G36gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT18), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G64gat), .B(G92gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(G169gat), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT96), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G183gat), .A2(G190gat), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(KEYINPUT79), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT79), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(G183gat), .A3(G190gat), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT23), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(KEYINPUT23), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G183gat), .A2(G190gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n322_), .B1(new_n330_), .B2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n331_), .ZN(new_n333_));
  OAI211_X1 g132(.A(KEYINPUT96), .B(new_n333_), .C1(new_n327_), .C2(new_n329_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n321_), .B1(new_n332_), .B2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n325_), .B1(G183gat), .B2(G190gat), .ZN(new_n336_));
  NOR2_X1   g135(.A1(new_n323_), .A2(KEYINPUT79), .ZN(new_n337_));
  OAI21_X1  g136(.A(KEYINPUT23), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT23), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n323_), .A2(new_n339_), .ZN(new_n340_));
  AND2_X1   g139(.A1(new_n338_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(G169gat), .ZN(new_n342_));
  INV_X1    g141(.A(G176gat), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n345_));
  NOR2_X1   g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  NOR3_X1   g145(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n347_));
  NOR2_X1   g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  XNOR2_X1  g147(.A(KEYINPUT26), .B(G190gat), .ZN(new_n349_));
  INV_X1    g148(.A(G183gat), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n350_), .A2(KEYINPUT25), .ZN(new_n351_));
  OR2_X1    g150(.A1(new_n350_), .A2(KEYINPUT25), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n349_), .A2(new_n351_), .A3(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n341_), .A2(new_n348_), .A3(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n354_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n274_), .B1(new_n335_), .B2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT20), .ZN(new_n357_));
  INV_X1    g156(.A(new_n347_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n358_), .B1(new_n344_), .B2(new_n345_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n349_), .A2(new_n352_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n351_), .A2(new_n361_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n350_), .A2(KEYINPUT78), .A3(KEYINPUT25), .ZN(new_n363_));
  AND2_X1   g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n359_), .B1(new_n360_), .B2(new_n364_), .ZN(new_n365_));
  OAI21_X1  g164(.A(new_n339_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(new_n328_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n338_), .A2(new_n333_), .A3(new_n340_), .ZN(new_n368_));
  AOI22_X1  g167(.A1(new_n365_), .A2(new_n367_), .B1(new_n368_), .B2(new_n320_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n357_), .B1(new_n295_), .B2(new_n369_), .ZN(new_n370_));
  XOR2_X1   g169(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n371_));
  NAND2_X1  g170(.A1(G226gat), .A2(G233gat), .ZN(new_n372_));
  XNOR2_X1  g171(.A(new_n371_), .B(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT95), .ZN(new_n374_));
  AND3_X1   g173(.A1(new_n356_), .A2(new_n370_), .A3(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n368_), .A2(new_n320_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n349_), .A2(new_n352_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n362_), .A2(new_n363_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n348_), .B1(new_n377_), .B2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n376_), .B1(new_n379_), .B2(new_n330_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n357_), .B1(new_n274_), .B2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(KEYINPUT96), .B1(new_n367_), .B2(new_n333_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n334_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n320_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n384_), .A2(new_n295_), .A3(new_n354_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n373_), .B1(new_n381_), .B2(new_n385_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n318_), .B1(new_n375_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n374_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n295_), .B1(new_n384_), .B2(new_n354_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT20), .B1(new_n274_), .B2(new_n380_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n388_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n381_), .A2(new_n385_), .A3(new_n373_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n318_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n391_), .A2(new_n392_), .A3(new_n393_), .ZN(new_n394_));
  AND3_X1   g193(.A1(new_n387_), .A2(KEYINPUT27), .A3(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT97), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n394_), .A2(new_n396_), .ZN(new_n397_));
  NAND4_X1  g196(.A1(new_n391_), .A2(KEYINPUT97), .A3(new_n392_), .A4(new_n393_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n391_), .A2(new_n392_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n318_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n397_), .A2(new_n398_), .A3(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT27), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n395_), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(G127gat), .B(G134gat), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G113gat), .B(G120gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n407_), .A2(KEYINPUT31), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT81), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT31), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n409_), .B1(new_n406_), .B2(new_n410_), .ZN(new_n411_));
  XOR2_X1   g210(.A(G15gat), .B(G43gat), .Z(new_n412_));
  OR3_X1    g211(.A1(new_n408_), .A2(new_n411_), .A3(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n412_), .B1(new_n408_), .B2(new_n411_), .ZN(new_n414_));
  AND2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(G227gat), .A2(G233gat), .ZN(new_n416_));
  XOR2_X1   g215(.A(new_n416_), .B(KEYINPUT80), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT30), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n380_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n369_), .A2(new_n418_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  XNOR2_X1  g221(.A(G71gat), .B(G99gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n423_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n420_), .A2(new_n421_), .A3(new_n425_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n415_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n427_));
  AOI21_X1  g226(.A(new_n415_), .B1(new_n424_), .B2(new_n426_), .ZN(new_n428_));
  NOR2_X1   g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G1gat), .B(G29gat), .ZN(new_n430_));
  XNOR2_X1  g229(.A(new_n430_), .B(G85gat), .ZN(new_n431_));
  XNOR2_X1  g230(.A(KEYINPUT0), .B(G57gat), .ZN(new_n432_));
  XOR2_X1   g231(.A(new_n431_), .B(new_n432_), .Z(new_n433_));
  INV_X1    g232(.A(KEYINPUT98), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n244_), .A2(new_n407_), .A3(new_n434_), .A4(new_n245_), .ZN(new_n435_));
  NOR3_X1   g234(.A1(new_n226_), .A2(new_n227_), .A3(new_n406_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT98), .B1(new_n407_), .B2(new_n242_), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT4), .ZN(new_n439_));
  NAND2_X1  g238(.A1(G225gat), .A2(G233gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n244_), .A2(new_n407_), .A3(new_n245_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n441_), .B1(new_n442_), .B2(KEYINPUT4), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n438_), .A2(new_n440_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n433_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n433_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n443_), .B1(new_n438_), .B2(KEYINPUT4), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n447_), .A2(new_n450_), .ZN(new_n451_));
  AND2_X1   g250(.A1(new_n429_), .A2(new_n451_), .ZN(new_n452_));
  AND3_X1   g251(.A1(new_n314_), .A2(new_n403_), .A3(new_n452_), .ZN(new_n453_));
  OAI211_X1 g252(.A(KEYINPUT32), .B(new_n393_), .C1(new_n375_), .C2(new_n386_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n393_), .A2(KEYINPUT32), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n391_), .A2(new_n392_), .A3(new_n455_), .ZN(new_n456_));
  OAI211_X1 g255(.A(new_n454_), .B(new_n456_), .C1(new_n447_), .C2(new_n450_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT4), .ZN(new_n458_));
  INV_X1    g257(.A(new_n242_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n434_), .B1(new_n459_), .B2(new_n406_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n442_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n458_), .B1(new_n461_), .B2(new_n435_), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n440_), .B1(new_n442_), .B2(KEYINPUT4), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT99), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT99), .ZN(new_n465_));
  INV_X1    g264(.A(new_n463_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n439_), .A2(new_n465_), .A3(new_n466_), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n433_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n464_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NOR3_X1   g268(.A1(new_n448_), .A2(KEYINPUT33), .A3(new_n449_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT33), .ZN(new_n471_));
  INV_X1    g270(.A(new_n433_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n472_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n471_), .B1(new_n445_), .B2(new_n473_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n469_), .B1(new_n470_), .B2(new_n474_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n457_), .B1(new_n475_), .B2(new_n401_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n476_), .A2(new_n314_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n305_), .A2(new_n313_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n401_), .A2(new_n402_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n395_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n478_), .A2(new_n479_), .A3(new_n451_), .A4(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n477_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n429_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n453_), .B1(new_n482_), .B2(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G229gat), .A2(G233gat), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G43gat), .B(G50gat), .ZN(new_n486_));
  INV_X1    g285(.A(new_n486_), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G29gat), .B(G36gat), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n488_), .A2(KEYINPUT71), .ZN(new_n489_));
  INV_X1    g288(.A(G36gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(G29gat), .ZN(new_n491_));
  INV_X1    g290(.A(G29gat), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(G36gat), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n491_), .A2(new_n493_), .A3(KEYINPUT71), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n487_), .B1(new_n489_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n491_), .A2(new_n493_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT71), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n488_), .A2(KEYINPUT71), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(new_n486_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n495_), .A2(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G15gat), .B(G22gat), .ZN(new_n502_));
  INV_X1    g301(.A(G1gat), .ZN(new_n503_));
  INV_X1    g302(.A(G8gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT14), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G1gat), .B(G8gat), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  OR2_X1    g307(.A1(new_n501_), .A2(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n501_), .A2(new_n508_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT76), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n509_), .A2(KEYINPUT76), .A3(new_n510_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n485_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n515_));
  AND3_X1   g314(.A1(new_n495_), .A2(KEYINPUT15), .A3(new_n500_), .ZN(new_n516_));
  AOI21_X1  g315(.A(KEYINPUT15), .B1(new_n495_), .B2(new_n500_), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n508_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n509_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n485_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n515_), .A2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G113gat), .B(G141gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G169gat), .B(G197gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n524_), .B(new_n525_), .Z(new_n526_));
  INV_X1    g325(.A(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(KEYINPUT77), .ZN(new_n529_));
  OR3_X1    g328(.A1(new_n515_), .A2(new_n522_), .A3(new_n527_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n528_), .A2(new_n529_), .A3(new_n530_), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n523_), .A2(KEYINPUT77), .A3(new_n527_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n484_), .A2(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G85gat), .A2(G92gat), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  NOR2_X1   g335(.A1(G85gat), .A2(G92gat), .ZN(new_n537_));
  NOR2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n538_), .A2(KEYINPUT9), .ZN(new_n539_));
  NAND2_X1  g338(.A1(G99gat), .A2(G106gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT6), .ZN(new_n541_));
  OR2_X1    g340(.A1(new_n535_), .A2(KEYINPUT9), .ZN(new_n542_));
  AND2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  XOR2_X1   g342(.A(KEYINPUT10), .B(G99gat), .Z(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NOR3_X1   g344(.A1(new_n545_), .A2(KEYINPUT65), .A3(G106gat), .ZN(new_n546_));
  INV_X1    g345(.A(KEYINPUT65), .ZN(new_n547_));
  INV_X1    g346(.A(G106gat), .ZN(new_n548_));
  AOI21_X1  g347(.A(new_n547_), .B1(new_n544_), .B2(new_n548_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n539_), .B(new_n543_), .C1(new_n546_), .C2(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT6), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n551_), .A2(KEYINPUT66), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT66), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(KEYINPUT6), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n552_), .A2(new_n554_), .A3(new_n540_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n540_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT7), .ZN(new_n557_));
  INV_X1    g356(.A(G99gat), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(new_n548_), .ZN(new_n559_));
  OAI21_X1  g358(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(new_n560_), .ZN(new_n561_));
  NOR3_X1   g360(.A1(new_n555_), .A2(new_n556_), .A3(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n538_), .ZN(new_n563_));
  OAI21_X1  g362(.A(KEYINPUT8), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  AND2_X1   g363(.A1(new_n559_), .A2(new_n560_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(new_n541_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT8), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n566_), .A2(new_n567_), .A3(new_n538_), .ZN(new_n568_));
  AOI21_X1  g367(.A(KEYINPUT68), .B1(new_n564_), .B2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n540_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n553_), .A2(KEYINPUT6), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n551_), .A2(KEYINPUT66), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n552_), .A2(new_n554_), .A3(new_n540_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n565_), .A2(new_n573_), .A3(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n567_), .B1(new_n575_), .B2(new_n538_), .ZN(new_n576_));
  INV_X1    g375(.A(KEYINPUT68), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n538_), .A2(new_n567_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n578_), .B1(new_n541_), .B2(new_n565_), .ZN(new_n579_));
  NOR3_X1   g378(.A1(new_n576_), .A2(new_n577_), .A3(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n550_), .B1(new_n569_), .B2(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G57gat), .B(G64gat), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n582_), .A2(KEYINPUT11), .ZN(new_n583_));
  XOR2_X1   g382(.A(G71gat), .B(G78gat), .Z(new_n584_));
  OR2_X1    g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n582_), .A2(KEYINPUT11), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n583_), .A2(new_n584_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n589_), .A2(KEYINPUT12), .ZN(new_n590_));
  INV_X1    g389(.A(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n556_), .A2(new_n561_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n563_), .B1(new_n592_), .B2(new_n574_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n568_), .B1(new_n593_), .B2(new_n567_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n594_), .A2(new_n550_), .A3(new_n588_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT12), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n594_), .A2(new_n550_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(new_n589_), .ZN(new_n598_));
  AOI22_X1  g397(.A1(new_n581_), .A2(new_n591_), .B1(new_n596_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G230gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n600_), .B(KEYINPUT64), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n599_), .A2(new_n601_), .ZN(new_n602_));
  OR2_X1    g401(.A1(new_n595_), .A2(KEYINPUT67), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n595_), .A2(KEYINPUT67), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n603_), .A2(new_n598_), .A3(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n601_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  XOR2_X1   g407(.A(G120gat), .B(G148gat), .Z(new_n609_));
  XNOR2_X1  g408(.A(G176gat), .B(G204gat), .ZN(new_n610_));
  XNOR2_X1  g409(.A(new_n609_), .B(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT69), .B(KEYINPUT5), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n608_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n613_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n602_), .A2(new_n607_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n614_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT70), .ZN(new_n618_));
  OAI21_X1  g417(.A(new_n617_), .B1(new_n618_), .B2(KEYINPUT13), .ZN(new_n619_));
  XOR2_X1   g418(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n620_));
  NAND3_X1  g419(.A1(new_n614_), .A2(new_n616_), .A3(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n622_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G190gat), .B(G218gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(G134gat), .B(G162gat), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT36), .ZN(new_n627_));
  INV_X1    g426(.A(new_n518_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n581_), .A2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT73), .ZN(new_n630_));
  NAND2_X1  g429(.A1(G232gat), .A2(G233gat), .ZN(new_n631_));
  XOR2_X1   g430(.A(new_n631_), .B(KEYINPUT34), .Z(new_n632_));
  INV_X1    g431(.A(KEYINPUT35), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT72), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n594_), .A2(new_n550_), .ZN(new_n637_));
  AND2_X1   g436(.A1(new_n495_), .A2(new_n500_), .ZN(new_n638_));
  AOI21_X1  g437(.A(new_n636_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n632_), .A2(new_n633_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n629_), .A2(new_n630_), .A3(new_n639_), .A4(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n630_), .ZN(new_n642_));
  OAI21_X1  g441(.A(KEYINPUT73), .B1(new_n632_), .B2(new_n633_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n577_), .B1(new_n576_), .B2(new_n579_), .ZN(new_n644_));
  OAI211_X1 g443(.A(KEYINPUT68), .B(new_n568_), .C1(new_n593_), .C2(new_n567_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n518_), .B1(new_n646_), .B2(new_n550_), .ZN(new_n647_));
  OAI21_X1  g446(.A(new_n635_), .B1(new_n597_), .B2(new_n501_), .ZN(new_n648_));
  OAI211_X1 g447(.A(new_n642_), .B(new_n643_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n626_), .A2(KEYINPUT36), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n641_), .A2(new_n649_), .A3(new_n651_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n641_), .B2(new_n649_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n627_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT74), .ZN(new_n655_));
  OAI21_X1  g454(.A(KEYINPUT37), .B1(new_n653_), .B2(new_n655_), .ZN(new_n656_));
  AND2_X1   g455(.A1(new_n654_), .A2(new_n656_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n654_), .A2(new_n656_), .ZN(new_n658_));
  NOR2_X1   g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(G231gat), .A2(G233gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n508_), .B(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(new_n589_), .ZN(new_n662_));
  XOR2_X1   g461(.A(G127gat), .B(G155gat), .Z(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT16), .ZN(new_n664_));
  XNOR2_X1  g463(.A(G183gat), .B(G211gat), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n664_), .B(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT17), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n662_), .A2(new_n668_), .ZN(new_n669_));
  XNOR2_X1  g468(.A(new_n669_), .B(KEYINPUT75), .ZN(new_n670_));
  AND2_X1   g469(.A1(new_n666_), .A2(new_n667_), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n662_), .A2(new_n668_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n670_), .A2(new_n672_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n623_), .A2(new_n659_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n534_), .A2(new_n674_), .ZN(new_n675_));
  XOR2_X1   g474(.A(new_n675_), .B(KEYINPUT100), .Z(new_n676_));
  INV_X1    g475(.A(new_n451_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n676_), .A2(new_n503_), .A3(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT38), .ZN(new_n679_));
  OR2_X1    g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n484_), .A2(new_n654_), .ZN(new_n681_));
  INV_X1    g480(.A(new_n533_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n673_), .ZN(new_n683_));
  NAND4_X1  g482(.A1(new_n681_), .A2(new_n682_), .A3(new_n683_), .A4(new_n622_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G1gat), .B1(new_n684_), .B2(new_n451_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n678_), .A2(new_n679_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n680_), .A2(new_n685_), .A3(new_n686_), .ZN(G1324gat));
  OAI21_X1  g486(.A(G8gat), .B1(new_n684_), .B2(new_n403_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT39), .ZN(new_n689_));
  INV_X1    g488(.A(new_n403_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n676_), .A2(new_n504_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(G1325gat));
  OAI21_X1  g493(.A(G15gat), .B1(new_n684_), .B2(new_n483_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT41), .ZN(new_n696_));
  NOR3_X1   g495(.A1(new_n675_), .A2(G15gat), .A3(new_n483_), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1326gat));
  OAI21_X1  g497(.A(G22gat), .B1(new_n684_), .B2(new_n314_), .ZN(new_n699_));
  XOR2_X1   g498(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n700_));
  XNOR2_X1  g499(.A(new_n699_), .B(new_n700_), .ZN(new_n701_));
  NOR2_X1   g500(.A1(new_n314_), .A2(G22gat), .ZN(new_n702_));
  XOR2_X1   g501(.A(new_n702_), .B(KEYINPUT103), .Z(new_n703_));
  OAI21_X1  g502(.A(new_n701_), .B1(new_n675_), .B2(new_n703_), .ZN(G1327gat));
  NAND2_X1  g503(.A1(new_n673_), .A2(new_n654_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n623_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n534_), .A2(new_n706_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n707_), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n708_), .A2(new_n492_), .A3(new_n677_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT104), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n710_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n653_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n641_), .A2(new_n649_), .A3(new_n651_), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n712_), .A2(new_n713_), .B1(KEYINPUT36), .B2(new_n626_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n656_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n714_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n654_), .A2(new_n656_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n716_), .A2(KEYINPUT104), .A3(new_n717_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n711_), .A2(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(KEYINPUT43), .B1(new_n484_), .B2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT43), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n659_), .A2(new_n721_), .ZN(new_n722_));
  OAI21_X1  g521(.A(KEYINPUT105), .B1(new_n484_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n716_), .A2(new_n717_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n724_), .A2(KEYINPUT43), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n429_), .B1(new_n477_), .B2(new_n481_), .ZN(new_n727_));
  OAI211_X1 g526(.A(new_n725_), .B(new_n726_), .C1(new_n727_), .C2(new_n453_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n720_), .A2(new_n723_), .A3(new_n728_), .ZN(new_n729_));
  NOR3_X1   g528(.A1(new_n623_), .A2(new_n533_), .A3(new_n683_), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n729_), .A2(KEYINPUT44), .A3(new_n730_), .ZN(new_n731_));
  AOI21_X1  g530(.A(KEYINPUT44), .B1(new_n729_), .B2(new_n730_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n731_), .A2(new_n732_), .A3(new_n451_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n709_), .B1(new_n733_), .B2(new_n492_), .ZN(G1328gat));
  NOR3_X1   g533(.A1(new_n707_), .A2(G36gat), .A3(new_n403_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT45), .Z(new_n736_));
  NOR2_X1   g535(.A1(new_n731_), .A2(new_n732_), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT106), .B1(new_n737_), .B2(new_n690_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n729_), .A2(new_n730_), .ZN(new_n739_));
  INV_X1    g538(.A(KEYINPUT44), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n739_), .A2(new_n740_), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n729_), .A2(new_n730_), .A3(KEYINPUT44), .ZN(new_n742_));
  NAND4_X1  g541(.A1(new_n741_), .A2(KEYINPUT106), .A3(new_n690_), .A4(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n743_), .A2(G36gat), .ZN(new_n744_));
  OAI21_X1  g543(.A(new_n736_), .B1(new_n738_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT107), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT46), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(KEYINPUT107), .A2(KEYINPUT46), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n745_), .A2(new_n748_), .A3(new_n749_), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n741_), .A2(new_n690_), .A3(new_n742_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n753_), .A2(G36gat), .A3(new_n743_), .ZN(new_n754_));
  NAND4_X1  g553(.A1(new_n754_), .A2(new_n746_), .A3(new_n747_), .A4(new_n736_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n750_), .A2(new_n755_), .ZN(G1329gat));
  NAND3_X1  g555(.A1(new_n737_), .A2(G43gat), .A3(new_n429_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n707_), .A2(new_n483_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n757_), .B1(G43gat), .B2(new_n758_), .ZN(new_n759_));
  XNOR2_X1  g558(.A(new_n759_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g559(.A(G50gat), .B1(new_n708_), .B2(new_n478_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n478_), .A2(G50gat), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n761_), .B1(new_n737_), .B2(new_n762_), .ZN(G1331gat));
  NOR2_X1   g562(.A1(new_n484_), .A2(new_n682_), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n764_), .A2(new_n724_), .A3(new_n683_), .A4(new_n623_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT108), .Z(new_n766_));
  INV_X1    g565(.A(G57gat), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n766_), .A2(new_n767_), .A3(new_n677_), .ZN(new_n768_));
  NAND4_X1  g567(.A1(new_n681_), .A2(new_n533_), .A3(new_n683_), .A4(new_n623_), .ZN(new_n769_));
  OAI21_X1  g568(.A(G57gat), .B1(new_n769_), .B2(new_n451_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(G1332gat));
  OAI21_X1  g570(.A(G64gat), .B1(new_n769_), .B2(new_n403_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT109), .ZN(new_n773_));
  INV_X1    g572(.A(new_n773_), .ZN(new_n774_));
  OR2_X1    g573(.A1(new_n774_), .A2(KEYINPUT48), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n774_), .A2(KEYINPUT48), .ZN(new_n776_));
  INV_X1    g575(.A(G64gat), .ZN(new_n777_));
  NAND3_X1  g576(.A1(new_n766_), .A2(new_n777_), .A3(new_n690_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n775_), .A2(new_n776_), .A3(new_n778_), .ZN(G1333gat));
  NOR2_X1   g578(.A1(new_n483_), .A2(G71gat), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT110), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n766_), .A2(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(G71gat), .B1(new_n769_), .B2(new_n483_), .ZN(new_n783_));
  XNOR2_X1  g582(.A(new_n783_), .B(KEYINPUT49), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n782_), .A2(new_n784_), .ZN(G1334gat));
  INV_X1    g584(.A(G78gat), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n766_), .A2(new_n786_), .A3(new_n478_), .ZN(new_n787_));
  OAI21_X1  g586(.A(G78gat), .B1(new_n769_), .B2(new_n314_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT50), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n787_), .A2(new_n789_), .ZN(G1335gat));
  NOR2_X1   g589(.A1(new_n622_), .A2(new_n705_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n764_), .A2(new_n791_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(G85gat), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n793_), .A2(new_n794_), .A3(new_n677_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n622_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n796_));
  AND2_X1   g595(.A1(new_n729_), .A2(new_n796_), .ZN(new_n797_));
  AND2_X1   g596(.A1(new_n797_), .A2(KEYINPUT111), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(KEYINPUT111), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n798_), .A2(new_n799_), .A3(new_n451_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n795_), .B1(new_n800_), .B2(new_n794_), .ZN(new_n801_));
  XNOR2_X1  g600(.A(new_n801_), .B(KEYINPUT112), .ZN(G1336gat));
  INV_X1    g601(.A(G92gat), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n793_), .A2(new_n803_), .A3(new_n690_), .ZN(new_n804_));
  NOR3_X1   g603(.A1(new_n798_), .A2(new_n799_), .A3(new_n403_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n803_), .ZN(G1337gat));
  AOI21_X1  g605(.A(new_n558_), .B1(new_n797_), .B2(new_n429_), .ZN(new_n807_));
  NOR2_X1   g606(.A1(new_n483_), .A2(new_n545_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n807_), .B1(new_n793_), .B2(new_n808_), .ZN(new_n809_));
  XNOR2_X1  g608(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n809_), .B(new_n810_), .ZN(G1338gat));
  NAND3_X1  g610(.A1(new_n793_), .A2(new_n548_), .A3(new_n478_), .ZN(new_n812_));
  XNOR2_X1  g611(.A(new_n812_), .B(KEYINPUT114), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n729_), .A2(new_n478_), .A3(new_n796_), .ZN(new_n814_));
  AOI21_X1  g613(.A(KEYINPUT115), .B1(new_n814_), .B2(G106gat), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n813_), .A2(new_n817_), .ZN(new_n818_));
  AND3_X1   g617(.A1(new_n814_), .A2(KEYINPUT115), .A3(G106gat), .ZN(new_n819_));
  NOR3_X1   g618(.A1(new_n819_), .A2(new_n815_), .A3(new_n816_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n821_), .B(new_n822_), .ZN(G1339gat));
  NAND2_X1  g622(.A1(new_n674_), .A2(new_n533_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825_));
  XNOR2_X1  g624(.A(new_n824_), .B(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n599_), .A2(KEYINPUT55), .A3(new_n601_), .ZN(new_n827_));
  AND2_X1   g626(.A1(new_n596_), .A2(new_n598_), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n590_), .B1(new_n646_), .B2(new_n550_), .ZN(new_n829_));
  OAI21_X1  g628(.A(new_n606_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n827_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(KEYINPUT55), .B1(new_n599_), .B2(new_n601_), .ZN(new_n832_));
  OAI211_X1 g631(.A(KEYINPUT56), .B(new_n613_), .C1(new_n831_), .C2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT119), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n833_), .A2(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n613_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT56), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n602_), .A2(new_n839_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n840_), .A2(new_n830_), .A3(new_n827_), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n841_), .A2(KEYINPUT119), .A3(KEYINPUT56), .A4(new_n613_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n835_), .A2(new_n838_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n513_), .A2(new_n514_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n485_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n846_), .A3(new_n527_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n485_), .B1(new_n520_), .B2(KEYINPUT117), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(KEYINPUT117), .B2(new_n520_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n521_), .B1(new_n513_), .B2(new_n514_), .ZN(new_n850_));
  OAI21_X1  g649(.A(KEYINPUT116), .B1(new_n850_), .B2(new_n526_), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n847_), .A2(new_n849_), .A3(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT118), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(new_n854_));
  NAND4_X1  g653(.A1(new_n847_), .A2(new_n851_), .A3(new_n849_), .A4(KEYINPUT118), .ZN(new_n855_));
  AND4_X1   g654(.A1(new_n530_), .A2(new_n854_), .A3(new_n616_), .A4(new_n855_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n843_), .A2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT58), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n724_), .B1(new_n857_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n860_));
  NAND4_X1  g659(.A1(new_n843_), .A2(new_n856_), .A3(new_n860_), .A4(KEYINPUT58), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n843_), .A2(new_n856_), .A3(KEYINPUT58), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT120), .ZN(new_n863_));
  NAND3_X1  g662(.A1(new_n859_), .A2(new_n861_), .A3(new_n863_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n531_), .A2(new_n532_), .A3(new_n616_), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n838_), .B2(new_n833_), .ZN(new_n866_));
  AND4_X1   g665(.A1(new_n530_), .A2(new_n617_), .A3(new_n854_), .A4(new_n855_), .ZN(new_n867_));
  OAI21_X1  g666(.A(new_n714_), .B1(new_n866_), .B2(new_n867_), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT57), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n864_), .A2(new_n870_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n868_), .A2(new_n869_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n826_), .B1(new_n873_), .B2(new_n673_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n314_), .A2(new_n403_), .A3(new_n677_), .A4(new_n429_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(G113gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n682_), .ZN(new_n878_));
  OAI21_X1  g677(.A(KEYINPUT59), .B1(new_n874_), .B2(new_n875_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n872_), .B1(new_n871_), .B2(new_n880_), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n864_), .A2(KEYINPUT121), .A3(new_n870_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n683_), .B1(new_n881_), .B2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n883_), .A2(new_n826_), .ZN(new_n884_));
  OR2_X1    g683(.A1(new_n875_), .A2(KEYINPUT59), .ZN(new_n885_));
  OAI211_X1 g684(.A(new_n879_), .B(new_n682_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n878_), .B1(new_n887_), .B2(new_n877_), .ZN(G1340gat));
  INV_X1    g687(.A(G120gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n889_), .B1(new_n622_), .B2(KEYINPUT60), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n876_), .B(new_n890_), .C1(KEYINPUT60), .C2(new_n889_), .ZN(new_n891_));
  OAI211_X1 g690(.A(new_n879_), .B(new_n623_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n892_));
  INV_X1    g691(.A(new_n892_), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n891_), .B1(new_n893_), .B2(new_n889_), .ZN(G1341gat));
  INV_X1    g693(.A(G127gat), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n876_), .A2(new_n895_), .A3(new_n683_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n879_), .B(new_n683_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  OAI21_X1  g697(.A(new_n896_), .B1(new_n898_), .B2(new_n895_), .ZN(G1342gat));
  INV_X1    g698(.A(G134gat), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n876_), .A2(new_n900_), .A3(new_n654_), .ZN(new_n901_));
  OAI211_X1 g700(.A(new_n879_), .B(new_n659_), .C1(new_n884_), .C2(new_n885_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n902_), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n901_), .B1(new_n903_), .B2(new_n900_), .ZN(G1343gat));
  NOR2_X1   g703(.A1(new_n874_), .A2(new_n429_), .ZN(new_n905_));
  NOR3_X1   g704(.A1(new_n690_), .A2(new_n451_), .A3(new_n314_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n907_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n908_), .A2(new_n204_), .A3(new_n682_), .ZN(new_n909_));
  OAI21_X1  g708(.A(G141gat), .B1(new_n907_), .B2(new_n533_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n909_), .A2(new_n910_), .ZN(G1344gat));
  NAND3_X1  g710(.A1(new_n908_), .A2(new_n205_), .A3(new_n623_), .ZN(new_n912_));
  OAI21_X1  g711(.A(G148gat), .B1(new_n907_), .B2(new_n622_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(G1345gat));
  XNOR2_X1  g713(.A(KEYINPUT61), .B(G155gat), .ZN(new_n915_));
  OR3_X1    g714(.A1(new_n907_), .A2(new_n673_), .A3(new_n915_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n907_), .B2(new_n673_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1346gat));
  INV_X1    g717(.A(G162gat), .ZN(new_n919_));
  NOR2_X1   g718(.A1(new_n719_), .A2(new_n919_), .ZN(new_n920_));
  XOR2_X1   g719(.A(new_n920_), .B(KEYINPUT122), .Z(new_n921_));
  NAND3_X1  g720(.A1(new_n905_), .A2(new_n654_), .A3(new_n906_), .ZN(new_n922_));
  AOI22_X1  g721(.A1(new_n908_), .A2(new_n921_), .B1(new_n922_), .B2(new_n919_), .ZN(G1347gat));
  NOR3_X1   g722(.A1(new_n478_), .A2(new_n483_), .A3(new_n677_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n690_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n925_), .ZN(new_n926_));
  OAI211_X1 g725(.A(new_n682_), .B(new_n926_), .C1(new_n883_), .C2(new_n826_), .ZN(new_n927_));
  OAI211_X1 g726(.A(KEYINPUT62), .B(new_n342_), .C1(new_n927_), .C2(KEYINPUT22), .ZN(new_n928_));
  INV_X1    g727(.A(new_n928_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n927_), .A2(KEYINPUT62), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(new_n342_), .ZN(new_n931_));
  OAI21_X1  g730(.A(KEYINPUT62), .B1(new_n927_), .B2(KEYINPUT22), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n929_), .B1(new_n931_), .B2(new_n932_), .ZN(G1348gat));
  NOR2_X1   g732(.A1(new_n884_), .A2(new_n925_), .ZN(new_n934_));
  AOI21_X1  g733(.A(G176gat), .B1(new_n934_), .B2(new_n623_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n936_));
  NOR2_X1   g735(.A1(new_n874_), .A2(new_n925_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n622_), .A2(new_n343_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n936_), .B1(new_n937_), .B2(new_n938_), .ZN(new_n939_));
  AND3_X1   g738(.A1(new_n937_), .A2(new_n936_), .A3(new_n938_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n935_), .A2(new_n939_), .A3(new_n940_), .ZN(G1349gat));
  AOI21_X1  g740(.A(G183gat), .B1(new_n937_), .B2(new_n683_), .ZN(new_n942_));
  NAND2_X1  g741(.A1(new_n352_), .A2(new_n351_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n683_), .A2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n942_), .B1(new_n934_), .B2(new_n945_), .ZN(G1350gat));
  NAND3_X1  g745(.A1(new_n934_), .A2(new_n349_), .A3(new_n654_), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n659_), .B(new_n926_), .C1(new_n883_), .C2(new_n826_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT124), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n948_), .A2(new_n949_), .A3(G190gat), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n949_), .B1(new_n948_), .B2(G190gat), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n947_), .B1(new_n950_), .B2(new_n951_), .ZN(G1351gat));
  NAND3_X1  g751(.A1(new_n690_), .A2(new_n451_), .A3(new_n478_), .ZN(new_n953_));
  NOR3_X1   g752(.A1(new_n874_), .A2(new_n429_), .A3(new_n953_), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n954_), .A2(new_n682_), .ZN(new_n955_));
  XNOR2_X1  g754(.A(new_n955_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g755(.A1(new_n954_), .A2(new_n623_), .ZN(new_n957_));
  XNOR2_X1  g756(.A(new_n957_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n683_), .B1(new_n959_), .B2(new_n248_), .ZN(new_n960_));
  XOR2_X1   g759(.A(new_n960_), .B(KEYINPUT125), .Z(new_n961_));
  INV_X1    g760(.A(KEYINPUT126), .ZN(new_n962_));
  OAI21_X1  g761(.A(new_n962_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n963_));
  NAND3_X1  g762(.A1(new_n959_), .A2(new_n248_), .A3(KEYINPUT126), .ZN(new_n964_));
  AOI22_X1  g763(.A1(new_n954_), .A2(new_n961_), .B1(new_n963_), .B2(new_n964_), .ZN(new_n965_));
  AND2_X1   g764(.A1(new_n954_), .A2(new_n961_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n965_), .B1(new_n966_), .B2(new_n964_), .ZN(G1354gat));
  NAND2_X1  g766(.A1(new_n954_), .A2(new_n654_), .ZN(new_n968_));
  XNOR2_X1  g767(.A(KEYINPUT127), .B(G218gat), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n724_), .A2(new_n969_), .ZN(new_n970_));
  AOI22_X1  g769(.A1(new_n968_), .A2(new_n969_), .B1(new_n954_), .B2(new_n970_), .ZN(G1355gat));
endmodule


