//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n891_, new_n892_, new_n893_,
    new_n894_, new_n896_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n916_, new_n917_,
    new_n918_, new_n920_, new_n921_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n942_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT18), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204_));
  XOR2_X1   g003(.A(new_n203_), .B(new_n204_), .Z(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XNOR2_X1  g005(.A(G197gat), .B(G204gat), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT21), .ZN(new_n208_));
  NOR2_X1   g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(G218gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(G211gat), .ZN(new_n211_));
  INV_X1    g010(.A(G211gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(G218gat), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n211_), .A2(new_n213_), .A3(KEYINPUT91), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT91), .ZN(new_n215_));
  NOR2_X1   g014(.A1(new_n212_), .A2(G218gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n210_), .A2(G211gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n215_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n209_), .A2(new_n214_), .A3(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n214_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT89), .ZN(new_n221_));
  INV_X1    g020(.A(G197gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n221_), .B1(new_n222_), .B2(G204gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n222_), .A2(G204gat), .ZN(new_n224_));
  INV_X1    g023(.A(G204gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n225_), .A2(KEYINPUT89), .A3(G197gat), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n223_), .A2(new_n224_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT21), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n220_), .A2(new_n228_), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT90), .B1(new_n207_), .B2(new_n208_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n225_), .A2(G197gat), .ZN(new_n231_));
  AND4_X1   g030(.A1(KEYINPUT90), .A2(new_n231_), .A3(new_n224_), .A4(new_n208_), .ZN(new_n232_));
  NOR2_X1   g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n219_), .B1(new_n229_), .B2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT23), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n236_), .A2(G183gat), .A3(G190gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(G183gat), .A2(G190gat), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT23), .ZN(new_n241_));
  NAND4_X1  g040(.A1(new_n236_), .A2(KEYINPUT80), .A3(G183gat), .A4(G190gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(new_n239_), .A2(new_n241_), .A3(new_n242_), .ZN(new_n243_));
  NOR3_X1   g042(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(G169gat), .A2(G176gat), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n245_), .A2(KEYINPUT24), .ZN(new_n246_));
  INV_X1    g045(.A(G169gat), .ZN(new_n247_));
  INV_X1    g046(.A(G176gat), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n244_), .B1(new_n246_), .B2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT26), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(G190gat), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n252_), .A2(KEYINPUT79), .ZN(new_n253_));
  INV_X1    g052(.A(G190gat), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT26), .ZN(new_n255_));
  INV_X1    g054(.A(G183gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT25), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n253_), .A2(new_n255_), .A3(new_n257_), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT78), .B1(new_n256_), .B2(KEYINPUT25), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT78), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT25), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n260_), .A2(new_n261_), .A3(G183gat), .ZN(new_n262_));
  OAI211_X1 g061(.A(new_n259_), .B(new_n262_), .C1(KEYINPUT79), .C2(new_n252_), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n243_), .B(new_n250_), .C1(new_n258_), .C2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(KEYINPUT81), .B(G169gat), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT22), .ZN(new_n266_));
  OAI21_X1  g065(.A(KEYINPUT82), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n247_), .A2(KEYINPUT81), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT81), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G169gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n268_), .A2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(new_n272_), .A3(KEYINPUT22), .ZN(new_n273_));
  AOI21_X1  g072(.A(G176gat), .B1(new_n266_), .B2(G169gat), .ZN(new_n274_));
  AND3_X1   g073(.A1(new_n267_), .A2(new_n273_), .A3(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n241_), .A2(new_n237_), .A3(KEYINPUT83), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n256_), .A2(new_n254_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT83), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n278_), .A2(new_n236_), .A3(G183gat), .A4(G190gat), .ZN(new_n279_));
  NAND3_X1  g078(.A1(new_n276_), .A2(new_n277_), .A3(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n280_), .A2(new_n245_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n264_), .B1(new_n275_), .B2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT84), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n266_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n274_), .B1(new_n284_), .B2(new_n272_), .ZN(new_n285_));
  NOR3_X1   g084(.A1(new_n265_), .A2(KEYINPUT82), .A3(new_n266_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n280_), .B(new_n245_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT84), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n287_), .A2(new_n288_), .A3(new_n264_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n235_), .B1(new_n283_), .B2(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G226gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n291_), .B(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n243_), .A2(new_n277_), .ZN(new_n294_));
  XNOR2_X1  g093(.A(KEYINPUT22), .B(G169gat), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT94), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n245_), .A2(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(KEYINPUT94), .A2(G169gat), .A3(G176gat), .ZN(new_n298_));
  AOI22_X1  g097(.A1(new_n295_), .A2(new_n248_), .B1(new_n297_), .B2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n261_), .A2(G183gat), .ZN(new_n301_));
  NAND4_X1  g100(.A1(new_n252_), .A2(new_n255_), .A3(new_n257_), .A4(new_n301_), .ZN(new_n302_));
  NAND4_X1  g101(.A1(new_n302_), .A2(new_n279_), .A3(new_n276_), .A4(new_n250_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT20), .B1(new_n304_), .B2(new_n234_), .ZN(new_n305_));
  NOR3_X1   g104(.A1(new_n290_), .A2(new_n293_), .A3(new_n305_), .ZN(new_n306_));
  INV_X1    g105(.A(new_n293_), .ZN(new_n307_));
  NAND3_X1  g106(.A1(new_n283_), .A2(new_n289_), .A3(new_n235_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT20), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n309_), .B1(new_n304_), .B2(new_n234_), .ZN(new_n310_));
  AOI21_X1  g109(.A(new_n307_), .B1(new_n308_), .B2(new_n310_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n206_), .B1(new_n306_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT95), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n287_), .A2(new_n288_), .A3(new_n264_), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n288_), .B1(new_n287_), .B2(new_n264_), .ZN(new_n315_));
  NOR3_X1   g114(.A1(new_n314_), .A2(new_n315_), .A3(new_n234_), .ZN(new_n316_));
  INV_X1    g115(.A(new_n310_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n293_), .B1(new_n316_), .B2(new_n317_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n234_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n305_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n319_), .A2(new_n307_), .A3(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n318_), .A2(new_n205_), .A3(new_n321_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n312_), .A2(new_n313_), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT27), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n318_), .A2(new_n321_), .ZN(new_n325_));
  NAND3_X1  g124(.A1(new_n325_), .A2(KEYINPUT95), .A3(new_n206_), .ZN(new_n326_));
  NAND3_X1  g125(.A1(new_n323_), .A2(new_n324_), .A3(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT97), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n293_), .B1(new_n290_), .B2(new_n305_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n308_), .A2(new_n310_), .A3(new_n307_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n328_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n319_), .A2(new_n320_), .ZN(new_n332_));
  AOI21_X1  g131(.A(KEYINPUT97), .B1(new_n332_), .B2(new_n293_), .ZN(new_n333_));
  OAI21_X1  g132(.A(new_n206_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n334_));
  AND2_X1   g133(.A1(new_n322_), .A2(KEYINPUT27), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  AND2_X1   g135(.A1(new_n327_), .A2(new_n336_), .ZN(new_n337_));
  AOI21_X1  g136(.A(KEYINPUT92), .B1(G228gat), .B2(G233gat), .ZN(new_n338_));
  AND3_X1   g137(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n339_));
  AOI21_X1  g138(.A(KEYINPUT87), .B1(G155gat), .B2(G162gat), .ZN(new_n340_));
  OAI21_X1  g139(.A(KEYINPUT1), .B1(new_n339_), .B2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(G155gat), .A2(G162gat), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT87), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT1), .ZN(new_n345_));
  NAND3_X1  g144(.A1(KEYINPUT87), .A2(G155gat), .A3(G162gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n344_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  INV_X1    g146(.A(G155gat), .ZN(new_n348_));
  INV_X1    g147(.A(G162gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n341_), .A2(new_n347_), .A3(new_n350_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(G141gat), .A2(G148gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(G141gat), .A2(G148gat), .ZN(new_n354_));
  AND2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n351_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(G141gat), .ZN(new_n357_));
  INV_X1    g156(.A(G148gat), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n357_), .A2(new_n358_), .A3(KEYINPUT88), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT3), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n352_), .A2(KEYINPUT88), .A3(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT2), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n354_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n365_));
  NAND4_X1  g164(.A1(new_n360_), .A2(new_n362_), .A3(new_n364_), .A4(new_n365_), .ZN(new_n366_));
  AOI22_X1  g165(.A1(new_n344_), .A2(new_n346_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n356_), .A2(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT28), .B1(new_n369_), .B2(KEYINPUT29), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n369_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n338_), .B1(new_n371_), .B2(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n372_), .ZN(new_n374_));
  INV_X1    g173(.A(new_n338_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n374_), .A2(new_n370_), .A3(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(G106gat), .ZN(new_n378_));
  NAND3_X1  g177(.A1(KEYINPUT92), .A2(G228gat), .A3(G233gat), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n220_), .B(new_n228_), .C1(new_n230_), .C2(new_n232_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n380_), .B1(new_n381_), .B2(new_n219_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n369_), .A2(KEYINPUT29), .ZN(new_n383_));
  INV_X1    g182(.A(G78gat), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n384_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n378_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n234_), .A2(new_n379_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT29), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n389_), .B1(new_n356_), .B2(new_n368_), .ZN(new_n390_));
  OAI21_X1  g189(.A(G78gat), .B1(new_n388_), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n382_), .A2(new_n383_), .A3(new_n384_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n391_), .A2(G106gat), .A3(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(G22gat), .B(G50gat), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n387_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n395_), .B1(new_n387_), .B2(new_n393_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n377_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NOR3_X1   g197(.A1(new_n385_), .A2(new_n386_), .A3(new_n378_), .ZN(new_n399_));
  AOI21_X1  g198(.A(G106gat), .B1(new_n391_), .B2(new_n392_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n394_), .B1(new_n399_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n377_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n387_), .A2(new_n393_), .A3(new_n395_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n398_), .A2(new_n404_), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G1gat), .B(G29gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n406_), .B(G85gat), .ZN(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT0), .B(G57gat), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT96), .ZN(new_n410_));
  INV_X1    g209(.A(G134gat), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(G127gat), .ZN(new_n412_));
  INV_X1    g211(.A(G127gat), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n413_), .A2(G134gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n412_), .A2(new_n414_), .A3(KEYINPUT85), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G113gat), .B(G120gat), .ZN(new_n419_));
  AND3_X1   g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n419_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n421_));
  NOR2_X1   g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n422_), .A2(new_n369_), .ZN(new_n423_));
  OAI211_X1 g222(.A(new_n356_), .B(new_n368_), .C1(new_n420_), .C2(new_n421_), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n423_), .A2(KEYINPUT4), .A3(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n422_), .A2(new_n369_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(G225gat), .A2(G233gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n427_), .A2(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n410_), .B1(new_n425_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n431_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n423_), .A2(KEYINPUT4), .A3(new_n424_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n433_), .A2(KEYINPUT96), .A3(new_n429_), .A4(new_n427_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n423_), .A2(new_n424_), .A3(new_n428_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n409_), .B1(new_n432_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n409_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n431_), .A2(new_n438_), .A3(new_n435_), .A4(new_n434_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G71gat), .B(G99gat), .ZN(new_n442_));
  INV_X1    g241(.A(G43gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT30), .ZN(new_n445_));
  OR2_X1    g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n444_), .A2(new_n445_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(G227gat), .A2(G233gat), .ZN(new_n448_));
  INV_X1    g247(.A(G15gat), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n448_), .B(new_n449_), .ZN(new_n450_));
  AND3_X1   g249(.A1(new_n446_), .A2(new_n447_), .A3(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n450_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n453_), .A2(new_n283_), .A3(new_n289_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT86), .ZN(new_n455_));
  OAI22_X1  g254(.A1(new_n451_), .A2(new_n452_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(new_n455_), .A3(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT31), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT31), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n454_), .A2(new_n455_), .A3(new_n459_), .A4(new_n456_), .ZN(new_n460_));
  AND3_X1   g259(.A1(new_n458_), .A2(new_n422_), .A3(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n422_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n462_));
  NOR2_X1   g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  AND4_X1   g262(.A1(new_n337_), .A2(new_n405_), .A3(new_n441_), .A4(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n323_), .A2(new_n326_), .ZN(new_n465_));
  AND3_X1   g264(.A1(new_n423_), .A2(new_n424_), .A3(new_n429_), .ZN(new_n466_));
  AND2_X1   g265(.A1(new_n427_), .A2(new_n428_), .ZN(new_n467_));
  AOI211_X1 g266(.A(new_n438_), .B(new_n466_), .C1(new_n433_), .C2(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n436_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT33), .ZN(new_n470_));
  NAND4_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n438_), .A4(new_n431_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n439_), .A2(KEYINPUT33), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n468_), .B1(new_n471_), .B2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n465_), .A2(new_n473_), .ZN(new_n474_));
  AND2_X1   g273(.A1(new_n205_), .A2(KEYINPUT32), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n475_), .B1(new_n331_), .B2(new_n333_), .ZN(new_n476_));
  OAI211_X1 g275(.A(new_n476_), .B(new_n440_), .C1(new_n325_), .C2(new_n475_), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n474_), .A2(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n405_), .ZN(new_n479_));
  NOR3_X1   g278(.A1(new_n396_), .A2(new_n397_), .A3(new_n377_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n402_), .B1(new_n401_), .B2(new_n403_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n482_), .A2(new_n327_), .A3(new_n336_), .A4(new_n441_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(KEYINPUT98), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n405_), .A2(new_n440_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT98), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n327_), .A4(new_n336_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n479_), .A2(new_n484_), .A3(new_n487_), .ZN(new_n488_));
  INV_X1    g287(.A(new_n463_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n464_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G29gat), .B(G36gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G43gat), .B(G50gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n491_), .B(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n493_), .B(KEYINPUT15), .ZN(new_n494_));
  XNOR2_X1  g293(.A(G1gat), .B(G8gat), .ZN(new_n495_));
  OR2_X1    g294(.A1(new_n495_), .A2(KEYINPUT75), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(KEYINPUT75), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  XNOR2_X1  g297(.A(G15gat), .B(G22gat), .ZN(new_n499_));
  INV_X1    g298(.A(G1gat), .ZN(new_n500_));
  INV_X1    g299(.A(G8gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT14), .B1(new_n500_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n499_), .A2(new_n502_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n498_), .A2(new_n503_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n496_), .A2(new_n502_), .A3(new_n499_), .A4(new_n497_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(new_n494_), .A2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508_));
  INV_X1    g307(.A(new_n493_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n507_), .B(new_n508_), .C1(new_n506_), .C2(new_n509_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n504_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n509_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n512_));
  OAI211_X1 g311(.A(G229gat), .B(G233gat), .C1(new_n511_), .C2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n510_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G113gat), .B(G141gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(G169gat), .B(G197gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(new_n515_), .B(new_n516_), .Z(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n514_), .B(new_n518_), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n519_), .B(KEYINPUT77), .Z(new_n520_));
  NOR2_X1   g319(.A1(new_n490_), .A2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(G231gat), .A2(G233gat), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n506_), .B(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(G71gat), .B(G78gat), .Z(new_n524_));
  XNOR2_X1  g323(.A(G57gat), .B(G64gat), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n524_), .B1(KEYINPUT11), .B2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT68), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n525_), .A2(new_n527_), .A3(KEYINPUT11), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n527_), .B1(new_n525_), .B2(KEYINPUT11), .ZN(new_n529_));
  OR3_X1    g328(.A1(new_n526_), .A2(new_n528_), .A3(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n526_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n523_), .B(new_n532_), .ZN(new_n533_));
  XOR2_X1   g332(.A(G127gat), .B(G155gat), .Z(new_n534_));
  XNOR2_X1  g333(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n534_), .B(new_n535_), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G183gat), .B(G211gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT17), .ZN(new_n539_));
  OAI21_X1  g338(.A(KEYINPUT69), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n533_), .A2(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n541_), .B1(new_n539_), .B2(new_n538_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n533_), .A2(new_n540_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT37), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G190gat), .B(G218gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G134gat), .B(G162gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n548_), .B(KEYINPUT36), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G99gat), .A2(G106gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(G99gat), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT7), .ZN(new_n555_));
  OAI211_X1 g354(.A(new_n554_), .B(new_n378_), .C1(new_n555_), .C2(KEYINPUT67), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT67), .ZN(new_n557_));
  OAI21_X1  g356(.A(new_n556_), .B1(new_n557_), .B2(KEYINPUT7), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n555_), .A2(new_n554_), .A3(new_n378_), .A4(KEYINPUT67), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n553_), .A2(new_n558_), .A3(new_n559_), .ZN(new_n560_));
  XOR2_X1   g359(.A(G85gat), .B(G92gat), .Z(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT8), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT8), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n560_), .A2(new_n564_), .A3(new_n561_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(KEYINPUT9), .A2(G85gat), .ZN(new_n566_));
  XNOR2_X1  g365(.A(KEYINPUT64), .B(G85gat), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT9), .ZN(new_n568_));
  AND2_X1   g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(G92gat), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n566_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n566_), .A2(new_n570_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT65), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT10), .B(G99gat), .ZN(new_n575_));
  OR2_X1    g374(.A1(new_n575_), .A2(G106gat), .ZN(new_n576_));
  AND2_X1   g375(.A1(new_n553_), .A2(new_n576_), .ZN(new_n577_));
  AOI22_X1  g376(.A1(new_n563_), .A2(new_n565_), .B1(new_n574_), .B2(new_n577_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n578_), .A2(new_n493_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n577_), .A2(new_n574_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n565_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n564_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n580_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n583_), .A2(new_n494_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n585_));
  NAND2_X1  g384(.A1(G232gat), .A2(G233gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT35), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n579_), .A2(new_n584_), .A3(new_n590_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n588_), .A2(new_n589_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n592_), .ZN(new_n594_));
  NAND4_X1  g393(.A1(new_n579_), .A2(new_n584_), .A3(new_n594_), .A4(new_n590_), .ZN(new_n595_));
  AOI21_X1  g394(.A(new_n550_), .B1(new_n593_), .B2(new_n595_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n548_), .A2(KEYINPUT36), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n593_), .A2(new_n598_), .A3(new_n595_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n545_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n599_), .ZN(new_n601_));
  NOR3_X1   g400(.A1(new_n601_), .A2(new_n596_), .A3(KEYINPUT37), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n544_), .B1(new_n600_), .B2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT12), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n530_), .A2(KEYINPUT69), .A3(new_n531_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  AOI21_X1  g405(.A(KEYINPUT69), .B1(new_n530_), .B2(new_n531_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n604_), .B1(new_n608_), .B2(new_n578_), .ZN(new_n609_));
  INV_X1    g408(.A(G230gat), .ZN(new_n610_));
  INV_X1    g409(.A(G233gat), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n608_), .A2(new_n578_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n532_), .A2(new_n604_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n583_), .A2(new_n615_), .ZN(new_n616_));
  NAND4_X1  g415(.A1(new_n609_), .A2(new_n613_), .A3(new_n614_), .A4(new_n616_), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n608_), .A2(new_n578_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n607_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(new_n605_), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(new_n583_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n612_), .B1(new_n618_), .B2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n617_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT70), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT72), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n617_), .A2(new_n622_), .A3(KEYINPUT70), .ZN(new_n627_));
  XOR2_X1   g426(.A(G120gat), .B(G148gat), .Z(new_n628_));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n628_), .B(new_n629_), .ZN(new_n630_));
  XNOR2_X1  g429(.A(KEYINPUT71), .B(KEYINPUT5), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n630_), .B(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n625_), .A2(new_n626_), .A3(new_n627_), .A4(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n617_), .A2(new_n622_), .A3(new_n632_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n632_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n637_));
  AOI21_X1  g436(.A(new_n626_), .B1(new_n637_), .B2(new_n627_), .ZN(new_n638_));
  INV_X1    g437(.A(KEYINPUT13), .ZN(new_n639_));
  AND2_X1   g438(.A1(new_n639_), .A2(KEYINPUT73), .ZN(new_n640_));
  NOR2_X1   g439(.A1(new_n639_), .A2(KEYINPUT73), .ZN(new_n641_));
  OAI22_X1  g440(.A1(new_n636_), .A2(new_n638_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n637_), .A2(new_n627_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT72), .ZN(new_n644_));
  INV_X1    g443(.A(new_n641_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n644_), .A2(new_n635_), .A3(new_n634_), .A4(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n603_), .B1(new_n642_), .B2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n521_), .A2(new_n647_), .ZN(new_n648_));
  NOR3_X1   g447(.A1(new_n648_), .A2(G1gat), .A3(new_n441_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT99), .ZN(new_n650_));
  OR2_X1    g449(.A1(new_n650_), .A2(KEYINPUT38), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n650_), .A2(KEYINPUT38), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n601_), .A2(new_n596_), .ZN(new_n653_));
  NOR2_X1   g452(.A1(new_n490_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n519_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n544_), .ZN(new_n656_));
  AOI211_X1 g455(.A(new_n655_), .B(new_n656_), .C1(new_n642_), .C2(new_n646_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n654_), .A2(new_n657_), .ZN(new_n658_));
  OR2_X1    g457(.A1(new_n658_), .A2(KEYINPUT100), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(KEYINPUT100), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n441_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n661_));
  OAI211_X1 g460(.A(new_n651_), .B(new_n652_), .C1(new_n500_), .C2(new_n661_), .ZN(G1324gat));
  INV_X1    g461(.A(new_n337_), .ZN(new_n663_));
  NAND4_X1  g462(.A1(new_n521_), .A2(new_n501_), .A3(new_n663_), .A4(new_n647_), .ZN(new_n664_));
  NOR2_X1   g463(.A1(new_n658_), .A2(new_n337_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n501_), .B1(new_n665_), .B2(KEYINPUT101), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT39), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT101), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n668_), .B1(new_n658_), .B2(new_n337_), .ZN(new_n669_));
  AND3_X1   g468(.A1(new_n666_), .A2(new_n667_), .A3(new_n669_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n667_), .B1(new_n666_), .B2(new_n669_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n664_), .B1(new_n670_), .B2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT40), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(KEYINPUT40), .B(new_n664_), .C1(new_n670_), .C2(new_n671_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1325gat));
  NAND2_X1  g475(.A1(new_n659_), .A2(new_n660_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n677_), .A2(new_n463_), .ZN(new_n678_));
  AND3_X1   g477(.A1(new_n678_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(KEYINPUT41), .B1(new_n678_), .B2(G15gat), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n463_), .A2(new_n449_), .ZN(new_n681_));
  OAI22_X1  g480(.A1(new_n679_), .A2(new_n680_), .B1(new_n648_), .B2(new_n681_), .ZN(G1326gat));
  AOI21_X1  g481(.A(new_n405_), .B1(new_n659_), .B2(new_n660_), .ZN(new_n683_));
  INV_X1    g482(.A(G22gat), .ZN(new_n684_));
  OR2_X1    g483(.A1(new_n683_), .A2(new_n684_), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n685_), .A2(KEYINPUT42), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(KEYINPUT42), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n482_), .A2(new_n684_), .ZN(new_n688_));
  OAI22_X1  g487(.A1(new_n686_), .A2(new_n687_), .B1(new_n648_), .B2(new_n688_), .ZN(G1327gat));
  INV_X1    g488(.A(new_n602_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT37), .B1(new_n601_), .B2(new_n596_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT43), .B1(new_n490_), .B2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n600_), .A2(new_n602_), .ZN(new_n695_));
  AOI22_X1  g494(.A1(new_n405_), .A2(new_n478_), .B1(new_n483_), .B2(KEYINPUT98), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n463_), .B1(new_n696_), .B2(new_n487_), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n694_), .B(new_n695_), .C1(new_n697_), .C2(new_n464_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n693_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n642_), .A2(new_n646_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n700_), .A2(new_n519_), .A3(new_n656_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(KEYINPUT44), .B1(new_n699_), .B2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT44), .ZN(new_n704_));
  AOI211_X1 g503(.A(new_n704_), .B(new_n701_), .C1(new_n693_), .C2(new_n698_), .ZN(new_n705_));
  NOR3_X1   g504(.A1(new_n703_), .A2(new_n705_), .A3(new_n441_), .ZN(new_n706_));
  INV_X1    g505(.A(G29gat), .ZN(new_n707_));
  INV_X1    g506(.A(new_n653_), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n708_), .A2(new_n544_), .ZN(new_n709_));
  AND2_X1   g508(.A1(new_n700_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n521_), .A2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n440_), .A2(new_n707_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT102), .ZN(new_n713_));
  OAI22_X1  g512(.A1(new_n706_), .A2(new_n707_), .B1(new_n711_), .B2(new_n713_), .ZN(G1328gat));
  INV_X1    g513(.A(KEYINPUT46), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n715_), .A2(KEYINPUT103), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT104), .Z(new_n717_));
  INV_X1    g516(.A(new_n717_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n337_), .A2(G36gat), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n719_), .B1(new_n711_), .B2(new_n721_), .ZN(new_n722_));
  NAND4_X1  g521(.A1(new_n521_), .A2(KEYINPUT45), .A3(new_n710_), .A4(new_n720_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n722_), .A2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n699_), .A2(new_n702_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n725_), .A2(new_n704_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n699_), .A2(KEYINPUT44), .A3(new_n702_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n726_), .A2(new_n663_), .A3(new_n727_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n724_), .B1(new_n728_), .B2(G36gat), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n715_), .A2(KEYINPUT103), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n718_), .B1(new_n729_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n730_), .ZN(new_n732_));
  INV_X1    g531(.A(G36gat), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n703_), .A2(new_n705_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n733_), .B1(new_n734_), .B2(new_n663_), .ZN(new_n735_));
  OAI211_X1 g534(.A(new_n732_), .B(new_n717_), .C1(new_n735_), .C2(new_n724_), .ZN(new_n736_));
  AND2_X1   g535(.A1(new_n731_), .A2(new_n736_), .ZN(G1329gat));
  NAND3_X1  g536(.A1(new_n734_), .A2(G43gat), .A3(new_n463_), .ZN(new_n738_));
  OAI21_X1  g537(.A(new_n443_), .B1(new_n711_), .B2(new_n489_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g540(.A1(new_n734_), .A2(G50gat), .A3(new_n482_), .ZN(new_n742_));
  INV_X1    g541(.A(G50gat), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n743_), .B1(new_n711_), .B2(new_n405_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n742_), .A2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(G1331gat));
  INV_X1    g546(.A(G57gat), .ZN(new_n748_));
  INV_X1    g547(.A(new_n520_), .ZN(new_n749_));
  NOR3_X1   g548(.A1(new_n700_), .A2(new_n749_), .A3(new_n656_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n654_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n654_), .A2(KEYINPUT106), .A3(new_n750_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n748_), .B1(new_n755_), .B2(new_n440_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n490_), .A2(new_n519_), .ZN(new_n757_));
  INV_X1    g556(.A(new_n700_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n603_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n757_), .A2(new_n758_), .A3(new_n759_), .ZN(new_n760_));
  NOR3_X1   g559(.A1(new_n760_), .A2(G57gat), .A3(new_n441_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n756_), .A2(new_n761_), .ZN(G1332gat));
  OR3_X1    g561(.A1(new_n760_), .A2(G64gat), .A3(new_n337_), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n753_), .A2(new_n663_), .A3(new_n754_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT48), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n764_), .A2(new_n765_), .A3(G64gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n764_), .B2(G64gat), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n763_), .B1(new_n766_), .B2(new_n767_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT107), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n768_), .B(new_n769_), .ZN(G1333gat));
  INV_X1    g569(.A(KEYINPUT49), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n755_), .A2(new_n463_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n772_), .B2(G71gat), .ZN(new_n773_));
  INV_X1    g572(.A(G71gat), .ZN(new_n774_));
  AOI211_X1 g573(.A(KEYINPUT49), .B(new_n774_), .C1(new_n755_), .C2(new_n463_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n463_), .A2(new_n774_), .ZN(new_n776_));
  OAI22_X1  g575(.A1(new_n773_), .A2(new_n775_), .B1(new_n760_), .B2(new_n776_), .ZN(G1334gat));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n755_), .A2(new_n482_), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n778_), .B1(new_n779_), .B2(G78gat), .ZN(new_n780_));
  AOI211_X1 g579(.A(KEYINPUT50), .B(new_n384_), .C1(new_n755_), .C2(new_n482_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n482_), .A2(new_n384_), .ZN(new_n782_));
  OAI22_X1  g581(.A1(new_n780_), .A2(new_n781_), .B1(new_n760_), .B2(new_n782_), .ZN(G1335gat));
  NAND3_X1  g582(.A1(new_n757_), .A2(new_n758_), .A3(new_n709_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  AOI21_X1  g584(.A(G85gat), .B1(new_n785_), .B2(new_n440_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n642_), .A2(new_n646_), .A3(new_n655_), .A4(new_n656_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n787_), .B1(new_n693_), .B2(new_n698_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n788_), .ZN(new_n789_));
  AND2_X1   g588(.A1(new_n789_), .A2(KEYINPUT108), .ZN(new_n790_));
  NOR2_X1   g589(.A1(new_n789_), .A2(KEYINPUT108), .ZN(new_n791_));
  NOR2_X1   g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n441_), .A2(new_n567_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n786_), .B1(new_n792_), .B2(new_n793_), .ZN(G1336gat));
  NAND3_X1  g593(.A1(new_n785_), .A2(new_n570_), .A3(new_n663_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n790_), .A2(new_n791_), .A3(new_n337_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n795_), .B1(new_n796_), .B2(new_n570_), .ZN(G1337gat));
  OAI21_X1  g596(.A(G99gat), .B1(new_n789_), .B2(new_n489_), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n489_), .A2(new_n575_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n784_), .B2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(KEYINPUT109), .A2(KEYINPUT51), .ZN(new_n801_));
  XOR2_X1   g600(.A(new_n800_), .B(new_n801_), .Z(G1338gat));
  NAND3_X1  g601(.A1(new_n785_), .A2(new_n378_), .A3(new_n482_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804_));
  AOI211_X1 g603(.A(new_n405_), .B(new_n787_), .C1(new_n693_), .C2(new_n698_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n378_), .B1(new_n805_), .B2(KEYINPUT110), .ZN(new_n806_));
  AOI21_X1  g605(.A(KEYINPUT110), .B1(new_n788_), .B2(new_n482_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n804_), .B1(new_n806_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n787_), .ZN(new_n810_));
  NAND4_X1  g609(.A1(new_n699_), .A2(KEYINPUT110), .A3(new_n482_), .A4(new_n810_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(G106gat), .ZN(new_n812_));
  NOR3_X1   g611(.A1(new_n812_), .A2(new_n807_), .A3(KEYINPUT52), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n803_), .B1(new_n809_), .B2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(KEYINPUT53), .ZN(new_n815_));
  INV_X1    g614(.A(KEYINPUT53), .ZN(new_n816_));
  OAI211_X1 g615(.A(new_n816_), .B(new_n803_), .C1(new_n809_), .C2(new_n813_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n815_), .A2(new_n817_), .ZN(G1339gat));
  NOR4_X1   g617(.A1(new_n663_), .A2(new_n489_), .A3(new_n482_), .A4(new_n441_), .ZN(new_n819_));
  INV_X1    g618(.A(new_n819_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n510_), .A2(new_n513_), .A3(new_n517_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n508_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n518_), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n823_), .A2(KEYINPUT114), .ZN(new_n824_));
  NOR2_X1   g623(.A1(new_n512_), .A2(new_n508_), .ZN(new_n825_));
  AOI22_X1  g624(.A1(new_n823_), .A2(KEYINPUT114), .B1(new_n507_), .B2(new_n825_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n821_), .B1(new_n824_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n635_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT115), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n635_), .A2(new_n827_), .A3(KEYINPUT115), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833_));
  NAND2_X1  g632(.A1(new_n617_), .A2(new_n833_), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n609_), .A2(KEYINPUT55), .A3(new_n614_), .A4(new_n616_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n613_), .A2(KEYINPUT113), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n834_), .A2(new_n835_), .A3(new_n837_), .ZN(new_n838_));
  AND4_X1   g637(.A1(KEYINPUT55), .A2(new_n609_), .A3(new_n614_), .A4(new_n616_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n632_), .B1(new_n839_), .B2(new_n836_), .ZN(new_n840_));
  AND3_X1   g639(.A1(new_n838_), .A2(new_n840_), .A3(KEYINPUT56), .ZN(new_n841_));
  AOI21_X1  g640(.A(KEYINPUT56), .B1(new_n838_), .B2(new_n840_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n832_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT58), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n832_), .B(KEYINPUT58), .C1(new_n841_), .C2(new_n842_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n845_), .A2(new_n695_), .A3(new_n846_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n827_), .B1(new_n636_), .B2(new_n638_), .ZN(new_n848_));
  AND3_X1   g647(.A1(new_n635_), .A2(new_n519_), .A3(KEYINPUT112), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT112), .B1(new_n635_), .B2(new_n519_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n849_), .A2(new_n850_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n851_), .B1(new_n841_), .B2(new_n842_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n653_), .B1(new_n848_), .B2(new_n852_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n847_), .B1(new_n853_), .B2(KEYINPUT57), .ZN(new_n854_));
  AND2_X1   g653(.A1(new_n853_), .A2(KEYINPUT57), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n656_), .B1(new_n854_), .B2(new_n855_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(KEYINPUT111), .B(KEYINPUT54), .ZN(new_n857_));
  AND4_X1   g656(.A1(new_n520_), .A2(new_n700_), .A3(new_n759_), .A4(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n857_), .B1(new_n647_), .B2(new_n520_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AOI21_X1  g659(.A(new_n820_), .B1(new_n856_), .B2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(G113gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n861_), .A2(new_n862_), .A3(new_n519_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n856_), .A2(new_n860_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n864_), .A2(KEYINPUT116), .A3(new_n819_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n861_), .A2(KEYINPUT116), .A3(KEYINPUT59), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n520_), .B1(new_n867_), .B2(new_n868_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n863_), .B1(new_n869_), .B2(new_n862_), .ZN(G1340gat));
  XNOR2_X1  g669(.A(KEYINPUT117), .B(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(new_n700_), .B2(KEYINPUT60), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n861_), .B(new_n872_), .C1(KEYINPUT60), .C2(new_n871_), .ZN(new_n873_));
  AND4_X1   g672(.A1(KEYINPUT116), .A2(new_n864_), .A3(KEYINPUT59), .A4(new_n819_), .ZN(new_n874_));
  AOI21_X1  g673(.A(KEYINPUT59), .B1(new_n861_), .B2(KEYINPUT116), .ZN(new_n875_));
  OAI211_X1 g674(.A(KEYINPUT118), .B(new_n758_), .C1(new_n874_), .C2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(new_n871_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n867_), .A2(new_n868_), .ZN(new_n879_));
  AOI21_X1  g678(.A(KEYINPUT118), .B1(new_n879_), .B2(new_n758_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n873_), .B1(new_n878_), .B2(new_n880_), .ZN(G1341gat));
  AOI21_X1  g680(.A(G127gat), .B1(new_n861_), .B2(new_n544_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(KEYINPUT119), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n656_), .A2(new_n413_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n883_), .B1(new_n879_), .B2(new_n884_), .ZN(G1342gat));
  AOI21_X1  g684(.A(G134gat), .B1(new_n861_), .B2(new_n653_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(KEYINPUT120), .ZN(new_n887_));
  XNOR2_X1  g686(.A(KEYINPUT121), .B(G134gat), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n692_), .A2(new_n888_), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n887_), .B1(new_n879_), .B2(new_n889_), .ZN(G1343gat));
  AOI21_X1  g689(.A(new_n463_), .B1(new_n856_), .B2(new_n860_), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n891_), .A2(new_n337_), .A3(new_n482_), .A4(new_n440_), .ZN(new_n892_));
  NOR2_X1   g691(.A1(new_n892_), .A2(new_n655_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT122), .B(G141gat), .ZN(new_n894_));
  XNOR2_X1  g693(.A(new_n893_), .B(new_n894_), .ZN(G1344gat));
  NOR2_X1   g694(.A1(new_n892_), .A2(new_n700_), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n896_), .B(new_n358_), .ZN(G1345gat));
  NOR2_X1   g696(.A1(new_n892_), .A2(new_n656_), .ZN(new_n898_));
  XOR2_X1   g697(.A(KEYINPUT61), .B(G155gat), .Z(new_n899_));
  XNOR2_X1  g698(.A(new_n898_), .B(new_n899_), .ZN(G1346gat));
  OAI21_X1  g699(.A(G162gat), .B1(new_n892_), .B2(new_n692_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n653_), .A2(new_n349_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n901_), .B1(new_n892_), .B2(new_n902_), .ZN(G1347gat));
  NOR4_X1   g702(.A1(new_n489_), .A2(new_n337_), .A3(new_n482_), .A4(new_n440_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n864_), .A2(new_n519_), .A3(new_n904_), .ZN(new_n905_));
  AOI21_X1  g704(.A(KEYINPUT124), .B1(new_n905_), .B2(G169gat), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n907_));
  INV_X1    g706(.A(new_n905_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n906_), .A2(new_n907_), .B1(new_n908_), .B2(new_n295_), .ZN(new_n909_));
  OR2_X1    g708(.A1(new_n906_), .A2(new_n907_), .ZN(new_n910_));
  AND3_X1   g709(.A1(new_n905_), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n911_));
  OAI21_X1  g710(.A(new_n909_), .B1(new_n910_), .B2(new_n911_), .ZN(G1348gat));
  NAND2_X1  g711(.A1(new_n864_), .A2(new_n904_), .ZN(new_n913_));
  NOR2_X1   g712(.A1(new_n913_), .A2(new_n700_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(new_n914_), .B(new_n248_), .ZN(G1349gat));
  NOR2_X1   g714(.A1(new_n913_), .A2(new_n656_), .ZN(new_n916_));
  NOR2_X1   g715(.A1(new_n916_), .A2(G183gat), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n257_), .A2(new_n301_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n917_), .B1(new_n918_), .B2(new_n916_), .ZN(G1350gat));
  OAI21_X1  g718(.A(G190gat), .B1(new_n913_), .B2(new_n692_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n653_), .A2(new_n252_), .A3(new_n255_), .ZN(new_n921_));
  OAI21_X1  g720(.A(new_n920_), .B1(new_n913_), .B2(new_n921_), .ZN(G1351gat));
  NOR3_X1   g721(.A1(new_n337_), .A2(new_n405_), .A3(new_n440_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n848_), .A2(new_n852_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n924_), .A2(new_n708_), .ZN(new_n925_));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n926_));
  AOI21_X1  g725(.A(new_n692_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n925_), .A2(new_n926_), .B1(new_n846_), .B2(new_n927_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n853_), .A2(KEYINPUT57), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n544_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n930_));
  NAND2_X1  g729(.A1(new_n647_), .A2(new_n520_), .ZN(new_n931_));
  INV_X1    g730(.A(new_n857_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  NAND3_X1  g732(.A1(new_n647_), .A2(new_n520_), .A3(new_n857_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n933_), .A2(new_n934_), .ZN(new_n935_));
  OAI211_X1 g734(.A(new_n489_), .B(new_n923_), .C1(new_n930_), .C2(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(KEYINPUT125), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n891_), .A2(new_n938_), .A3(new_n923_), .ZN(new_n939_));
  AOI21_X1  g738(.A(new_n655_), .B1(new_n937_), .B2(new_n939_), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(new_n222_), .ZN(G1352gat));
  AOI21_X1  g740(.A(new_n700_), .B1(new_n937_), .B2(new_n939_), .ZN(new_n942_));
  XNOR2_X1  g741(.A(new_n942_), .B(new_n225_), .ZN(G1353gat));
  NAND2_X1  g742(.A1(new_n937_), .A2(new_n939_), .ZN(new_n944_));
  OR2_X1    g743(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n945_));
  NAND2_X1  g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  AND4_X1   g745(.A1(new_n544_), .A2(new_n944_), .A3(new_n945_), .A4(new_n946_), .ZN(new_n947_));
  AOI21_X1  g746(.A(new_n945_), .B1(new_n944_), .B2(new_n544_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n947_), .A2(new_n948_), .ZN(G1354gat));
  AOI211_X1 g748(.A(new_n210_), .B(new_n692_), .C1(new_n937_), .C2(new_n939_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n708_), .B1(new_n937_), .B2(new_n939_), .ZN(new_n951_));
  INV_X1    g750(.A(KEYINPUT126), .ZN(new_n952_));
  AOI21_X1  g751(.A(G218gat), .B1(new_n951_), .B2(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n936_), .A2(KEYINPUT125), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n938_), .B1(new_n891_), .B2(new_n923_), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n653_), .B1(new_n954_), .B2(new_n955_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n956_), .A2(KEYINPUT126), .ZN(new_n957_));
  AOI21_X1  g756(.A(new_n950_), .B1(new_n953_), .B2(new_n957_), .ZN(G1355gat));
endmodule


