//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n588_, new_n589_, new_n590_, new_n591_, new_n593_, new_n594_,
    new_n595_, new_n596_, new_n597_, new_n598_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n692_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n788_, new_n789_,
    new_n790_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n803_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n813_, new_n814_, new_n815_, new_n816_,
    new_n817_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n844_, new_n845_,
    new_n846_, new_n848_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n863_, new_n864_, new_n865_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_;
  XOR2_X1   g000(.A(G190gat), .B(G218gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(G134gat), .B(G162gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT36), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G29gat), .B(G36gat), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT71), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G43gat), .B(G50gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  XOR2_X1   g011(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n213_));
  XNOR2_X1  g012(.A(new_n212_), .B(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G99gat), .ZN(new_n216_));
  INV_X1    g015(.A(G106gat), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n216_), .A2(new_n217_), .A3(KEYINPUT66), .A4(KEYINPUT7), .ZN(new_n218_));
  NAND2_X1  g017(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n219_), .B1(G99gat), .B2(G106gat), .ZN(new_n220_));
  NOR2_X1   g019(.A1(KEYINPUT66), .A2(KEYINPUT7), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n218_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT6), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT64), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT6), .ZN(new_n226_));
  AND2_X1   g025(.A1(G99gat), .A2(G106gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n224_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(new_n227_), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n225_), .A2(KEYINPUT6), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n223_), .A2(KEYINPUT64), .ZN(new_n231_));
  OAI21_X1  g030(.A(new_n229_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n222_), .A2(new_n228_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT8), .ZN(new_n234_));
  INV_X1    g033(.A(G85gat), .ZN(new_n235_));
  INV_X1    g034(.A(G92gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(G85gat), .A2(G92gat), .ZN(new_n238_));
  AND3_X1   g037(.A1(new_n237_), .A2(KEYINPUT67), .A3(new_n238_), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n233_), .A2(new_n234_), .A3(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n234_), .B1(new_n233_), .B2(new_n239_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n232_), .A2(new_n228_), .ZN(new_n242_));
  OR2_X1    g041(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n243_));
  NAND2_X1  g042(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(new_n217_), .A3(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n237_), .A2(KEYINPUT9), .A3(new_n238_), .ZN(new_n246_));
  OR2_X1    g045(.A1(new_n238_), .A2(KEYINPUT9), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT65), .ZN(new_n249_));
  NOR3_X1   g048(.A1(new_n242_), .A2(new_n248_), .A3(new_n249_), .ZN(new_n250_));
  AND3_X1   g049(.A1(new_n245_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n251_));
  AND3_X1   g050(.A1(new_n224_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n227_), .B1(new_n224_), .B2(new_n226_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT65), .B1(new_n251_), .B2(new_n254_), .ZN(new_n255_));
  OAI22_X1  g054(.A1(new_n240_), .A2(new_n241_), .B1(new_n250_), .B2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(KEYINPUT69), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n251_), .A2(new_n254_), .A3(KEYINPUT65), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n249_), .B1(new_n242_), .B2(new_n248_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n261_));
  OAI211_X1 g060(.A(new_n260_), .B(new_n261_), .C1(new_n241_), .C2(new_n240_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(new_n262_), .ZN(new_n263_));
  OAI21_X1  g062(.A(KEYINPUT73), .B1(new_n215_), .B2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT73), .ZN(new_n265_));
  NAND4_X1  g064(.A1(new_n214_), .A2(new_n265_), .A3(new_n257_), .A4(new_n262_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n264_), .A2(new_n266_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n241_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n233_), .A2(new_n234_), .A3(new_n239_), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n268_), .A2(new_n269_), .B1(new_n259_), .B2(new_n258_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n212_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(G232gat), .A2(G233gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(KEYINPUT34), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(KEYINPUT35), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n274_), .B1(new_n267_), .B2(KEYINPUT74), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n273_), .A2(KEYINPUT35), .ZN(new_n276_));
  OAI211_X1 g075(.A(new_n267_), .B(new_n271_), .C1(new_n275_), .C2(new_n276_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n267_), .A2(new_n271_), .ZN(new_n278_));
  AND2_X1   g077(.A1(new_n267_), .A2(KEYINPUT74), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n278_), .B1(new_n279_), .B2(new_n274_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n208_), .B1(new_n277_), .B2(new_n280_), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n277_), .A2(new_n280_), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n206_), .B(KEYINPUT36), .Z(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n282_), .B(KEYINPUT37), .C1(new_n283_), .C2(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(KEYINPUT77), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n285_), .B1(new_n283_), .B2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n277_), .A2(new_n280_), .A3(KEYINPUT77), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n281_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n286_), .B1(new_n290_), .B2(KEYINPUT37), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G57gat), .B(G64gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(KEYINPUT11), .ZN(new_n293_));
  XOR2_X1   g092(.A(G71gat), .B(G78gat), .Z(new_n294_));
  OR2_X1    g093(.A1(new_n293_), .A2(new_n294_), .ZN(new_n295_));
  NOR2_X1   g094(.A1(new_n292_), .A2(KEYINPUT11), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n293_), .A2(new_n294_), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n295_), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G231gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT78), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G15gat), .B(G22gat), .ZN(new_n302_));
  INV_X1    g101(.A(G1gat), .ZN(new_n303_));
  INV_X1    g102(.A(G8gat), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT14), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n302_), .A2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G1gat), .B(G8gat), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n306_), .B(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n301_), .B(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT17), .ZN(new_n310_));
  XOR2_X1   g109(.A(G127gat), .B(G155gat), .Z(new_n311_));
  XNOR2_X1  g110(.A(new_n311_), .B(KEYINPUT16), .ZN(new_n312_));
  XNOR2_X1  g111(.A(G183gat), .B(G211gat), .ZN(new_n313_));
  XNOR2_X1  g112(.A(new_n312_), .B(new_n313_), .ZN(new_n314_));
  OR3_X1    g113(.A1(new_n309_), .A2(new_n310_), .A3(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n314_), .B(KEYINPUT17), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n309_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(new_n291_), .A2(new_n318_), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n319_), .B(KEYINPUT79), .Z(new_n320_));
  INV_X1    g119(.A(KEYINPUT82), .ZN(new_n321_));
  INV_X1    g120(.A(G169gat), .ZN(new_n322_));
  INV_X1    g121(.A(G176gat), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n322_), .A3(new_n323_), .ZN(new_n324_));
  OAI21_X1  g123(.A(KEYINPUT82), .B1(G169gat), .B2(G176gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G169gat), .A2(G176gat), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT24), .ZN(new_n328_));
  OR3_X1    g127(.A1(new_n326_), .A2(KEYINPUT83), .A3(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(KEYINPUT83), .B1(new_n326_), .B2(new_n328_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT24), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(KEYINPUT25), .B(G183gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT26), .B(G190gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n334_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G183gat), .A2(G190gat), .ZN(new_n337_));
  XNOR2_X1  g136(.A(new_n337_), .B(KEYINPUT23), .ZN(new_n338_));
  AND2_X1   g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n331_), .A2(new_n333_), .A3(new_n339_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n338_), .B1(G183gat), .B2(G190gat), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT84), .B(G176gat), .ZN(new_n342_));
  XNOR2_X1  g141(.A(KEYINPUT22), .B(G169gat), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n341_), .A2(new_n327_), .A3(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n340_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G71gat), .B(G99gat), .ZN(new_n347_));
  INV_X1    g146(.A(G43gat), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n346_), .B(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G127gat), .B(G134gat), .Z(new_n351_));
  XOR2_X1   g150(.A(G113gat), .B(G120gat), .Z(new_n352_));
  XOR2_X1   g151(.A(new_n351_), .B(new_n352_), .Z(new_n353_));
  INV_X1    g152(.A(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n350_), .B(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(G227gat), .A2(G233gat), .ZN(new_n356_));
  XOR2_X1   g155(.A(new_n356_), .B(G15gat), .Z(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(KEYINPUT30), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(KEYINPUT31), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n355_), .A2(new_n359_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n360_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT92), .ZN(new_n364_));
  INV_X1    g163(.A(G197gat), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n365_), .A2(G204gat), .ZN(new_n366_));
  INV_X1    g165(.A(G204gat), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n367_), .A2(G197gat), .ZN(new_n368_));
  AND2_X1   g167(.A1(new_n366_), .A2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(KEYINPUT86), .ZN(new_n370_));
  OAI211_X1 g169(.A(new_n370_), .B(KEYINPUT21), .C1(KEYINPUT86), .C2(new_n366_), .ZN(new_n371_));
  XOR2_X1   g170(.A(G211gat), .B(G218gat), .Z(new_n372_));
  INV_X1    g171(.A(KEYINPUT21), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n372_), .B1(new_n373_), .B2(new_n369_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n371_), .A2(new_n374_), .ZN(new_n375_));
  OR2_X1    g174(.A1(new_n369_), .A2(KEYINPUT87), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n369_), .A2(KEYINPUT87), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n376_), .A2(new_n377_), .A3(KEYINPUT21), .A4(new_n372_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n375_), .A2(new_n378_), .ZN(new_n379_));
  OAI21_X1  g178(.A(KEYINPUT20), .B1(new_n346_), .B2(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT90), .ZN(new_n381_));
  AND3_X1   g180(.A1(new_n344_), .A2(new_n381_), .A3(new_n327_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n381_), .B1(new_n344_), .B2(new_n327_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n341_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT91), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n328_), .A2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n327_), .A2(KEYINPUT88), .A3(KEYINPUT24), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n388_), .A2(new_n324_), .A3(new_n325_), .A4(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT89), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n390_), .A2(new_n391_), .A3(new_n336_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n391_), .B1(new_n390_), .B2(new_n336_), .ZN(new_n393_));
  OAI211_X1 g192(.A(new_n338_), .B(new_n333_), .C1(new_n392_), .C2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(KEYINPUT91), .B(new_n341_), .C1(new_n382_), .C2(new_n383_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n386_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n380_), .B1(new_n379_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT19), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n364_), .B1(new_n397_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n396_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n379_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(KEYINPUT92), .B(new_n399_), .C1(new_n404_), .C2(new_n380_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n401_), .A2(new_n405_), .ZN(new_n406_));
  XOR2_X1   g205(.A(G8gat), .B(G36gat), .Z(new_n407_));
  XNOR2_X1  g206(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n407_), .B(new_n408_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G64gat), .B(G92gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT20), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n413_), .B1(new_n346_), .B2(new_n379_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n414_), .B(new_n400_), .C1(new_n396_), .C2(new_n379_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n406_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n403_), .A2(new_n394_), .A3(new_n384_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n400_), .B1(new_n414_), .B2(new_n417_), .ZN(new_n418_));
  AOI22_X1  g217(.A1(new_n397_), .A2(new_n400_), .B1(new_n418_), .B2(KEYINPUT96), .ZN(new_n419_));
  OR2_X1    g218(.A1(new_n418_), .A2(KEYINPUT96), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n412_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT97), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n416_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n419_), .A2(new_n420_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n424_), .A2(new_n422_), .A3(new_n411_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT27), .ZN(new_n426_));
  OAI21_X1  g225(.A(KEYINPUT98), .B1(new_n423_), .B2(new_n426_), .ZN(new_n427_));
  OR2_X1    g226(.A1(new_n421_), .A2(new_n422_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT27), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n429_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT98), .ZN(new_n431_));
  NAND4_X1  g230(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .A4(new_n416_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n427_), .A2(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n412_), .B1(new_n406_), .B2(new_n415_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n415_), .ZN(new_n435_));
  AOI211_X1 g234(.A(new_n411_), .B(new_n435_), .C1(new_n401_), .C2(new_n405_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n429_), .B1(new_n434_), .B2(new_n436_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT99), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT99), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n439_), .B(new_n429_), .C1(new_n434_), .C2(new_n436_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n438_), .A2(new_n440_), .ZN(new_n441_));
  XOR2_X1   g240(.A(G155gat), .B(G162gat), .Z(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT85), .ZN(new_n443_));
  OR2_X1    g242(.A1(G141gat), .A2(G148gat), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n444_), .A2(KEYINPUT3), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G141gat), .A2(G148gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT2), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n444_), .A2(KEYINPUT3), .ZN(new_n450_));
  NAND4_X1  g249(.A1(new_n445_), .A2(new_n448_), .A3(new_n449_), .A4(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n443_), .A2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(G155gat), .ZN(new_n453_));
  INV_X1    g252(.A(G162gat), .ZN(new_n454_));
  OAI21_X1  g253(.A(KEYINPUT1), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n455_), .B1(G155gat), .B2(G162gat), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n453_), .A2(new_n454_), .A3(KEYINPUT1), .ZN(new_n457_));
  OAI211_X1 g256(.A(new_n446_), .B(new_n444_), .C1(new_n456_), .C2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n452_), .A2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n459_), .A2(KEYINPUT29), .ZN(new_n460_));
  XOR2_X1   g259(.A(new_n460_), .B(KEYINPUT28), .Z(new_n461_));
  AOI21_X1  g260(.A(new_n403_), .B1(new_n459_), .B2(KEYINPUT29), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n461_), .B(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G228gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(G78gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n464_), .B(new_n465_), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(new_n217_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G22gat), .B(G50gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(new_n463_), .B(new_n469_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n459_), .A2(new_n353_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n354_), .A2(new_n452_), .A3(new_n458_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n471_), .A2(new_n472_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(G225gat), .A2(G233gat), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n473_), .A2(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n471_), .A2(KEYINPUT4), .A3(new_n472_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT4), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n459_), .A2(new_n478_), .A3(new_n353_), .ZN(new_n479_));
  AOI21_X1  g278(.A(new_n474_), .B1(new_n477_), .B2(new_n479_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n476_), .A2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(G1gat), .B(G29gat), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n482_), .B(G85gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT0), .B(G57gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(new_n483_), .B(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  XNOR2_X1  g285(.A(new_n481_), .B(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n470_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n433_), .A2(new_n441_), .A3(new_n488_), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n406_), .A2(new_n415_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(new_n411_), .ZN(new_n491_));
  OAI21_X1  g290(.A(new_n486_), .B1(new_n476_), .B2(new_n480_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT33), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT33), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n494_), .B(new_n486_), .C1(new_n476_), .C2(new_n480_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n486_), .B1(new_n473_), .B2(new_n475_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n477_), .A2(new_n474_), .A3(new_n479_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT94), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT94), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n496_), .A2(new_n497_), .A3(new_n500_), .ZN(new_n501_));
  AOI22_X1  g300(.A1(new_n493_), .A2(new_n495_), .B1(new_n499_), .B2(new_n501_), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n491_), .A2(new_n416_), .A3(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT95), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND4_X1  g304(.A1(new_n491_), .A2(KEYINPUT95), .A3(new_n416_), .A4(new_n502_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n412_), .A2(KEYINPUT32), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n424_), .A2(new_n507_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n487_), .B(new_n508_), .C1(new_n490_), .C2(new_n507_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n505_), .A2(new_n506_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(new_n470_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n363_), .B1(new_n489_), .B2(new_n511_), .ZN(new_n512_));
  NOR2_X1   g311(.A1(new_n362_), .A2(new_n487_), .ZN(new_n513_));
  AND4_X1   g312(.A1(new_n433_), .A2(new_n441_), .A3(new_n470_), .A4(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n270_), .A2(new_n298_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT68), .ZN(new_n517_));
  AND2_X1   g316(.A1(G230gat), .A2(G233gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n270_), .A2(new_n298_), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT68), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n519_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n517_), .B(new_n518_), .C1(new_n521_), .C2(new_n516_), .ZN(new_n522_));
  OAI211_X1 g321(.A(new_n295_), .B(KEYINPUT12), .C1(new_n296_), .C2(new_n297_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n257_), .A2(new_n262_), .A3(new_n524_), .ZN(new_n525_));
  XOR2_X1   g324(.A(KEYINPUT70), .B(KEYINPUT12), .Z(new_n526_));
  OAI21_X1  g325(.A(new_n526_), .B1(new_n270_), .B2(new_n298_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n518_), .B1(new_n270_), .B2(new_n298_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n525_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n522_), .A2(new_n529_), .ZN(new_n530_));
  XOR2_X1   g329(.A(G120gat), .B(G148gat), .Z(new_n531_));
  XNOR2_X1  g330(.A(new_n531_), .B(KEYINPUT5), .ZN(new_n532_));
  XNOR2_X1  g331(.A(G176gat), .B(G204gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  OR2_X1    g333(.A1(new_n530_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n530_), .A2(new_n534_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT13), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n535_), .A2(KEYINPUT13), .A3(new_n536_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n308_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n212_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G229gat), .A2(G233gat), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n543_), .A2(new_n545_), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n214_), .A2(new_n308_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n212_), .A2(new_n542_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n548_), .A2(new_n544_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n546_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(G113gat), .B(G141gat), .Z(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT80), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G169gat), .B(G197gat), .ZN(new_n553_));
  XOR2_X1   g352(.A(new_n552_), .B(new_n553_), .Z(new_n554_));
  XNOR2_X1  g353(.A(new_n550_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT81), .ZN(new_n556_));
  NOR3_X1   g355(.A1(new_n515_), .A2(new_n541_), .A3(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n320_), .A2(new_n557_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n487_), .A2(new_n303_), .ZN(new_n559_));
  INV_X1    g358(.A(KEYINPUT102), .ZN(new_n560_));
  XNOR2_X1  g359(.A(KEYINPUT100), .B(KEYINPUT38), .ZN(new_n561_));
  OAI22_X1  g360(.A1(new_n558_), .A2(new_n559_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n561_), .A2(new_n560_), .ZN(new_n563_));
  OR2_X1    g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n562_), .A2(new_n563_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT101), .ZN(new_n566_));
  OR2_X1    g365(.A1(new_n512_), .A2(new_n514_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n290_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n566_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n566_), .B(new_n568_), .C1(new_n512_), .C2(new_n514_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n569_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n555_), .ZN(new_n573_));
  NOR3_X1   g372(.A1(new_n541_), .A2(new_n318_), .A3(new_n573_), .ZN(new_n574_));
  AND3_X1   g373(.A1(new_n572_), .A2(new_n487_), .A3(new_n574_), .ZN(new_n575_));
  OAI211_X1 g374(.A(new_n564_), .B(new_n565_), .C1(new_n303_), .C2(new_n575_), .ZN(G1324gat));
  NAND2_X1  g375(.A1(new_n433_), .A2(new_n441_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n320_), .A2(new_n304_), .A3(new_n577_), .A4(new_n557_), .ZN(new_n578_));
  OAI211_X1 g377(.A(new_n577_), .B(new_n574_), .C1(new_n569_), .C2(new_n571_), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT39), .ZN(new_n580_));
  AND3_X1   g379(.A1(new_n579_), .A2(new_n580_), .A3(G8gat), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n580_), .B1(new_n579_), .B2(G8gat), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n578_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT40), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  OAI211_X1 g384(.A(new_n578_), .B(KEYINPUT40), .C1(new_n581_), .C2(new_n582_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(G1325gat));
  OR3_X1    g386(.A1(new_n558_), .A2(G15gat), .A3(new_n362_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n572_), .A2(new_n363_), .A3(new_n574_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n589_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n590_));
  AOI21_X1  g389(.A(KEYINPUT41), .B1(new_n589_), .B2(G15gat), .ZN(new_n591_));
  OAI21_X1  g390(.A(new_n588_), .B1(new_n590_), .B2(new_n591_), .ZN(G1326gat));
  OR3_X1    g391(.A1(new_n558_), .A2(G22gat), .A3(new_n470_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n470_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n572_), .A2(new_n594_), .A3(new_n574_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT42), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n595_), .A2(new_n596_), .A3(G22gat), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n595_), .B2(G22gat), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n593_), .B1(new_n597_), .B2(new_n598_), .ZN(G1327gat));
  NAND2_X1  g398(.A1(new_n290_), .A2(new_n318_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n557_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n487_), .ZN(new_n603_));
  OR3_X1    g402(.A1(new_n602_), .A2(G29gat), .A3(new_n603_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n291_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT43), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT43), .ZN(new_n607_));
  OAI211_X1 g406(.A(new_n607_), .B(new_n291_), .C1(new_n512_), .C2(new_n514_), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n606_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n541_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n610_), .A2(new_n318_), .A3(new_n555_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT103), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n609_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT44), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n614_), .A2(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n609_), .A2(KEYINPUT44), .A3(new_n613_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n616_), .A2(new_n487_), .A3(new_n617_), .ZN(new_n618_));
  AND3_X1   g417(.A1(new_n618_), .A2(KEYINPUT104), .A3(G29gat), .ZN(new_n619_));
  AOI21_X1  g418(.A(KEYINPUT104), .B1(new_n618_), .B2(G29gat), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n604_), .B1(new_n619_), .B2(new_n620_), .ZN(G1328gat));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n622_), .A2(KEYINPUT46), .ZN(new_n623_));
  INV_X1    g422(.A(G36gat), .ZN(new_n624_));
  AOI21_X1  g423(.A(KEYINPUT44), .B1(new_n609_), .B2(new_n613_), .ZN(new_n625_));
  AOI211_X1 g424(.A(new_n615_), .B(new_n612_), .C1(new_n606_), .C2(new_n608_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n624_), .B1(new_n627_), .B2(new_n577_), .ZN(new_n628_));
  INV_X1    g427(.A(new_n602_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT45), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n577_), .A2(new_n624_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n629_), .A2(new_n630_), .A3(new_n632_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT45), .B1(new_n602_), .B2(new_n631_), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n623_), .B1(new_n628_), .B2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(new_n623_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(new_n634_), .ZN(new_n638_));
  AND3_X1   g437(.A1(new_n616_), .A2(new_n577_), .A3(new_n617_), .ZN(new_n639_));
  OAI211_X1 g438(.A(new_n637_), .B(new_n638_), .C1(new_n639_), .C2(new_n624_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(G1329gat));
  NOR4_X1   g440(.A1(new_n625_), .A2(new_n626_), .A3(new_n348_), .A4(new_n362_), .ZN(new_n642_));
  AOI21_X1  g441(.A(G43gat), .B1(new_n629_), .B2(new_n363_), .ZN(new_n643_));
  OAI21_X1  g442(.A(KEYINPUT47), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n627_), .A2(G43gat), .A3(new_n363_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT47), .ZN(new_n646_));
  INV_X1    g445(.A(new_n643_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n645_), .A2(new_n646_), .A3(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n644_), .A2(new_n648_), .ZN(G1330gat));
  OR3_X1    g448(.A1(new_n602_), .A2(G50gat), .A3(new_n470_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n627_), .A2(KEYINPUT106), .A3(new_n594_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n651_), .A2(G50gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(KEYINPUT106), .B1(new_n627_), .B2(new_n594_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n650_), .B1(new_n652_), .B2(new_n653_), .ZN(G1331gat));
  NOR3_X1   g453(.A1(new_n515_), .A2(new_n610_), .A3(new_n555_), .ZN(new_n655_));
  AND2_X1   g454(.A1(new_n320_), .A2(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(G57gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n656_), .A2(new_n657_), .A3(new_n487_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n318_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n556_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n660_), .A2(new_n610_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n572_), .A2(new_n487_), .A3(new_n661_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n658_), .B1(new_n662_), .B2(new_n657_), .ZN(G1332gat));
  INV_X1    g462(.A(G64gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n656_), .A2(new_n664_), .A3(new_n577_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n572_), .A2(new_n577_), .A3(new_n661_), .ZN(new_n666_));
  XNOR2_X1  g465(.A(KEYINPUT107), .B(KEYINPUT48), .ZN(new_n667_));
  AND3_X1   g466(.A1(new_n666_), .A2(G64gat), .A3(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n667_), .B1(new_n666_), .B2(G64gat), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(G1333gat));
  INV_X1    g469(.A(G71gat), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n656_), .A2(new_n671_), .A3(new_n363_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n572_), .A2(new_n363_), .A3(new_n661_), .ZN(new_n673_));
  INV_X1    g472(.A(KEYINPUT49), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n673_), .A2(new_n674_), .A3(G71gat), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n674_), .B1(new_n673_), .B2(G71gat), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n672_), .B1(new_n675_), .B2(new_n676_), .ZN(G1334gat));
  NAND3_X1  g476(.A1(new_n656_), .A2(new_n465_), .A3(new_n594_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n572_), .A2(new_n594_), .A3(new_n661_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT50), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n679_), .A2(new_n680_), .A3(G78gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n680_), .B1(new_n679_), .B2(G78gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n678_), .B1(new_n681_), .B2(new_n682_), .ZN(G1335gat));
  NAND2_X1  g482(.A1(new_n655_), .A2(new_n601_), .ZN(new_n684_));
  INV_X1    g483(.A(new_n684_), .ZN(new_n685_));
  NAND3_X1  g484(.A1(new_n685_), .A2(new_n235_), .A3(new_n487_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n610_), .A2(new_n555_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n318_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n688_), .B1(new_n606_), .B2(new_n608_), .ZN(new_n689_));
  AND2_X1   g488(.A1(new_n689_), .A2(new_n487_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n686_), .B1(new_n690_), .B2(new_n235_), .ZN(G1336gat));
  AOI21_X1  g490(.A(G92gat), .B1(new_n685_), .B2(new_n577_), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n577_), .A2(G92gat), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT108), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n692_), .B1(new_n689_), .B2(new_n694_), .ZN(G1337gat));
  INV_X1    g494(.A(KEYINPUT109), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(KEYINPUT51), .ZN(new_n697_));
  AND3_X1   g496(.A1(new_n363_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n697_), .B1(new_n684_), .B2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n689_), .A2(new_n363_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(G99gat), .B2(new_n701_), .ZN(new_n702_));
  NOR2_X1   g501(.A1(new_n696_), .A2(KEYINPUT51), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n702_), .B(new_n703_), .ZN(G1338gat));
  NAND3_X1  g503(.A1(new_n685_), .A2(new_n217_), .A3(new_n594_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n689_), .A2(new_n594_), .ZN(new_n706_));
  NOR2_X1   g505(.A1(KEYINPUT110), .A2(KEYINPUT52), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n217_), .B1(KEYINPUT110), .B2(KEYINPUT52), .ZN(new_n708_));
  AND3_X1   g507(.A1(new_n706_), .A2(new_n707_), .A3(new_n708_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n707_), .B1(new_n706_), .B2(new_n708_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n705_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n711_), .A2(KEYINPUT53), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT53), .ZN(new_n713_));
  OAI211_X1 g512(.A(new_n713_), .B(new_n705_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n712_), .A2(new_n714_), .ZN(G1339gat));
  INV_X1    g514(.A(new_n556_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n660_), .A2(new_n541_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n717_), .B(new_n286_), .C1(new_n290_), .C2(KEYINPUT37), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT54), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n718_), .B(new_n719_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n550_), .A2(new_n554_), .ZN(new_n721_));
  OAI211_X1 g520(.A(new_n548_), .B(new_n545_), .C1(new_n215_), .C2(new_n542_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n554_), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n721_), .B1(new_n722_), .B2(new_n724_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n537_), .A2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n525_), .A2(new_n527_), .A3(new_n519_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n529_), .A2(KEYINPUT55), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT55), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n525_), .A2(new_n730_), .A3(new_n527_), .A4(new_n528_), .ZN(new_n731_));
  AOI221_X4 g530(.A(new_n727_), .B1(new_n728_), .B2(new_n518_), .C1(new_n729_), .C2(new_n731_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n729_), .A2(new_n731_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n728_), .A2(new_n518_), .ZN(new_n734_));
  AOI21_X1  g533(.A(KEYINPUT111), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  OAI211_X1 g534(.A(KEYINPUT56), .B(new_n534_), .C1(new_n732_), .C2(new_n735_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n534_), .B1(new_n732_), .B2(new_n735_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT56), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n737_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n738_), .B1(new_n737_), .B2(new_n739_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n736_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n555_), .A2(new_n535_), .ZN(new_n743_));
  INV_X1    g542(.A(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n726_), .B1(new_n742_), .B2(new_n744_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT57), .ZN(new_n746_));
  OR3_X1    g545(.A1(new_n745_), .A2(new_n746_), .A3(new_n290_), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(new_n290_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n725_), .A2(new_n535_), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT113), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT114), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n737_), .B2(new_n739_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n736_), .ZN(new_n753_));
  NOR2_X1   g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n737_), .A2(new_n751_), .A3(new_n739_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n750_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT58), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  OAI211_X1 g557(.A(KEYINPUT58), .B(new_n750_), .C1(new_n754_), .C2(new_n755_), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n758_), .A2(new_n291_), .A3(new_n759_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n747_), .A2(new_n748_), .A3(new_n760_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n720_), .B1(new_n761_), .B2(new_n318_), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n577_), .A2(new_n594_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n603_), .A2(new_n362_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT59), .B1(new_n762_), .B2(new_n765_), .ZN(new_n766_));
  NOR3_X1   g565(.A1(new_n745_), .A2(new_n746_), .A3(new_n290_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n760_), .A2(new_n748_), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(KEYINPUT115), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n760_), .A2(new_n748_), .A3(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n659_), .B1(new_n769_), .B2(new_n771_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n772_), .A2(new_n720_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n765_), .A2(KEYINPUT59), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n716_), .B(new_n766_), .C1(new_n773_), .C2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(G113gat), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n762_), .A2(new_n765_), .ZN(new_n778_));
  INV_X1    g577(.A(new_n778_), .ZN(new_n779_));
  OR3_X1    g578(.A1(new_n779_), .A2(G113gat), .A3(new_n573_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n777_), .A2(new_n780_), .ZN(G1340gat));
  OAI211_X1 g580(.A(new_n541_), .B(new_n766_), .C1(new_n773_), .C2(new_n775_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(G120gat), .ZN(new_n783_));
  INV_X1    g582(.A(G120gat), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n784_), .B1(new_n610_), .B2(KEYINPUT60), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n778_), .B(new_n785_), .C1(KEYINPUT60), .C2(new_n784_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n783_), .A2(new_n786_), .ZN(G1341gat));
  OAI211_X1 g586(.A(new_n659_), .B(new_n766_), .C1(new_n773_), .C2(new_n775_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(G127gat), .ZN(new_n789_));
  OR3_X1    g588(.A1(new_n779_), .A2(G127gat), .A3(new_n318_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(G1342gat));
  AOI21_X1  g590(.A(G134gat), .B1(new_n778_), .B2(new_n290_), .ZN(new_n792_));
  OR2_X1    g591(.A1(new_n772_), .A2(new_n720_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n793_), .A2(new_n774_), .B1(new_n779_), .B2(KEYINPUT59), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n291_), .A2(G134gat), .ZN(new_n795_));
  XOR2_X1   g594(.A(new_n795_), .B(KEYINPUT116), .Z(new_n796_));
  AOI21_X1  g595(.A(new_n792_), .B1(new_n794_), .B2(new_n796_), .ZN(G1343gat));
  NOR2_X1   g596(.A1(new_n470_), .A2(new_n363_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n433_), .A2(new_n441_), .A3(new_n487_), .A4(new_n798_), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n799_), .B(KEYINPUT117), .ZN(new_n800_));
  INV_X1    g599(.A(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n762_), .A2(new_n801_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n555_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(G141gat), .ZN(G1344gat));
  XNOR2_X1  g603(.A(KEYINPUT118), .B(G148gat), .ZN(new_n805_));
  INV_X1    g604(.A(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n318_), .B1(new_n768_), .B2(new_n767_), .ZN(new_n807_));
  INV_X1    g606(.A(new_n720_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(new_n800_), .ZN(new_n810_));
  NOR3_X1   g609(.A1(new_n810_), .A2(KEYINPUT119), .A3(new_n610_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n812_), .B1(new_n802_), .B2(new_n541_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n806_), .B1(new_n811_), .B2(new_n813_), .ZN(new_n814_));
  OAI21_X1  g613(.A(KEYINPUT119), .B1(new_n810_), .B2(new_n610_), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n802_), .A2(new_n812_), .A3(new_n541_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n816_), .A3(new_n805_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n817_), .ZN(G1345gat));
  NAND2_X1  g617(.A1(new_n802_), .A2(new_n659_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(KEYINPUT61), .B(G155gat), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(G1346gat));
  AOI21_X1  g620(.A(G162gat), .B1(new_n802_), .B2(new_n290_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n291_), .A2(G162gat), .ZN(new_n823_));
  XOR2_X1   g622(.A(new_n823_), .B(KEYINPUT120), .Z(new_n824_));
  AOI21_X1  g623(.A(new_n822_), .B1(new_n802_), .B2(new_n824_), .ZN(G1347gat));
  NAND2_X1  g624(.A1(new_n577_), .A2(new_n513_), .ZN(new_n826_));
  NOR2_X1   g625(.A1(new_n826_), .A2(new_n594_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n555_), .B(new_n827_), .C1(new_n772_), .C2(new_n720_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n322_), .B1(new_n829_), .B2(KEYINPUT62), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n828_), .A2(new_n830_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n829_), .A2(KEYINPUT62), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n831_), .A2(new_n832_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n828_), .B(new_n830_), .C1(new_n829_), .C2(KEYINPUT62), .ZN(new_n834_));
  NAND4_X1  g633(.A1(new_n793_), .A2(new_n343_), .A3(new_n555_), .A4(new_n827_), .ZN(new_n835_));
  NAND3_X1  g634(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .ZN(G1348gat));
  NOR2_X1   g635(.A1(new_n762_), .A2(new_n594_), .ZN(new_n837_));
  NOR3_X1   g636(.A1(new_n826_), .A2(new_n323_), .A3(new_n610_), .ZN(new_n838_));
  AND2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n827_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(new_n773_), .A2(new_n840_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(new_n541_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n839_), .B1(new_n842_), .B2(new_n342_), .ZN(G1349gat));
  NOR2_X1   g642(.A1(new_n826_), .A2(new_n318_), .ZN(new_n844_));
  AOI21_X1  g643(.A(G183gat), .B1(new_n837_), .B2(new_n844_), .ZN(new_n845_));
  NOR2_X1   g644(.A1(new_n318_), .A2(new_n334_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n845_), .B1(new_n841_), .B2(new_n846_), .ZN(G1350gat));
  NAND3_X1  g646(.A1(new_n793_), .A2(new_n291_), .A3(new_n827_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n848_), .A2(G190gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n841_), .A2(new_n290_), .A3(new_n335_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n849_), .A2(new_n850_), .ZN(G1351gat));
  XNOR2_X1  g650(.A(KEYINPUT123), .B(G197gat), .ZN(new_n852_));
  INV_X1    g651(.A(KEYINPUT122), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n577_), .A2(new_n603_), .A3(new_n798_), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n762_), .B2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n854_), .ZN(new_n856_));
  NAND3_X1  g655(.A1(new_n809_), .A2(KEYINPUT122), .A3(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n852_), .B1(new_n858_), .B2(new_n555_), .ZN(new_n859_));
  AND2_X1   g658(.A1(new_n365_), .A2(KEYINPUT123), .ZN(new_n860_));
  AOI211_X1 g659(.A(new_n573_), .B(new_n860_), .C1(new_n855_), .C2(new_n857_), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n859_), .A2(new_n861_), .ZN(G1352gat));
  OAI211_X1 g661(.A(new_n858_), .B(new_n541_), .C1(KEYINPUT124), .C2(new_n367_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n610_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT124), .B(G204gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n863_), .B1(new_n864_), .B2(new_n865_), .ZN(G1353gat));
  AOI21_X1  g665(.A(new_n318_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n867_));
  XNOR2_X1  g666(.A(new_n867_), .B(KEYINPUT125), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n858_), .A2(new_n868_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT126), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n869_), .A2(new_n872_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n858_), .A2(new_n871_), .A3(new_n868_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n873_), .A2(new_n874_), .ZN(G1354gat));
  NAND2_X1  g674(.A1(new_n858_), .A2(new_n290_), .ZN(new_n876_));
  INV_X1    g675(.A(G218gat), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n291_), .A2(G218gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n878_), .B(KEYINPUT127), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n876_), .A2(new_n877_), .B1(new_n858_), .B2(new_n879_), .ZN(G1355gat));
endmodule


