//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n771_, new_n772_,
    new_n774_, new_n775_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n814_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n822_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n907_, new_n909_, new_n910_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n960_, new_n961_,
    new_n962_, new_n963_, new_n964_, new_n965_, new_n966_, new_n967_,
    new_n968_, new_n969_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_;
  NAND2_X1  g000(.A1(G99gat), .A2(G106gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT6), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(G85gat), .B(G92gat), .Z(new_n205_));
  AOI21_X1  g004(.A(new_n204_), .B1(KEYINPUT9), .B2(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT10), .B(G99gat), .Z(new_n207_));
  INV_X1    g006(.A(G106gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT64), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XOR2_X1   g010(.A(KEYINPUT65), .B(G85gat), .Z(new_n212_));
  INV_X1    g011(.A(KEYINPUT9), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n212_), .A2(new_n213_), .A3(G92gat), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n207_), .A2(KEYINPUT64), .A3(new_n208_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n206_), .A2(new_n211_), .A3(new_n214_), .A4(new_n215_), .ZN(new_n216_));
  NOR2_X1   g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT7), .ZN(new_n218_));
  XNOR2_X1  g017(.A(new_n217_), .B(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n205_), .B1(new_n219_), .B2(new_n204_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(KEYINPUT8), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT8), .ZN(new_n222_));
  XNOR2_X1  g021(.A(new_n217_), .B(KEYINPUT7), .ZN(new_n223_));
  XNOR2_X1  g022(.A(new_n202_), .B(KEYINPUT6), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  AOI21_X1  g024(.A(new_n222_), .B1(new_n225_), .B2(new_n205_), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n216_), .B1(new_n221_), .B2(new_n226_), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT66), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  OAI211_X1 g028(.A(new_n216_), .B(KEYINPUT66), .C1(new_n221_), .C2(new_n226_), .ZN(new_n230_));
  XNOR2_X1  g029(.A(G57gat), .B(G64gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT11), .ZN(new_n232_));
  XOR2_X1   g031(.A(G71gat), .B(G78gat), .Z(new_n233_));
  OR2_X1    g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n231_), .A2(KEYINPUT11), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n232_), .A2(new_n233_), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n234_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n229_), .A2(new_n230_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n237_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n227_), .A2(new_n239_), .A3(KEYINPUT12), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n237_), .B1(new_n229_), .B2(new_n230_), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n238_), .B(new_n240_), .C1(new_n241_), .C2(KEYINPUT12), .ZN(new_n242_));
  NAND2_X1  g041(.A1(G230gat), .A2(G233gat), .ZN(new_n243_));
  INV_X1    g042(.A(new_n243_), .ZN(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT67), .B1(new_n242_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n220_), .B(KEYINPUT8), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT66), .B1(new_n246_), .B2(new_n216_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n230_), .ZN(new_n248_));
  OAI21_X1  g047(.A(new_n239_), .B1(new_n247_), .B2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(new_n238_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n250_), .A2(new_n244_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n238_), .A2(new_n240_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT12), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n249_), .A2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT67), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n252_), .A2(new_n254_), .A3(new_n255_), .A4(new_n243_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n245_), .A2(new_n251_), .A3(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G120gat), .B(G148gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n258_), .B(KEYINPUT5), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G176gat), .B(G204gat), .ZN(new_n260_));
  XOR2_X1   g059(.A(new_n259_), .B(new_n260_), .Z(new_n261_));
  NAND2_X1  g060(.A1(new_n257_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n261_), .ZN(new_n263_));
  NAND4_X1  g062(.A1(new_n245_), .A2(new_n256_), .A3(new_n251_), .A4(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n262_), .A2(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT13), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n262_), .A2(KEYINPUT13), .A3(new_n264_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  XOR2_X1   g069(.A(G127gat), .B(G155gat), .Z(new_n271_));
  XNOR2_X1  g070(.A(new_n271_), .B(KEYINPUT16), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G183gat), .B(G211gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G1gat), .B(G8gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n276_), .B(KEYINPUT70), .ZN(new_n277_));
  INV_X1    g076(.A(G15gat), .ZN(new_n278_));
  INV_X1    g077(.A(G22gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G15gat), .A2(G22gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(G1gat), .A2(G8gat), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n280_), .A2(new_n281_), .B1(KEYINPUT14), .B2(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n277_), .B(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  OR2_X1    g084(.A1(new_n236_), .A2(new_n235_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G231gat), .A2(G233gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(new_n287_), .A3(new_n234_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n287_), .B1(new_n286_), .B2(new_n234_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n285_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n237_), .A2(G231gat), .A3(G233gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n292_), .A2(new_n284_), .A3(new_n288_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT71), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n275_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT17), .B1(new_n294_), .B2(new_n275_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  OAI211_X1 g097(.A(KEYINPUT17), .B(new_n275_), .C1(new_n294_), .C2(new_n295_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G113gat), .B(G141gat), .Z(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(KEYINPUT74), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G169gat), .B(G197gat), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n302_), .B(new_n303_), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n304_), .A2(KEYINPUT73), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G29gat), .B(G36gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT68), .ZN(new_n307_));
  XNOR2_X1  g106(.A(G43gat), .B(G50gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XOR2_X1   g108(.A(new_n309_), .B(new_n284_), .Z(new_n310_));
  NAND2_X1  g109(.A1(G229gat), .A2(G233gat), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n310_), .A2(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n285_), .A2(new_n309_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(new_n311_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n309_), .B(KEYINPUT15), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n316_), .B1(new_n317_), .B2(new_n284_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n305_), .B1(new_n314_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n284_), .ZN(new_n320_));
  NAND3_X1  g119(.A1(new_n320_), .A2(new_n315_), .A3(new_n311_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n305_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(new_n322_), .A3(new_n313_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n319_), .A2(new_n323_), .ZN(new_n324_));
  NAND3_X1  g123(.A1(new_n270_), .A2(new_n300_), .A3(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G127gat), .B(G134gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G113gat), .B(G120gat), .ZN(new_n327_));
  OR2_X1    g126(.A1(new_n326_), .A2(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n326_), .A2(new_n327_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT79), .ZN(new_n331_));
  NAND2_X1  g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332_));
  AND2_X1   g131(.A1(KEYINPUT75), .A2(KEYINPUT23), .ZN(new_n333_));
  NOR2_X1   g132(.A1(KEYINPUT75), .A2(KEYINPUT23), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n332_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n335_));
  OAI21_X1  g134(.A(new_n335_), .B1(KEYINPUT23), .B2(new_n332_), .ZN(new_n336_));
  NOR3_X1   g135(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n337_));
  AND2_X1   g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338_));
  NOR2_X1   g137(.A1(G169gat), .A2(G176gat), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n337_), .B1(new_n340_), .B2(KEYINPUT24), .ZN(new_n341_));
  INV_X1    g140(.A(G183gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n342_), .A2(KEYINPUT25), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT25), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(G183gat), .ZN(new_n345_));
  INV_X1    g144(.A(G190gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n346_), .A2(KEYINPUT26), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT26), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n348_), .A2(G190gat), .ZN(new_n349_));
  NAND4_X1  g148(.A1(new_n343_), .A2(new_n345_), .A3(new_n347_), .A4(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n336_), .A2(new_n341_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n352_));
  AND2_X1   g151(.A1(KEYINPUT76), .A2(G169gat), .ZN(new_n353_));
  NOR2_X1   g152(.A1(KEYINPUT76), .A2(G169gat), .ZN(new_n354_));
  OAI211_X1 g153(.A(new_n352_), .B(KEYINPUT22), .C1(new_n353_), .C2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT22), .ZN(new_n356_));
  AOI21_X1  g155(.A(G176gat), .B1(new_n356_), .B2(G169gat), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n355_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT76), .B(G169gat), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n352_), .B1(new_n359_), .B2(KEYINPUT22), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n332_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n362_), .B1(new_n333_), .B2(new_n334_), .ZN(new_n363_));
  NOR2_X1   g162(.A1(G183gat), .A2(G190gat), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n363_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(G169gat), .A2(G176gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  OAI21_X1  g169(.A(new_n351_), .B1(new_n361_), .B2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT30), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT75), .B(KEYINPUT23), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n366_), .B1(new_n374_), .B2(new_n362_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n338_), .B1(new_n375_), .B2(new_n365_), .ZN(new_n376_));
  OAI21_X1  g175(.A(KEYINPUT22), .B1(new_n353_), .B2(new_n354_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(KEYINPUT77), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n378_), .A2(new_n355_), .A3(new_n357_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT30), .B1(new_n380_), .B2(new_n351_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n331_), .B1(new_n373_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n339_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n383_), .A2(KEYINPUT24), .A3(new_n369_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n337_), .ZN(new_n385_));
  AND3_X1   g184(.A1(new_n350_), .A2(new_n384_), .A3(new_n385_), .ZN(new_n386_));
  AOI22_X1  g185(.A1(new_n376_), .A2(new_n379_), .B1(new_n386_), .B2(new_n336_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(KEYINPUT30), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n371_), .A2(new_n372_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n388_), .A2(KEYINPUT79), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n382_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G227gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(G71gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(G99gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XOR2_X1   g195(.A(G15gat), .B(G43gat), .Z(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT78), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n396_), .B(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n391_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(KEYINPUT31), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n390_), .A2(new_n399_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n399_), .B1(new_n382_), .B2(new_n390_), .ZN(new_n405_));
  AND2_X1   g204(.A1(new_n390_), .A2(new_n399_), .ZN(new_n406_));
  OAI21_X1  g205(.A(KEYINPUT31), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n408_));
  AND3_X1   g207(.A1(new_n404_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n409_));
  AOI21_X1  g208(.A(new_n408_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n330_), .B1(new_n409_), .B2(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n404_), .A2(new_n407_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n412_), .A2(KEYINPUT80), .ZN(new_n413_));
  INV_X1    g212(.A(new_n330_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n404_), .A2(new_n407_), .A3(new_n408_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n413_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(G57gat), .B(G85gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(KEYINPUT94), .ZN(new_n418_));
  INV_X1    g217(.A(G1gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n418_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n421_));
  INV_X1    g220(.A(G29gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n420_), .B(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n426_), .B(KEYINPUT92), .Z(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(G155gat), .A2(G162gat), .ZN(new_n429_));
  NOR2_X1   g228(.A1(G155gat), .A2(G162gat), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n429_), .B1(new_n430_), .B2(KEYINPUT1), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT1), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n432_), .A2(KEYINPUT82), .A3(G155gat), .A4(G162gat), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT82), .ZN(new_n434_));
  OAI21_X1  g233(.A(new_n434_), .B1(new_n429_), .B2(KEYINPUT1), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n431_), .A2(new_n433_), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(G141gat), .ZN(new_n437_));
  INV_X1    g236(.A(G148gat), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n437_), .A2(new_n438_), .A3(KEYINPUT81), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT81), .ZN(new_n440_));
  OAI21_X1  g239(.A(new_n440_), .B1(G141gat), .B2(G148gat), .ZN(new_n441_));
  AOI22_X1  g240(.A1(new_n439_), .A2(new_n441_), .B1(G141gat), .B2(G148gat), .ZN(new_n442_));
  AND2_X1   g241(.A1(new_n436_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n429_), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n444_), .A2(new_n430_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n437_), .A2(new_n438_), .A3(KEYINPUT3), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT3), .ZN(new_n447_));
  OAI21_X1  g246(.A(new_n447_), .B1(G141gat), .B2(G148gat), .ZN(new_n448_));
  AOI21_X1  g247(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n449_));
  AOI22_X1  g248(.A1(new_n446_), .A2(new_n448_), .B1(new_n449_), .B2(KEYINPUT83), .ZN(new_n450_));
  AND3_X1   g249(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(G141gat), .A2(G148gat), .ZN(new_n452_));
  INV_X1    g251(.A(KEYINPUT2), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n452_), .A2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT83), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n451_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n445_), .B1(new_n450_), .B2(new_n456_), .ZN(new_n457_));
  OAI21_X1  g256(.A(KEYINPUT84), .B1(new_n443_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n445_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n446_), .A2(new_n448_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n449_), .A2(KEYINPUT83), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n463_));
  OAI21_X1  g262(.A(new_n463_), .B1(new_n449_), .B2(KEYINPUT83), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n459_), .B1(new_n462_), .B2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(KEYINPUT84), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n436_), .A2(new_n442_), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n458_), .A2(new_n468_), .A3(new_n414_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n443_), .A2(new_n457_), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n330_), .A2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n328_), .A2(KEYINPUT91), .A3(new_n329_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n470_), .A2(new_n472_), .A3(new_n473_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n469_), .A2(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n475_), .A2(KEYINPUT4), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT4), .ZN(new_n477_));
  NAND2_X1  g276(.A1(new_n469_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n428_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n469_), .A2(new_n426_), .A3(new_n474_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n480_), .A2(KEYINPUT95), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT95), .ZN(new_n482_));
  NAND4_X1  g281(.A1(new_n469_), .A2(new_n474_), .A3(new_n482_), .A4(new_n426_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n481_), .A2(new_n483_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n425_), .B1(new_n479_), .B2(new_n484_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n469_), .A2(new_n477_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n477_), .B1(new_n469_), .B2(new_n474_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n427_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n488_), .A2(new_n424_), .A3(new_n481_), .A4(new_n483_), .ZN(new_n489_));
  AND2_X1   g288(.A1(new_n485_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n411_), .A2(new_n416_), .A3(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G8gat), .B(G36gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(G64gat), .B(G92gat), .ZN(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT20), .ZN(new_n498_));
  INV_X1    g297(.A(G218gat), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n499_), .A2(G211gat), .ZN(new_n500_));
  INV_X1    g299(.A(G211gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(G218gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n500_), .A2(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(G197gat), .A2(G204gat), .ZN(new_n504_));
  NOR2_X1   g303(.A1(G197gat), .A2(G204gat), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n504_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT86), .ZN(new_n507_));
  NAND4_X1  g306(.A1(new_n503_), .A2(new_n506_), .A3(new_n507_), .A4(KEYINPUT21), .ZN(new_n508_));
  OR2_X1    g307(.A1(G197gat), .A2(G204gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(G197gat), .A2(G204gat), .ZN(new_n510_));
  NAND4_X1  g309(.A1(new_n509_), .A2(new_n507_), .A3(KEYINPUT21), .A4(new_n510_), .ZN(new_n511_));
  AND2_X1   g310(.A1(new_n500_), .A2(new_n502_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n511_), .A2(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT21), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n515_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(KEYINPUT85), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT85), .ZN(new_n518_));
  OAI211_X1 g317(.A(new_n518_), .B(new_n515_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n506_), .A2(KEYINPUT21), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n517_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n514_), .A2(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n498_), .B1(new_n387_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT89), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT22), .B(G169gat), .ZN(new_n525_));
  INV_X1    g324(.A(G176gat), .ZN(new_n526_));
  AOI21_X1  g325(.A(new_n338_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n332_), .A2(KEYINPUT23), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n528_), .B1(new_n374_), .B2(new_n332_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n527_), .B1(new_n529_), .B2(new_n364_), .ZN(new_n530_));
  INV_X1    g329(.A(KEYINPUT88), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n531_), .A2(KEYINPUT24), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT24), .ZN(new_n533_));
  NOR2_X1   g332(.A1(new_n533_), .A2(KEYINPUT88), .ZN(new_n534_));
  OAI211_X1 g333(.A(new_n369_), .B(new_n383_), .C1(new_n532_), .C2(new_n534_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(KEYINPUT88), .B(KEYINPUT24), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n339_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n375_), .A2(new_n350_), .A3(new_n535_), .A4(new_n537_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n530_), .A2(new_n538_), .ZN(new_n539_));
  OAI21_X1  g338(.A(new_n524_), .B1(new_n539_), .B2(new_n522_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(G226gat), .A2(G233gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT19), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n530_), .A2(new_n538_), .ZN(new_n544_));
  NOR3_X1   g343(.A1(new_n504_), .A2(new_n505_), .A3(new_n515_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n545_), .B1(KEYINPUT85), .B2(new_n516_), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n546_), .A2(new_n519_), .B1(new_n513_), .B2(new_n508_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n544_), .A2(new_n547_), .A3(KEYINPUT89), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n523_), .A2(new_n540_), .A3(new_n543_), .A4(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT98), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  AND3_X1   g350(.A1(new_n544_), .A2(new_n547_), .A3(KEYINPUT89), .ZN(new_n552_));
  AOI21_X1  g351(.A(KEYINPUT89), .B1(new_n544_), .B2(new_n547_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n554_), .A2(KEYINPUT98), .A3(new_n543_), .A4(new_n523_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n551_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n557_));
  OAI21_X1  g356(.A(KEYINPUT20), .B1(new_n544_), .B2(new_n547_), .ZN(new_n558_));
  AOI21_X1  g357(.A(new_n522_), .B1(new_n380_), .B2(new_n351_), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n557_), .B(new_n542_), .C1(new_n558_), .C2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n371_), .A2(new_n547_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n522_), .A2(new_n530_), .A3(new_n538_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n562_), .A2(KEYINPUT20), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n557_), .B1(new_n564_), .B2(new_n542_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n497_), .B1(new_n556_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT99), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  OAI211_X1 g368(.A(KEYINPUT99), .B(new_n497_), .C1(new_n556_), .C2(new_n566_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT27), .ZN(new_n571_));
  NAND4_X1  g370(.A1(new_n562_), .A2(KEYINPUT20), .A3(new_n563_), .A4(new_n543_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n523_), .A2(new_n540_), .A3(new_n548_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n573_), .B1(new_n542_), .B2(new_n574_), .ZN(new_n575_));
  AOI21_X1  g374(.A(new_n571_), .B1(new_n575_), .B2(new_n496_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n569_), .A2(new_n570_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n574_), .A2(new_n542_), .ZN(new_n578_));
  AND3_X1   g377(.A1(new_n578_), .A2(new_n496_), .A3(new_n572_), .ZN(new_n579_));
  AOI21_X1  g378(.A(new_n496_), .B1(new_n578_), .B2(new_n572_), .ZN(new_n580_));
  OAI21_X1  g379(.A(new_n571_), .B1(new_n579_), .B2(new_n580_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT87), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G22gat), .B(G50gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT28), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n458_), .A2(new_n468_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT29), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  AOI211_X1 g387(.A(KEYINPUT29), .B(new_n584_), .C1(new_n458_), .C2(new_n468_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n582_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n458_), .A2(KEYINPUT29), .A3(new_n468_), .ZN(new_n591_));
  AND2_X1   g390(.A1(G228gat), .A2(G233gat), .ZN(new_n592_));
  NOR2_X1   g391(.A1(new_n522_), .A2(new_n592_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n547_), .B1(new_n470_), .B2(new_n587_), .ZN(new_n594_));
  AOI22_X1  g393(.A1(new_n591_), .A2(new_n593_), .B1(new_n594_), .B2(new_n592_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n590_), .A2(new_n595_), .ZN(new_n596_));
  XOR2_X1   g395(.A(G78gat), .B(G106gat), .Z(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NOR2_X1   g397(.A1(new_n588_), .A2(new_n589_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n598_), .B1(new_n599_), .B2(KEYINPUT87), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n443_), .A2(new_n457_), .A3(KEYINPUT84), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n466_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n587_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n584_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n586_), .A2(new_n587_), .A3(new_n585_), .ZN(new_n605_));
  NAND4_X1  g404(.A1(new_n604_), .A2(KEYINPUT87), .A3(new_n605_), .A4(new_n598_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  OAI21_X1  g406(.A(new_n596_), .B1(new_n600_), .B2(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n604_), .A2(KEYINPUT87), .A3(new_n605_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n597_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n610_), .A2(new_n590_), .A3(new_n595_), .A4(new_n606_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n577_), .A2(new_n581_), .A3(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n491_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n570_), .A2(new_n576_), .ZN(new_n616_));
  OAI211_X1 g415(.A(new_n551_), .B(new_n555_), .C1(new_n565_), .C2(new_n561_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT99), .B1(new_n617_), .B2(new_n497_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n616_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n490_), .A2(new_n612_), .A3(new_n581_), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT100), .B1(new_n619_), .B2(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n485_), .A2(new_n489_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n496_), .A2(KEYINPUT32), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n617_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT96), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n575_), .A2(new_n626_), .A3(new_n623_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n578_), .A2(new_n572_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT96), .B1(new_n628_), .B2(new_n624_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n622_), .A2(new_n625_), .A3(new_n627_), .A4(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n579_), .A2(new_n580_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n489_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n484_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n634_), .A2(KEYINPUT33), .A3(new_n424_), .A4(new_n488_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n426_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n425_), .B(new_n636_), .C1(new_n428_), .C2(new_n475_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n631_), .A2(new_n633_), .A3(new_n635_), .A4(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n630_), .A2(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(new_n613_), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n622_), .B1(new_n611_), .B2(new_n608_), .ZN(new_n641_));
  INV_X1    g440(.A(KEYINPUT100), .ZN(new_n642_));
  NAND4_X1  g441(.A1(new_n577_), .A2(new_n641_), .A3(new_n642_), .A4(new_n581_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n621_), .A2(new_n640_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n411_), .A2(new_n416_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n615_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n229_), .A2(new_n230_), .A3(new_n309_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT15), .ZN(new_n650_));
  XNOR2_X1  g449(.A(new_n309_), .B(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n227_), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n649_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT35), .ZN(new_n654_));
  XNOR2_X1  g453(.A(G190gat), .B(G218gat), .ZN(new_n655_));
  XNOR2_X1  g454(.A(G134gat), .B(G162gat), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  AOI22_X1  g456(.A1(new_n653_), .A2(new_n654_), .B1(KEYINPUT36), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(KEYINPUT34), .B(KEYINPUT35), .ZN(new_n659_));
  NAND2_X1  g458(.A1(G232gat), .A2(G233gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n659_), .B(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT69), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n662_), .B1(new_n653_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n317_), .A2(new_n227_), .ZN(new_n665_));
  NAND4_X1  g464(.A1(new_n665_), .A2(KEYINPUT69), .A3(new_n649_), .A4(new_n661_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n658_), .A2(new_n664_), .A3(new_n666_), .ZN(new_n667_));
  NOR2_X1   g466(.A1(new_n657_), .A2(KEYINPUT36), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n668_), .ZN(new_n670_));
  NAND4_X1  g469(.A1(new_n658_), .A2(new_n664_), .A3(new_n670_), .A4(new_n666_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n669_), .A2(new_n671_), .ZN(new_n672_));
  NAND3_X1  g471(.A1(new_n647_), .A2(new_n648_), .A3(new_n672_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n672_), .ZN(new_n674_));
  OAI21_X1  g473(.A(KEYINPUT103), .B1(new_n646_), .B2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n325_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n676_), .A2(KEYINPUT104), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n678_));
  AOI211_X1 g477(.A(new_n678_), .B(new_n325_), .C1(new_n673_), .C2(new_n675_), .ZN(new_n679_));
  NOR2_X1   g478(.A1(new_n677_), .A2(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(G1gat), .B1(new_n680_), .B2(new_n490_), .ZN(new_n681_));
  AND3_X1   g480(.A1(new_n669_), .A2(KEYINPUT37), .A3(new_n671_), .ZN(new_n682_));
  AOI21_X1  g481(.A(KEYINPUT37), .B1(new_n669_), .B2(new_n671_), .ZN(new_n683_));
  AND3_X1   g482(.A1(new_n298_), .A2(KEYINPUT72), .A3(new_n299_), .ZN(new_n684_));
  AOI21_X1  g483(.A(KEYINPUT72), .B1(new_n298_), .B2(new_n299_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n684_), .A2(new_n685_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n682_), .A2(new_n683_), .A3(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n324_), .ZN(new_n689_));
  NOR4_X1   g488(.A1(new_n646_), .A2(new_n688_), .A3(new_n689_), .A4(new_n269_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n622_), .B(KEYINPUT101), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n690_), .A2(new_n419_), .A3(new_n692_), .ZN(new_n693_));
  XOR2_X1   g492(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n694_));
  XNOR2_X1  g493(.A(new_n693_), .B(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n681_), .A2(new_n695_), .ZN(G1324gat));
  INV_X1    g495(.A(G8gat), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n577_), .A2(new_n581_), .ZN(new_n698_));
  NAND3_X1  g497(.A1(new_n690_), .A2(new_n697_), .A3(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT39), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n676_), .A2(new_n698_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(G8gat), .ZN(new_n702_));
  AOI211_X1 g501(.A(KEYINPUT39), .B(new_n697_), .C1(new_n676_), .C2(new_n698_), .ZN(new_n703_));
  OAI21_X1  g502(.A(new_n699_), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(KEYINPUT40), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  OAI211_X1 g505(.A(KEYINPUT40), .B(new_n699_), .C1(new_n702_), .C2(new_n703_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1325gat));
  INV_X1    g507(.A(new_n645_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n690_), .A2(new_n278_), .A3(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n711_));
  AND3_X1   g510(.A1(new_n711_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT41), .B1(new_n711_), .B2(G15gat), .ZN(new_n713_));
  OAI21_X1  g512(.A(new_n710_), .B1(new_n712_), .B2(new_n713_), .ZN(G1326gat));
  NAND3_X1  g513(.A1(new_n690_), .A2(new_n279_), .A3(new_n612_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n612_), .B1(new_n677_), .B2(new_n679_), .ZN(new_n716_));
  XNOR2_X1  g515(.A(KEYINPUT105), .B(KEYINPUT42), .ZN(new_n717_));
  AND3_X1   g516(.A1(new_n716_), .A2(G22gat), .A3(new_n717_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n717_), .B1(new_n716_), .B2(G22gat), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n715_), .B1(new_n718_), .B2(new_n719_), .ZN(G1327gat));
  NOR2_X1   g519(.A1(new_n646_), .A2(new_n689_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n674_), .A2(new_n686_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n269_), .A2(new_n722_), .ZN(new_n723_));
  AND2_X1   g522(.A1(new_n721_), .A2(new_n723_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G29gat), .B1(new_n724_), .B2(new_n622_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n270_), .A2(new_n324_), .A3(new_n686_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n682_), .A2(new_n683_), .ZN(new_n729_));
  INV_X1    g528(.A(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n577_), .A2(new_n641_), .A3(new_n581_), .ZN(new_n731_));
  AOI22_X1  g530(.A1(new_n731_), .A2(KEYINPUT100), .B1(new_n613_), .B2(new_n639_), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n709_), .B1(new_n732_), .B2(new_n643_), .ZN(new_n733_));
  OAI211_X1 g532(.A(new_n728_), .B(new_n730_), .C1(new_n733_), .C2(new_n615_), .ZN(new_n734_));
  OAI21_X1  g533(.A(KEYINPUT43), .B1(new_n646_), .B2(new_n729_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n727_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n726_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  AOI211_X1 g537(.A(KEYINPUT106), .B(new_n727_), .C1(new_n734_), .C2(new_n735_), .ZN(new_n739_));
  NOR2_X1   g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n740_), .B1(KEYINPUT44), .B2(new_n736_), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n691_), .A2(new_n422_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n725_), .B1(new_n741_), .B2(new_n742_), .ZN(G1328gat));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n744_));
  INV_X1    g543(.A(new_n698_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n745_), .B1(new_n736_), .B2(KEYINPUT44), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n746_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n747_));
  AND2_X1   g546(.A1(KEYINPUT107), .A2(G36gat), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n750_));
  NOR2_X1   g549(.A1(new_n745_), .A2(G36gat), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n721_), .A2(new_n750_), .A3(new_n723_), .A4(new_n751_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT107), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n724_), .A2(new_n751_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(KEYINPUT45), .B2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n744_), .B1(new_n749_), .B2(new_n756_), .ZN(new_n757_));
  AOI211_X1 g556(.A(KEYINPUT46), .B(new_n755_), .C1(new_n747_), .C2(new_n748_), .ZN(new_n758_));
  NOR2_X1   g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1329gat));
  NAND2_X1  g558(.A1(new_n736_), .A2(KEYINPUT44), .ZN(new_n760_));
  INV_X1    g559(.A(G43gat), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n645_), .A2(new_n761_), .ZN(new_n762_));
  OAI211_X1 g561(.A(new_n760_), .B(new_n762_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n724_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n764_), .B2(new_n645_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n766_), .A2(KEYINPUT47), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT47), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n763_), .A2(new_n768_), .A3(new_n765_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(G1330gat));
  AOI21_X1  g569(.A(G50gat), .B1(new_n724_), .B2(new_n612_), .ZN(new_n771_));
  AND2_X1   g570(.A1(new_n612_), .A2(G50gat), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n741_), .B2(new_n772_), .ZN(G1331gat));
  NOR4_X1   g572(.A1(new_n646_), .A2(new_n688_), .A3(new_n270_), .A4(new_n324_), .ZN(new_n774_));
  AOI21_X1  g573(.A(G57gat), .B1(new_n774_), .B2(new_n692_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n686_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n269_), .A2(new_n689_), .A3(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n777_), .B1(new_n673_), .B2(new_n675_), .ZN(new_n778_));
  OR2_X1    g577(.A1(new_n778_), .A2(KEYINPUT108), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(KEYINPUT108), .ZN(new_n780_));
  AND2_X1   g579(.A1(new_n779_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(KEYINPUT109), .B(G57gat), .ZN(new_n782_));
  NOR2_X1   g581(.A1(new_n490_), .A2(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n775_), .B1(new_n781_), .B2(new_n783_), .ZN(G1332gat));
  INV_X1    g583(.A(G64gat), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n774_), .A2(new_n785_), .A3(new_n698_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n779_), .A2(new_n698_), .A3(new_n780_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT48), .ZN(new_n788_));
  AND3_X1   g587(.A1(new_n787_), .A2(new_n788_), .A3(G64gat), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n788_), .B1(new_n787_), .B2(G64gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n786_), .B1(new_n789_), .B2(new_n790_), .ZN(G1333gat));
  NAND3_X1  g590(.A1(new_n774_), .A2(new_n393_), .A3(new_n709_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n779_), .A2(new_n709_), .A3(new_n780_), .ZN(new_n793_));
  XOR2_X1   g592(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n794_));
  AND3_X1   g593(.A1(new_n793_), .A2(G71gat), .A3(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n794_), .B1(new_n793_), .B2(G71gat), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n792_), .B1(new_n795_), .B2(new_n796_), .ZN(G1334gat));
  INV_X1    g596(.A(G78gat), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n774_), .A2(new_n798_), .A3(new_n612_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n779_), .A2(new_n612_), .A3(new_n780_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n801_));
  AND3_X1   g600(.A1(new_n800_), .A2(G78gat), .A3(new_n801_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n801_), .B1(new_n800_), .B2(G78gat), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n799_), .B1(new_n802_), .B2(new_n803_), .ZN(G1335gat));
  NOR4_X1   g603(.A1(new_n646_), .A2(new_n324_), .A3(new_n270_), .A4(new_n722_), .ZN(new_n805_));
  AOI21_X1  g604(.A(G85gat), .B1(new_n805_), .B2(new_n692_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n269_), .A2(new_n689_), .A3(new_n686_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n807_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n808_));
  XOR2_X1   g607(.A(new_n808_), .B(KEYINPUT112), .Z(new_n809_));
  AND2_X1   g608(.A1(new_n622_), .A2(new_n212_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n806_), .B1(new_n809_), .B2(new_n810_), .ZN(G1336gat));
  AOI21_X1  g610(.A(G92gat), .B1(new_n805_), .B2(new_n698_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n698_), .A2(G92gat), .ZN(new_n813_));
  XOR2_X1   g612(.A(new_n813_), .B(KEYINPUT113), .Z(new_n814_));
  AOI21_X1  g613(.A(new_n812_), .B1(new_n809_), .B2(new_n814_), .ZN(G1337gat));
  NAND3_X1  g614(.A1(new_n805_), .A2(new_n207_), .A3(new_n709_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n816_), .B(KEYINPUT114), .ZN(new_n817_));
  AOI21_X1  g616(.A(new_n395_), .B1(new_n808_), .B2(new_n709_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  XNOR2_X1  g618(.A(KEYINPUT115), .B(KEYINPUT51), .ZN(new_n820_));
  XNOR2_X1  g619(.A(new_n819_), .B(new_n820_), .ZN(G1338gat));
  NAND3_X1  g620(.A1(new_n805_), .A2(new_n208_), .A3(new_n612_), .ZN(new_n822_));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n808_), .A2(new_n612_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n823_), .B1(new_n824_), .B2(G106gat), .ZN(new_n825_));
  AOI211_X1 g624(.A(KEYINPUT52), .B(new_n208_), .C1(new_n808_), .C2(new_n612_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n822_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  XNOR2_X1  g626(.A(new_n827_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g627(.A1(new_n687_), .A2(new_n268_), .A3(new_n689_), .A4(new_n267_), .ZN(new_n829_));
  XNOR2_X1  g628(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n830_));
  XNOR2_X1  g629(.A(new_n829_), .B(new_n830_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n832_), .A2(KEYINPUT57), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n304_), .B1(new_n314_), .B2(new_n318_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n311_), .B1(new_n285_), .B2(new_n309_), .ZN(new_n835_));
  AOI22_X1  g634(.A1(new_n320_), .A2(new_n835_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n834_), .B1(new_n836_), .B2(new_n304_), .ZN(new_n837_));
  AND2_X1   g636(.A1(new_n265_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT55), .ZN(new_n839_));
  NOR3_X1   g638(.A1(new_n242_), .A2(new_n839_), .A3(new_n244_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n243_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n245_), .A2(new_n839_), .A3(new_n256_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n261_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT56), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(KEYINPUT56), .A3(new_n261_), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n264_), .A2(new_n324_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n850_), .A2(KEYINPUT117), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n264_), .A2(new_n324_), .A3(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n851_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n838_), .B1(new_n849_), .B2(new_n855_), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n833_), .B1(new_n856_), .B2(new_n674_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n833_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n854_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n859_));
  OAI211_X1 g658(.A(new_n672_), .B(new_n858_), .C1(new_n859_), .C2(new_n838_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n837_), .A2(new_n264_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n861_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT58), .ZN(new_n863_));
  INV_X1    g662(.A(new_n861_), .ZN(new_n864_));
  AOI21_X1  g663(.A(KEYINPUT56), .B1(new_n844_), .B2(new_n261_), .ZN(new_n865_));
  AOI211_X1 g664(.A(new_n846_), .B(new_n263_), .C1(new_n842_), .C2(new_n843_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n864_), .B1(new_n865_), .B2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n863_), .A2(new_n869_), .A3(new_n730_), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n857_), .A2(new_n860_), .A3(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n300_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n831_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  NOR3_X1   g672(.A1(new_n614_), .A2(new_n645_), .A3(new_n691_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n875_), .ZN(new_n876_));
  INV_X1    g675(.A(G113gat), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n876_), .A2(new_n877_), .A3(new_n324_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n831_), .B1(new_n871_), .B2(new_n686_), .ZN(new_n879_));
  OR3_X1    g678(.A1(new_n879_), .A2(KEYINPUT59), .A3(new_n875_), .ZN(new_n880_));
  OAI21_X1  g679(.A(KEYINPUT59), .B1(new_n873_), .B2(new_n875_), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n880_), .A2(new_n324_), .A3(new_n881_), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n878_), .B1(new_n882_), .B2(new_n877_), .ZN(G1340gat));
  NAND3_X1  g682(.A1(new_n880_), .A2(new_n269_), .A3(new_n881_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(G120gat), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT60), .ZN(new_n886_));
  AOI21_X1  g685(.A(G120gat), .B1(new_n269_), .B2(new_n886_), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n887_), .A2(KEYINPUT119), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n889_), .B1(new_n886_), .B2(G120gat), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n876_), .B(new_n888_), .C1(new_n887_), .C2(new_n890_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n885_), .A2(new_n891_), .ZN(G1341gat));
  INV_X1    g691(.A(G127gat), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n876_), .A2(new_n893_), .A3(new_n776_), .ZN(new_n894_));
  AND3_X1   g693(.A1(new_n880_), .A2(new_n300_), .A3(new_n881_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n893_), .ZN(G1342gat));
  INV_X1    g695(.A(G134gat), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n876_), .A2(new_n897_), .A3(new_n674_), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n880_), .A2(new_n730_), .A3(new_n881_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n898_), .B1(new_n899_), .B2(new_n897_), .ZN(G1343gat));
  NOR4_X1   g699(.A1(new_n709_), .A2(new_n698_), .A3(new_n691_), .A4(new_n613_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n873_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n324_), .ZN(new_n904_));
  XOR2_X1   g703(.A(KEYINPUT120), .B(G141gat), .Z(new_n905_));
  XNOR2_X1  g704(.A(new_n904_), .B(new_n905_), .ZN(G1344gat));
  NAND2_X1  g705(.A1(new_n903_), .A2(new_n269_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g707(.A1(new_n903_), .A2(new_n776_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(KEYINPUT61), .B(G155gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n909_), .B(new_n910_), .ZN(G1346gat));
  NAND2_X1  g710(.A1(new_n871_), .A2(new_n872_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n831_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(new_n901_), .ZN(new_n915_));
  OAI21_X1  g714(.A(G162gat), .B1(new_n915_), .B2(new_n729_), .ZN(new_n916_));
  NOR4_X1   g715(.A1(new_n873_), .A2(G162gat), .A3(new_n672_), .A4(new_n902_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n916_), .A2(new_n918_), .A3(KEYINPUT121), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n920_));
  INV_X1    g719(.A(G162gat), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n921_), .B1(new_n903_), .B2(new_n730_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n920_), .B1(new_n922_), .B2(new_n917_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n919_), .A2(new_n923_), .ZN(G1347gat));
  NAND3_X1  g723(.A1(new_n709_), .A2(new_n698_), .A3(new_n691_), .ZN(new_n925_));
  NOR3_X1   g724(.A1(new_n879_), .A2(new_n612_), .A3(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n926_), .A2(new_n525_), .A3(new_n324_), .ZN(new_n927_));
  INV_X1    g726(.A(KEYINPUT62), .ZN(new_n928_));
  INV_X1    g727(.A(G169gat), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n925_), .A2(new_n689_), .ZN(new_n930_));
  XNOR2_X1  g729(.A(new_n930_), .B(KEYINPUT122), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n931_), .A2(new_n613_), .ZN(new_n932_));
  NAND2_X1  g731(.A1(new_n871_), .A2(new_n686_), .ZN(new_n933_));
  AOI21_X1  g732(.A(new_n932_), .B1(new_n933_), .B2(new_n913_), .ZN(new_n934_));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n929_), .B1(new_n934_), .B2(new_n935_), .ZN(new_n936_));
  OAI21_X1  g735(.A(KEYINPUT123), .B1(new_n879_), .B2(new_n932_), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n928_), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  AND2_X1   g737(.A1(new_n931_), .A2(new_n613_), .ZN(new_n939_));
  OAI21_X1  g738(.A(new_n672_), .B1(new_n859_), .B2(new_n838_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n729_), .B1(new_n862_), .B2(KEYINPUT58), .ZN(new_n941_));
  AOI22_X1  g740(.A1(new_n940_), .A2(new_n833_), .B1(new_n941_), .B2(new_n869_), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n776_), .B1(new_n942_), .B2(new_n860_), .ZN(new_n943_));
  OAI211_X1 g742(.A(new_n935_), .B(new_n939_), .C1(new_n943_), .C2(new_n831_), .ZN(new_n944_));
  AND4_X1   g743(.A1(new_n928_), .A2(new_n937_), .A3(new_n944_), .A4(G169gat), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n927_), .B1(new_n938_), .B2(new_n945_), .ZN(G1348gat));
  NOR3_X1   g745(.A1(new_n873_), .A2(new_n612_), .A3(new_n925_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n270_), .A2(new_n526_), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n947_), .A2(new_n948_), .A3(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(G176gat), .B1(new_n926_), .B2(new_n269_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n948_), .B1(new_n947_), .B2(new_n949_), .ZN(new_n952_));
  NOR3_X1   g751(.A1(new_n950_), .A2(new_n951_), .A3(new_n952_), .ZN(G1349gat));
  AOI21_X1  g752(.A(G183gat), .B1(new_n947_), .B2(new_n776_), .ZN(new_n954_));
  AOI21_X1  g753(.A(new_n872_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n954_), .B1(new_n926_), .B2(new_n955_), .ZN(G1350gat));
  NAND4_X1  g755(.A1(new_n926_), .A2(new_n674_), .A3(new_n347_), .A4(new_n349_), .ZN(new_n957_));
  AND2_X1   g756(.A1(new_n926_), .A2(new_n730_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n957_), .B1(new_n958_), .B2(new_n346_), .ZN(G1351gat));
  XNOR2_X1  g758(.A(KEYINPUT126), .B(G197gat), .ZN(new_n960_));
  NAND3_X1  g759(.A1(new_n645_), .A2(new_n698_), .A3(new_n641_), .ZN(new_n961_));
  INV_X1    g760(.A(new_n961_), .ZN(new_n962_));
  NAND3_X1  g761(.A1(new_n914_), .A2(KEYINPUT125), .A3(new_n962_), .ZN(new_n963_));
  INV_X1    g762(.A(KEYINPUT125), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n964_), .B1(new_n873_), .B2(new_n961_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n963_), .A2(new_n965_), .ZN(new_n966_));
  AOI21_X1  g765(.A(new_n960_), .B1(new_n966_), .B2(new_n324_), .ZN(new_n967_));
  INV_X1    g766(.A(new_n960_), .ZN(new_n968_));
  AOI211_X1 g767(.A(new_n689_), .B(new_n968_), .C1(new_n963_), .C2(new_n965_), .ZN(new_n969_));
  NOR2_X1   g768(.A1(new_n967_), .A2(new_n969_), .ZN(G1352gat));
  AOI21_X1  g769(.A(KEYINPUT125), .B1(new_n914_), .B2(new_n962_), .ZN(new_n971_));
  NOR3_X1   g770(.A1(new_n873_), .A2(new_n964_), .A3(new_n961_), .ZN(new_n972_));
  OAI21_X1  g771(.A(new_n269_), .B1(new_n971_), .B2(new_n972_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n973_), .A2(G204gat), .ZN(new_n974_));
  INV_X1    g773(.A(G204gat), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n966_), .A2(new_n975_), .A3(new_n269_), .ZN(new_n976_));
  NAND2_X1  g775(.A1(new_n974_), .A2(new_n976_), .ZN(G1353gat));
  OR2_X1    g776(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n978_), .B1(new_n966_), .B2(new_n300_), .ZN(new_n979_));
  XNOR2_X1  g778(.A(KEYINPUT63), .B(G211gat), .ZN(new_n980_));
  AOI211_X1 g779(.A(new_n872_), .B(new_n980_), .C1(new_n963_), .C2(new_n965_), .ZN(new_n981_));
  NOR2_X1   g780(.A1(new_n979_), .A2(new_n981_), .ZN(G1354gat));
  NAND3_X1  g781(.A1(new_n966_), .A2(new_n499_), .A3(new_n674_), .ZN(new_n983_));
  AOI21_X1  g782(.A(new_n729_), .B1(new_n963_), .B2(new_n965_), .ZN(new_n984_));
  OAI21_X1  g783(.A(new_n983_), .B1(new_n499_), .B2(new_n984_), .ZN(G1355gat));
endmodule


