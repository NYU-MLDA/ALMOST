//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 0 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n650_, new_n651_, new_n652_, new_n653_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n721_, new_n722_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n766_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n908_, new_n909_, new_n910_,
    new_n912_, new_n913_, new_n914_, new_n915_, new_n916_, new_n917_,
    new_n919_, new_n920_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_;
  XNOR2_X1  g000(.A(G211gat), .B(G218gat), .ZN(new_n202_));
  OR2_X1    g001(.A1(KEYINPUT93), .A2(G204gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(KEYINPUT93), .A2(G204gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n205_), .A2(G197gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT21), .ZN(new_n207_));
  AOI21_X1  g006(.A(new_n207_), .B1(G197gat), .B2(G204gat), .ZN(new_n208_));
  INV_X1    g007(.A(new_n208_), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G197gat), .A2(G204gat), .ZN(new_n210_));
  AOI21_X1  g009(.A(new_n210_), .B1(new_n205_), .B2(G197gat), .ZN(new_n211_));
  OAI221_X1 g010(.A(new_n202_), .B1(new_n206_), .B2(new_n209_), .C1(KEYINPUT21), .C2(new_n211_), .ZN(new_n212_));
  NOR2_X1   g011(.A1(new_n202_), .A2(new_n207_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(G141gat), .ZN(new_n216_));
  INV_X1    g015(.A(G148gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  OAI21_X1  g017(.A(new_n218_), .B1(KEYINPUT89), .B2(KEYINPUT3), .ZN(new_n219_));
  NOR2_X1   g018(.A1(KEYINPUT89), .A2(KEYINPUT3), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n220_), .A2(new_n216_), .A3(new_n217_), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n222_), .B1(new_n216_), .B2(new_n217_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n219_), .A2(new_n221_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(G155gat), .A2(G162gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n227_), .A2(KEYINPUT86), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT86), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n229_), .A2(G155gat), .A3(G162gat), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n226_), .B1(new_n228_), .B2(new_n230_), .ZN(new_n231_));
  AND3_X1   g030(.A1(new_n225_), .A2(KEYINPUT90), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(KEYINPUT90), .B1(new_n225_), .B2(new_n231_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n232_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT88), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n228_), .A2(new_n230_), .ZN(new_n236_));
  OAI22_X1  g035(.A1(new_n236_), .A2(KEYINPUT1), .B1(G155gat), .B2(G162gat), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT87), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n228_), .A2(new_n230_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT1), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n238_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n236_), .A2(KEYINPUT87), .A3(KEYINPUT1), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n237_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n218_), .A2(KEYINPUT85), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n218_), .A2(KEYINPUT85), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n244_), .A2(new_n245_), .B1(G141gat), .B2(G148gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n235_), .B1(new_n243_), .B2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(KEYINPUT87), .B1(new_n236_), .B2(KEYINPUT1), .ZN(new_n249_));
  AOI211_X1 g048(.A(new_n238_), .B(new_n240_), .C1(new_n228_), .C2(new_n230_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  OAI211_X1 g050(.A(KEYINPUT88), .B(new_n246_), .C1(new_n251_), .C2(new_n237_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n234_), .B1(new_n248_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT29), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n215_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G228gat), .A2(G233gat), .ZN(new_n256_));
  OR2_X1    g055(.A1(new_n211_), .A2(KEYINPUT21), .ZN(new_n257_));
  INV_X1    g056(.A(new_n202_), .ZN(new_n258_));
  AND2_X1   g057(.A1(new_n203_), .A2(new_n204_), .ZN(new_n259_));
  INV_X1    g058(.A(G197gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n258_), .B1(new_n261_), .B2(new_n208_), .ZN(new_n262_));
  AOI22_X1  g061(.A1(new_n257_), .A2(new_n262_), .B1(new_n211_), .B2(new_n213_), .ZN(new_n263_));
  OAI21_X1  g062(.A(new_n256_), .B1(new_n263_), .B2(KEYINPUT92), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n255_), .B(new_n264_), .ZN(new_n265_));
  INV_X1    g064(.A(new_n265_), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  XOR2_X1   g067(.A(G22gat), .B(G50gat), .Z(new_n269_));
  INV_X1    g068(.A(new_n269_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n253_), .A2(new_n254_), .A3(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n270_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n268_), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G78gat), .B(G106gat), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n248_), .A2(new_n252_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n234_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n277_), .A2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n269_), .B1(new_n279_), .B2(KEYINPUT29), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(new_n267_), .A3(new_n271_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n274_), .A2(new_n276_), .A3(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n276_), .B1(new_n274_), .B2(new_n281_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n266_), .B1(new_n283_), .B2(new_n284_), .ZN(new_n285_));
  NOR3_X1   g084(.A1(new_n272_), .A2(new_n268_), .A3(new_n273_), .ZN(new_n286_));
  AOI21_X1  g085(.A(new_n267_), .B1(new_n280_), .B2(new_n271_), .ZN(new_n287_));
  OAI21_X1  g086(.A(new_n275_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(new_n265_), .A3(new_n282_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  XOR2_X1   g089(.A(G8gat), .B(G36gat), .Z(new_n291_));
  XNOR2_X1  g090(.A(new_n291_), .B(KEYINPUT18), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G64gat), .B(G92gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(G183gat), .ZN(new_n295_));
  INV_X1    g094(.A(G190gat), .ZN(new_n296_));
  OAI21_X1  g095(.A(KEYINPUT23), .B1(new_n295_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT23), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n298_), .A2(G183gat), .A3(G190gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n297_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n300_), .B1(G183gat), .B2(G190gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT22), .B(G169gat), .ZN(new_n302_));
  INV_X1    g101(.A(G176gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n302_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT95), .ZN(new_n306_));
  INV_X1    g105(.A(KEYINPUT96), .ZN(new_n307_));
  AND3_X1   g106(.A1(new_n304_), .A2(new_n306_), .A3(new_n307_), .ZN(new_n308_));
  AOI21_X1  g107(.A(new_n307_), .B1(new_n304_), .B2(new_n306_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n301_), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n305_), .A2(KEYINPUT24), .ZN(new_n311_));
  NOR2_X1   g110(.A1(G169gat), .A2(G176gat), .ZN(new_n312_));
  MUX2_X1   g111(.A(new_n311_), .B(KEYINPUT24), .S(new_n312_), .Z(new_n313_));
  OR2_X1    g112(.A1(new_n299_), .A2(KEYINPUT82), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n297_), .A2(KEYINPUT82), .A3(new_n299_), .ZN(new_n315_));
  AND2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT25), .B(G183gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n317_), .B(KEYINPUT94), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT26), .B(G190gat), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  OAI211_X1 g119(.A(new_n313_), .B(new_n316_), .C1(new_n318_), .C2(new_n320_), .ZN(new_n321_));
  NAND3_X1  g120(.A1(new_n263_), .A2(new_n310_), .A3(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n323_), .B(G169gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n314_), .A2(new_n315_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G183gat), .A2(G190gat), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n324_), .B1(new_n325_), .B2(new_n326_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT81), .ZN(new_n328_));
  NOR2_X1   g127(.A1(new_n317_), .A2(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n328_), .B1(new_n295_), .B2(KEYINPUT25), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n319_), .A2(new_n330_), .ZN(new_n331_));
  OAI211_X1 g130(.A(new_n313_), .B(new_n300_), .C1(new_n329_), .C2(new_n331_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n327_), .A2(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n215_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G226gat), .A2(G233gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n335_), .B(KEYINPUT19), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n322_), .A2(new_n334_), .A3(KEYINPUT20), .A4(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT20), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n310_), .A2(new_n321_), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(new_n215_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n263_), .A2(new_n332_), .A3(new_n327_), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n294_), .B(new_n338_), .C1(new_n343_), .C2(new_n337_), .ZN(new_n344_));
  INV_X1    g143(.A(new_n294_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n338_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n337_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n345_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT27), .B1(new_n344_), .B2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT99), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n344_), .A2(KEYINPUT27), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n294_), .B(KEYINPUT98), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n322_), .A2(new_n334_), .A3(KEYINPUT20), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n353_), .A2(new_n336_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n341_), .A2(new_n342_), .A3(new_n337_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n352_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n356_));
  OAI21_X1  g155(.A(new_n350_), .B1(new_n351_), .B2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n356_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n358_), .A2(new_n344_), .A3(KEYINPUT99), .A4(KEYINPUT27), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n349_), .B1(new_n357_), .B2(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n290_), .A2(new_n360_), .ZN(new_n361_));
  XOR2_X1   g160(.A(G127gat), .B(G134gat), .Z(new_n362_));
  XOR2_X1   g161(.A(G113gat), .B(G120gat), .Z(new_n363_));
  XOR2_X1   g162(.A(new_n362_), .B(new_n363_), .Z(new_n364_));
  NAND2_X1  g163(.A1(new_n279_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n364_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n253_), .A2(new_n366_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(G225gat), .A2(G233gat), .ZN(new_n368_));
  NAND3_X1  g167(.A1(new_n365_), .A2(new_n367_), .A3(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(G1gat), .B(G29gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n370_), .B(G85gat), .ZN(new_n371_));
  XNOR2_X1  g170(.A(KEYINPUT0), .B(G57gat), .ZN(new_n372_));
  XOR2_X1   g171(.A(new_n371_), .B(new_n372_), .Z(new_n373_));
  NOR2_X1   g172(.A1(new_n253_), .A2(new_n366_), .ZN(new_n374_));
  AOI211_X1 g173(.A(new_n364_), .B(new_n234_), .C1(new_n248_), .C2(new_n252_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT4), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n374_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n279_), .A2(new_n376_), .A3(new_n364_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n368_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n378_), .A2(new_n379_), .ZN(new_n380_));
  OAI211_X1 g179(.A(new_n369_), .B(new_n373_), .C1(new_n377_), .C2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n365_), .A2(KEYINPUT4), .A3(new_n367_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n383_), .A2(new_n379_), .A3(new_n378_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n373_), .B1(new_n384_), .B2(new_n369_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n382_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G71gat), .B(G99gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(KEYINPUT83), .B(G43gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  XNOR2_X1  g188(.A(new_n333_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(new_n364_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(G227gat), .A2(G233gat), .ZN(new_n392_));
  INV_X1    g191(.A(G15gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n392_), .B(new_n393_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT30), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n395_), .B(KEYINPUT31), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n391_), .B(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n386_), .A2(new_n398_), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n361_), .A2(new_n399_), .ZN(new_n400_));
  NAND4_X1  g199(.A1(new_n360_), .A2(new_n285_), .A3(new_n386_), .A4(new_n289_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n346_), .A2(new_n347_), .ZN(new_n402_));
  AND2_X1   g201(.A1(new_n294_), .A2(KEYINPUT32), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n402_), .A2(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n354_), .A2(new_n355_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(new_n403_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n405_), .A2(new_n407_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n369_), .B1(new_n377_), .B2(new_n380_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n373_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n408_), .B1(new_n411_), .B2(new_n381_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT33), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n381_), .A2(new_n413_), .ZN(new_n414_));
  NAND4_X1  g213(.A1(new_n384_), .A2(KEYINPUT33), .A3(new_n369_), .A4(new_n373_), .ZN(new_n415_));
  AND2_X1   g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n344_), .A2(new_n348_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n365_), .A2(new_n367_), .A3(new_n379_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(new_n410_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n379_), .B1(new_n374_), .B2(new_n376_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n383_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT97), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n419_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n383_), .A2(new_n420_), .A3(KEYINPUT97), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n417_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  AOI21_X1  g224(.A(new_n412_), .B1(new_n416_), .B2(new_n425_), .ZN(new_n426_));
  INV_X1    g225(.A(new_n290_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n401_), .B1(new_n426_), .B2(new_n427_), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n397_), .B(KEYINPUT84), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n400_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G29gat), .B(G36gat), .Z(new_n431_));
  XOR2_X1   g230(.A(G43gat), .B(G50gat), .Z(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n433_), .B(KEYINPUT15), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G15gat), .B(G22gat), .ZN(new_n435_));
  INV_X1    g234(.A(G1gat), .ZN(new_n436_));
  INV_X1    g235(.A(G8gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT14), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT79), .ZN(new_n439_));
  OAI21_X1  g238(.A(new_n435_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n438_), .A2(new_n439_), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G1gat), .B(G8gat), .ZN(new_n442_));
  OR3_X1    g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n442_), .B1(new_n440_), .B2(new_n441_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n434_), .A2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n433_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(G229gat), .A2(G233gat), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n449_), .A3(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n450_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n433_), .B1(new_n443_), .B2(new_n444_), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n452_), .B1(new_n448_), .B2(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n451_), .A2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G113gat), .B(G141gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G169gat), .B(G197gat), .ZN(new_n457_));
  XOR2_X1   g256(.A(new_n456_), .B(new_n457_), .Z(new_n458_));
  INV_X1    g257(.A(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n455_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n451_), .A2(new_n454_), .A3(new_n458_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n460_), .A2(new_n461_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT80), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n460_), .A2(KEYINPUT80), .A3(new_n461_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n464_), .A2(new_n465_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n430_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT37), .ZN(new_n468_));
  NOR2_X1   g267(.A1(G85gat), .A2(G92gat), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G85gat), .A2(G92gat), .ZN(new_n470_));
  INV_X1    g269(.A(KEYINPUT9), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n470_), .A2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT65), .ZN(new_n473_));
  INV_X1    g272(.A(new_n470_), .ZN(new_n474_));
  OAI21_X1  g273(.A(new_n473_), .B1(new_n474_), .B2(KEYINPUT9), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n470_), .A2(KEYINPUT65), .A3(new_n471_), .ZN(new_n476_));
  AOI211_X1 g275(.A(new_n469_), .B(new_n472_), .C1(new_n475_), .C2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(G99gat), .ZN(new_n478_));
  INV_X1    g277(.A(G106gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT6), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(G99gat), .A3(G106gat), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(KEYINPUT10), .B(G99gat), .ZN(new_n484_));
  XNOR2_X1  g283(.A(KEYINPUT64), .B(G106gat), .ZN(new_n485_));
  OAI21_X1  g284(.A(new_n483_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n477_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT68), .ZN(new_n488_));
  NOR2_X1   g287(.A1(G99gat), .A2(G106gat), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT66), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT7), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT66), .ZN(new_n493_));
  AOI21_X1  g292(.A(new_n489_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n494_));
  AOI211_X1 g293(.A(G99gat), .B(G106gat), .C1(new_n490_), .C2(KEYINPUT7), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n488_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n491_), .A2(new_n489_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(KEYINPUT66), .B(KEYINPUT7), .ZN(new_n498_));
  OAI211_X1 g297(.A(KEYINPUT68), .B(new_n497_), .C1(new_n498_), .C2(new_n489_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT67), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n480_), .A2(new_n482_), .A3(new_n500_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n483_), .A2(KEYINPUT67), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n496_), .A2(new_n499_), .A3(new_n501_), .A4(new_n502_), .ZN(new_n503_));
  NOR2_X1   g302(.A1(new_n474_), .A2(new_n469_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n505_), .A2(KEYINPUT8), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n483_), .B(new_n497_), .C1(new_n489_), .C2(new_n498_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT8), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n507_), .A2(new_n508_), .A3(new_n504_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n487_), .B1(new_n506_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT35), .ZN(new_n511_));
  NAND2_X1  g310(.A1(G232gat), .A2(G233gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n512_), .B(KEYINPUT34), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  AOI22_X1  g313(.A1(new_n510_), .A2(new_n433_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n515_));
  NOR2_X1   g314(.A1(new_n514_), .A2(new_n511_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n487_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n508_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n509_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n521_), .A2(new_n434_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n515_), .A2(new_n517_), .A3(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n522_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n514_), .A2(new_n511_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n525_), .B1(new_n521_), .B2(new_n447_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n516_), .B1(new_n524_), .B2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n523_), .A2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G190gat), .B(G218gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(new_n529_), .B(KEYINPUT75), .ZN(new_n530_));
  XNOR2_X1  g329(.A(G134gat), .B(G162gat), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n532_), .A2(new_n533_), .ZN(new_n534_));
  XOR2_X1   g333(.A(new_n534_), .B(KEYINPUT76), .Z(new_n535_));
  NOR2_X1   g334(.A1(new_n528_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n532_), .B(new_n533_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n528_), .A2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n468_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT77), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n538_), .B1(new_n528_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n523_), .A2(new_n527_), .A3(KEYINPUT77), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n536_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  AOI21_X1  g345(.A(KEYINPUT78), .B1(new_n546_), .B2(new_n468_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n517_), .B1(new_n515_), .B2(new_n522_), .ZN(new_n548_));
  NOR3_X1   g347(.A1(new_n524_), .A2(new_n526_), .A3(new_n516_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n543_), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(new_n539_), .A3(new_n545_), .ZN(new_n551_));
  AND4_X1   g350(.A1(KEYINPUT78), .A2(new_n551_), .A3(new_n468_), .A4(new_n537_), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n542_), .B1(new_n547_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n554_));
  XNOR2_X1  g353(.A(G127gat), .B(G155gat), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT16), .ZN(new_n556_));
  XOR2_X1   g355(.A(G183gat), .B(G211gat), .Z(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  AND2_X1   g357(.A1(G231gat), .A2(G233gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n445_), .B(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G57gat), .B(G64gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G71gat), .B(G78gat), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n561_), .A2(new_n562_), .A3(KEYINPUT11), .ZN(new_n563_));
  INV_X1    g362(.A(new_n562_), .ZN(new_n564_));
  INV_X1    g363(.A(G64gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(G57gat), .ZN(new_n566_));
  INV_X1    g365(.A(G57gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(G64gat), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n566_), .A2(new_n568_), .A3(KEYINPUT11), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n561_), .A2(KEYINPUT11), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n563_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT71), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  AOI211_X1 g373(.A(new_n554_), .B(new_n558_), .C1(new_n560_), .C2(new_n574_), .ZN(new_n575_));
  OAI21_X1  g374(.A(new_n575_), .B1(new_n574_), .B2(new_n560_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n558_), .B(new_n554_), .ZN(new_n577_));
  INV_X1    g376(.A(new_n560_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT69), .ZN(new_n579_));
  OAI211_X1 g378(.A(new_n579_), .B(new_n563_), .C1(new_n570_), .C2(new_n571_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n566_), .A2(new_n568_), .ZN(new_n582_));
  INV_X1    g381(.A(KEYINPUT11), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n584_), .A2(new_n569_), .A3(new_n564_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n579_), .B1(new_n585_), .B2(new_n563_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n577_), .B1(new_n578_), .B2(new_n588_), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n589_), .B1(new_n578_), .B2(new_n588_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n576_), .A2(new_n590_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n587_), .B(new_n518_), .C1(new_n519_), .C2(new_n520_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n574_), .A2(KEYINPUT12), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n592_), .B1(new_n510_), .B2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(G230gat), .A2(G233gat), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AOI21_X1  g395(.A(KEYINPUT12), .B1(new_n521_), .B2(new_n588_), .ZN(new_n597_));
  OR3_X1    g396(.A1(new_n594_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n521_), .A2(new_n588_), .ZN(new_n599_));
  INV_X1    g398(.A(KEYINPUT70), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n599_), .A2(new_n600_), .A3(new_n592_), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n601_), .B(new_n596_), .C1(new_n600_), .C2(new_n599_), .ZN(new_n602_));
  XOR2_X1   g401(.A(G176gat), .B(G204gat), .Z(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT73), .ZN(new_n604_));
  XOR2_X1   g403(.A(G120gat), .B(G148gat), .Z(new_n605_));
  XNOR2_X1  g404(.A(new_n604_), .B(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n606_), .B(new_n607_), .Z(new_n608_));
  NAND3_X1  g407(.A1(new_n598_), .A2(new_n602_), .A3(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  AOI21_X1  g409(.A(new_n608_), .B1(new_n598_), .B2(new_n602_), .ZN(new_n611_));
  XOR2_X1   g410(.A(KEYINPUT74), .B(KEYINPUT13), .Z(new_n612_));
  OR3_X1    g411(.A1(new_n610_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  OAI22_X1  g412(.A1(new_n610_), .A2(new_n611_), .B1(KEYINPUT74), .B2(KEYINPUT13), .ZN(new_n614_));
  AOI21_X1  g413(.A(new_n591_), .B1(new_n613_), .B2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n467_), .A2(new_n553_), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(KEYINPUT100), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n616_), .B(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n386_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n618_), .A2(new_n436_), .A3(new_n619_), .ZN(new_n620_));
  XNOR2_X1  g419(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n621_));
  OR2_X1    g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n621_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n430_), .A2(new_n546_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n613_), .A2(new_n614_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n466_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  NOR2_X1   g426(.A1(new_n627_), .A2(new_n591_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n624_), .A2(new_n628_), .ZN(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(new_n619_), .ZN(new_n630_));
  OAI211_X1 g429(.A(new_n622_), .B(new_n623_), .C1(new_n436_), .C2(new_n630_), .ZN(G1324gat));
  INV_X1    g430(.A(new_n360_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n624_), .A2(new_n632_), .A3(new_n628_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(G8gat), .ZN(new_n634_));
  AND2_X1   g433(.A1(new_n634_), .A2(KEYINPUT102), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(KEYINPUT102), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT39), .ZN(new_n637_));
  OR3_X1    g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n360_), .A2(G8gat), .ZN(new_n639_));
  AOI22_X1  g438(.A1(new_n618_), .A2(new_n639_), .B1(new_n635_), .B2(new_n637_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n641_));
  AND3_X1   g440(.A1(new_n638_), .A2(new_n640_), .A3(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n641_), .B1(new_n638_), .B2(new_n640_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1325gat));
  INV_X1    g443(.A(new_n429_), .ZN(new_n645_));
  AOI21_X1  g444(.A(new_n393_), .B1(new_n629_), .B2(new_n645_), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n646_), .B(KEYINPUT41), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n618_), .A2(new_n393_), .A3(new_n645_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n647_), .A2(new_n648_), .ZN(G1326gat));
  INV_X1    g448(.A(G22gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n650_), .B1(new_n629_), .B2(new_n427_), .ZN(new_n651_));
  XOR2_X1   g450(.A(new_n651_), .B(KEYINPUT42), .Z(new_n652_));
  NAND3_X1  g451(.A1(new_n618_), .A2(new_n650_), .A3(new_n427_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1327gat));
  INV_X1    g453(.A(new_n546_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n591_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n655_), .A2(new_n656_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n625_), .A2(new_n657_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n467_), .A2(KEYINPUT105), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n401_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n421_), .A2(new_n422_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n419_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n661_), .A2(new_n424_), .A3(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(new_n417_), .ZN(new_n664_));
  NAND4_X1  g463(.A1(new_n663_), .A2(new_n414_), .A3(new_n664_), .A4(new_n415_), .ZN(new_n665_));
  OAI211_X1 g464(.A(new_n407_), .B(new_n405_), .C1(new_n382_), .C2(new_n385_), .ZN(new_n666_));
  AOI22_X1  g465(.A1(new_n665_), .A2(new_n666_), .B1(new_n289_), .B2(new_n285_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n429_), .B1(new_n660_), .B2(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(new_n400_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n670_), .A2(new_n626_), .A3(new_n658_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n659_), .A2(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(G29gat), .B1(new_n675_), .B2(new_n619_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT104), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n553_), .A2(new_n677_), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n551_), .A2(new_n537_), .A3(new_n468_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT78), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n546_), .A2(KEYINPUT78), .A3(new_n468_), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n541_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT104), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n678_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(KEYINPUT43), .B1(new_n685_), .B2(new_n430_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n681_), .A2(new_n682_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n687_), .A2(new_n688_), .A3(new_n542_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n689_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n686_), .A2(new_n691_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n627_), .A2(new_n656_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n692_), .A2(KEYINPUT44), .A3(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT44), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n665_), .A2(new_n666_), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n696_), .A2(new_n290_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n645_), .B1(new_n697_), .B2(new_n401_), .ZN(new_n698_));
  OAI211_X1 g497(.A(new_n678_), .B(new_n684_), .C1(new_n698_), .C2(new_n400_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n690_), .B1(new_n699_), .B2(KEYINPUT43), .ZN(new_n700_));
  INV_X1    g499(.A(new_n693_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n695_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n694_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AND2_X1   g503(.A1(new_n619_), .A2(G29gat), .ZN(new_n705_));
  AOI21_X1  g504(.A(new_n676_), .B1(new_n704_), .B2(new_n705_), .ZN(G1328gat));
  OAI21_X1  g505(.A(G36gat), .B1(new_n703_), .B2(new_n360_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n360_), .A2(G36gat), .ZN(new_n708_));
  NAND3_X1  g507(.A1(new_n659_), .A2(new_n673_), .A3(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT45), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n707_), .A2(new_n710_), .A3(KEYINPUT106), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n712_));
  AOI21_X1  g511(.A(KEYINPUT46), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(KEYINPUT46), .ZN(new_n714_));
  AOI22_X1  g513(.A1(new_n707_), .A2(new_n710_), .B1(KEYINPUT106), .B2(new_n714_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n713_), .A2(new_n715_), .ZN(G1329gat));
  NAND2_X1  g515(.A1(new_n398_), .A2(G43gat), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n674_), .A2(new_n429_), .ZN(new_n718_));
  OAI22_X1  g517(.A1(new_n703_), .A2(new_n717_), .B1(new_n718_), .B2(G43gat), .ZN(new_n719_));
  XNOR2_X1  g518(.A(new_n719_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g519(.A(G50gat), .B1(new_n675_), .B2(new_n427_), .ZN(new_n721_));
  AND2_X1   g520(.A1(new_n427_), .A2(G50gat), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n704_), .B2(new_n722_), .ZN(G1331gat));
  INV_X1    g522(.A(new_n625_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(new_n656_), .ZN(new_n725_));
  NOR4_X1   g524(.A1(new_n430_), .A2(new_n626_), .A3(new_n683_), .A4(new_n725_), .ZN(new_n726_));
  NAND3_X1  g525(.A1(new_n726_), .A2(new_n567_), .A3(new_n619_), .ZN(new_n727_));
  NOR4_X1   g526(.A1(new_n430_), .A2(new_n626_), .A3(new_n546_), .A4(new_n725_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n728_), .A2(new_n619_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n729_), .B2(new_n567_), .ZN(G1332gat));
  AOI21_X1  g529(.A(new_n565_), .B1(new_n728_), .B2(new_n632_), .ZN(new_n731_));
  XOR2_X1   g530(.A(new_n731_), .B(KEYINPUT48), .Z(new_n732_));
  NAND3_X1  g531(.A1(new_n726_), .A2(new_n565_), .A3(new_n632_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n732_), .A2(new_n733_), .ZN(G1333gat));
  INV_X1    g533(.A(G71gat), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n726_), .A2(new_n735_), .A3(new_n645_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n728_), .A2(new_n645_), .ZN(new_n737_));
  XOR2_X1   g536(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(G71gat), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n737_), .B2(G71gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  XOR2_X1   g540(.A(new_n741_), .B(KEYINPUT109), .Z(G1334gat));
  INV_X1    g541(.A(G78gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n728_), .B2(new_n427_), .ZN(new_n744_));
  XOR2_X1   g543(.A(new_n744_), .B(KEYINPUT50), .Z(new_n745_));
  NOR2_X1   g544(.A1(new_n290_), .A2(G78gat), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT110), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n726_), .A2(new_n747_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n745_), .A2(new_n748_), .ZN(G1335gat));
  NAND4_X1  g548(.A1(new_n670_), .A2(new_n466_), .A3(new_n724_), .A4(new_n657_), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n750_), .B(KEYINPUT111), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n619_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n625_), .A2(new_n626_), .A3(new_n656_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n755_), .B1(new_n686_), .B2(new_n691_), .ZN(new_n756_));
  XOR2_X1   g555(.A(new_n756_), .B(KEYINPUT112), .Z(new_n757_));
  AND2_X1   g556(.A1(new_n619_), .A2(G85gat), .ZN(new_n758_));
  AOI21_X1  g557(.A(new_n753_), .B1(new_n757_), .B2(new_n758_), .ZN(G1336gat));
  AOI21_X1  g558(.A(G92gat), .B1(new_n752_), .B2(new_n632_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n632_), .A2(G92gat), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n757_), .B2(new_n761_), .ZN(G1337gat));
  INV_X1    g561(.A(new_n756_), .ZN(new_n763_));
  OAI21_X1  g562(.A(G99gat), .B1(new_n763_), .B2(new_n429_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n397_), .A2(new_n484_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n751_), .B2(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n766_), .B(KEYINPUT51), .ZN(G1338gat));
  OR3_X1    g566(.A1(new_n751_), .A2(new_n290_), .A3(new_n485_), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT52), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n700_), .A2(new_n290_), .A3(new_n755_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n479_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(KEYINPUT104), .B1(new_n687_), .B2(new_n542_), .ZN(new_n773_));
  AOI211_X1 g572(.A(new_n677_), .B(new_n541_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n688_), .B1(new_n775_), .B2(new_n670_), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n427_), .B(new_n754_), .C1(new_n776_), .C2(new_n690_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT113), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n769_), .B1(new_n772_), .B2(new_n778_), .ZN(new_n779_));
  OAI21_X1  g578(.A(G106gat), .B1(new_n777_), .B2(KEYINPUT113), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n771_), .B1(new_n756_), .B2(new_n427_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(KEYINPUT52), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n768_), .B1(new_n779_), .B2(new_n782_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n783_), .A2(KEYINPUT53), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT53), .ZN(new_n785_));
  OAI211_X1 g584(.A(new_n785_), .B(new_n768_), .C1(new_n779_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n784_), .A2(new_n786_), .ZN(G1339gat));
  INV_X1    g586(.A(KEYINPUT118), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n553_), .A2(new_n466_), .A3(new_n615_), .ZN(new_n789_));
  XNOR2_X1  g588(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n790_));
  INV_X1    g589(.A(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n789_), .A2(new_n791_), .ZN(new_n792_));
  NAND4_X1  g591(.A1(new_n553_), .A2(new_n466_), .A3(new_n615_), .A4(new_n790_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n608_), .ZN(new_n795_));
  NOR3_X1   g594(.A1(new_n594_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n596_), .B1(new_n594_), .B2(new_n597_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n796_), .B1(KEYINPUT55), .B2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  NOR4_X1   g598(.A1(new_n594_), .A2(new_n597_), .A3(new_n799_), .A4(new_n596_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n795_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT56), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n797_), .A2(KEYINPUT55), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n598_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n800_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n807_), .A2(KEYINPUT56), .A3(new_n795_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n803_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n446_), .A2(new_n449_), .A3(new_n452_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n450_), .B1(new_n448_), .B2(new_n453_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n810_), .A2(new_n459_), .A3(new_n811_), .ZN(new_n812_));
  AND3_X1   g611(.A1(new_n609_), .A2(new_n461_), .A3(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n809_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT58), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n809_), .A2(KEYINPUT58), .A3(new_n813_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n816_), .A2(new_n683_), .A3(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n466_), .A2(new_n610_), .ZN(new_n819_));
  AOI21_X1  g618(.A(KEYINPUT56), .B1(new_n807_), .B2(new_n795_), .ZN(new_n820_));
  AOI211_X1 g619(.A(new_n802_), .B(new_n608_), .C1(new_n805_), .C2(new_n806_), .ZN(new_n821_));
  OAI21_X1  g620(.A(new_n819_), .B1(new_n820_), .B2(new_n821_), .ZN(new_n822_));
  OAI211_X1 g621(.A(new_n461_), .B(new_n812_), .C1(new_n610_), .C2(new_n611_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n546_), .B1(new_n822_), .B2(new_n823_), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n824_), .A2(KEYINPUT57), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n826_));
  INV_X1    g625(.A(new_n823_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n827_), .B1(new_n809_), .B2(new_n819_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n826_), .B1(new_n828_), .B2(new_n546_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n818_), .A2(new_n825_), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(new_n794_), .B1(new_n830_), .B2(new_n591_), .ZN(new_n831_));
  INV_X1    g630(.A(new_n361_), .ZN(new_n832_));
  NOR2_X1   g631(.A1(new_n386_), .A2(new_n397_), .ZN(new_n833_));
  XOR2_X1   g632(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n833_), .A3(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n831_), .A2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(G113gat), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n466_), .A2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n824_), .B2(KEYINPUT57), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT115), .B(new_n826_), .C1(new_n828_), .C2(new_n546_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n841_), .A2(new_n842_), .A3(new_n825_), .A4(new_n818_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n794_), .B1(new_n843_), .B2(new_n591_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n832_), .A2(new_n833_), .ZN(new_n845_));
  OAI21_X1  g644(.A(KEYINPUT59), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(KEYINPUT116), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT116), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n848_), .B(KEYINPUT59), .C1(new_n844_), .C2(new_n845_), .ZN(new_n849_));
  AOI211_X1 g648(.A(new_n836_), .B(new_n839_), .C1(new_n847_), .C2(new_n849_), .ZN(new_n850_));
  NOR2_X1   g649(.A1(new_n844_), .A2(new_n845_), .ZN(new_n851_));
  AOI21_X1  g650(.A(G113gat), .B1(new_n851_), .B2(new_n626_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n788_), .B1(new_n850_), .B2(new_n852_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n847_), .A2(new_n849_), .ZN(new_n854_));
  INV_X1    g653(.A(new_n836_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n854_), .A2(new_n855_), .A3(new_n838_), .ZN(new_n856_));
  INV_X1    g655(.A(new_n852_), .ZN(new_n857_));
  NAND3_X1  g656(.A1(new_n856_), .A2(KEYINPUT118), .A3(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n853_), .A2(new_n858_), .ZN(G1340gat));
  INV_X1    g658(.A(G120gat), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n860_), .B1(new_n625_), .B2(KEYINPUT60), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n851_), .B(new_n861_), .C1(KEYINPUT60), .C2(new_n860_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n724_), .B1(new_n831_), .B2(new_n835_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n863_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n864_));
  AND2_X1   g663(.A1(new_n864_), .A2(KEYINPUT119), .ZN(new_n865_));
  OAI21_X1  g664(.A(G120gat), .B1(new_n864_), .B2(KEYINPUT119), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n862_), .B1(new_n865_), .B2(new_n866_), .ZN(G1341gat));
  AOI21_X1  g666(.A(G127gat), .B1(new_n851_), .B2(new_n656_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n836_), .B1(new_n847_), .B2(new_n849_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n656_), .A2(G127gat), .ZN(new_n870_));
  XOR2_X1   g669(.A(new_n870_), .B(KEYINPUT120), .Z(new_n871_));
  AOI21_X1  g670(.A(new_n868_), .B1(new_n869_), .B2(new_n871_), .ZN(G1342gat));
  INV_X1    g671(.A(G134gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n851_), .A2(new_n873_), .A3(new_n546_), .ZN(new_n874_));
  AND2_X1   g673(.A1(new_n869_), .A2(new_n683_), .ZN(new_n875_));
  OAI21_X1  g674(.A(new_n874_), .B1(new_n875_), .B2(new_n873_), .ZN(G1343gat));
  NAND3_X1  g675(.A1(new_n429_), .A2(new_n619_), .A3(new_n360_), .ZN(new_n877_));
  NOR3_X1   g676(.A1(new_n844_), .A2(new_n290_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n626_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n724_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g681(.A(KEYINPUT61), .B(G155gat), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n878_), .A2(new_n656_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(KEYINPUT121), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n885_), .A2(KEYINPUT121), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n884_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n888_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n890_), .A2(new_n886_), .A3(new_n883_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(G1346gat));
  AOI21_X1  g691(.A(G162gat), .B1(new_n878_), .B2(new_n546_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n775_), .A2(G162gat), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n878_), .B2(new_n894_), .ZN(G1347gat));
  NOR2_X1   g694(.A1(new_n831_), .A2(new_n427_), .ZN(new_n896_));
  NOR3_X1   g695(.A1(new_n429_), .A2(new_n619_), .A3(new_n360_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n898_), .A2(new_n466_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n896_), .A2(new_n302_), .A3(new_n899_), .ZN(new_n900_));
  INV_X1    g699(.A(G169gat), .ZN(new_n901_));
  XOR2_X1   g700(.A(new_n899_), .B(KEYINPUT122), .Z(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n896_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904_));
  AND2_X1   g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n904_), .ZN(new_n906_));
  OAI21_X1  g705(.A(new_n900_), .B1(new_n905_), .B2(new_n906_), .ZN(G1348gat));
  NAND2_X1  g706(.A1(new_n896_), .A2(new_n897_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n724_), .A2(new_n303_), .ZN(new_n909_));
  NOR4_X1   g708(.A1(new_n844_), .A2(new_n427_), .A3(new_n625_), .A4(new_n898_), .ZN(new_n910_));
  OAI22_X1  g709(.A1(new_n908_), .A2(new_n909_), .B1(new_n910_), .B2(new_n303_), .ZN(G1349gat));
  NOR2_X1   g710(.A1(new_n898_), .A2(new_n591_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n896_), .A2(new_n318_), .A3(new_n912_), .ZN(new_n913_));
  AND2_X1   g712(.A1(new_n913_), .A2(KEYINPUT123), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n913_), .A2(KEYINPUT123), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n844_), .A2(new_n427_), .ZN(new_n916_));
  AOI21_X1  g715(.A(G183gat), .B1(new_n916_), .B2(new_n912_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n914_), .A2(new_n915_), .A3(new_n917_), .ZN(G1350gat));
  OAI21_X1  g717(.A(G190gat), .B1(new_n908_), .B2(new_n553_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n546_), .A2(new_n319_), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n908_), .B2(new_n920_), .ZN(G1351gat));
  NAND4_X1  g720(.A1(new_n427_), .A2(new_n386_), .A3(new_n632_), .A4(new_n429_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(new_n844_), .A2(new_n922_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n626_), .ZN(new_n924_));
  XNOR2_X1  g723(.A(new_n924_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g724(.A1(new_n923_), .A2(new_n724_), .ZN(new_n926_));
  MUX2_X1   g725(.A(new_n259_), .B(G204gat), .S(new_n926_), .Z(G1353gat));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(KEYINPUT124), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(KEYINPUT125), .ZN(new_n930_));
  NAND2_X1  g729(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n931_));
  NAND4_X1  g730(.A1(new_n923_), .A2(new_n656_), .A3(new_n930_), .A4(new_n931_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n929_), .A2(KEYINPUT125), .ZN(new_n933_));
  XNOR2_X1  g732(.A(new_n932_), .B(new_n933_), .ZN(G1354gat));
  NAND2_X1  g733(.A1(new_n923_), .A2(new_n546_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT126), .ZN(new_n936_));
  XOR2_X1   g735(.A(KEYINPUT127), .B(G218gat), .Z(new_n937_));
  NOR2_X1   g736(.A1(new_n553_), .A2(new_n937_), .ZN(new_n938_));
  AOI22_X1  g737(.A1(new_n936_), .A2(new_n937_), .B1(new_n923_), .B2(new_n938_), .ZN(G1355gat));
endmodule


