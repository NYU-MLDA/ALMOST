//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n750_, new_n751_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n786_, new_n787_, new_n789_, new_n790_, new_n791_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n797_, new_n798_,
    new_n799_, new_n800_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n810_,
    new_n811_, new_n812_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n901_, new_n902_, new_n903_, new_n904_, new_n905_,
    new_n906_, new_n907_, new_n909_, new_n911_, new_n912_, new_n914_,
    new_n915_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n940_, new_n941_,
    new_n943_, new_n944_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n957_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n972_, new_n973_, new_n974_, new_n975_;
  INV_X1    g000(.A(G169gat), .ZN(new_n202_));
  OAI21_X1  g001(.A(KEYINPUT22), .B1(new_n202_), .B2(KEYINPUT81), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT81), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT22), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(G169gat), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G169gat), .A2(G176gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  INV_X1    g009(.A(G183gat), .ZN(new_n211_));
  INV_X1    g010(.A(G190gat), .ZN(new_n212_));
  OAI21_X1  g011(.A(KEYINPUT23), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT82), .ZN(new_n214_));
  NOR2_X1   g013(.A1(new_n211_), .A2(KEYINPUT23), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n214_), .B1(new_n215_), .B2(G190gat), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT23), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n214_), .A2(new_n217_), .A3(G183gat), .A4(G190gat), .ZN(new_n218_));
  INV_X1    g017(.A(new_n218_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n213_), .B1(new_n216_), .B2(new_n219_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G183gat), .A2(G190gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n210_), .B1(new_n220_), .B2(new_n222_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n224_));
  AND2_X1   g023(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n225_));
  AND2_X1   g024(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n227_));
  OAI22_X1  g026(.A1(new_n224_), .A2(new_n225_), .B1(new_n226_), .B2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n217_), .A2(G183gat), .A3(G190gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n213_), .A2(new_n229_), .ZN(new_n230_));
  NOR3_X1   g029(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n231_));
  INV_X1    g030(.A(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n228_), .A2(new_n230_), .A3(new_n232_), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT80), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n209_), .A2(KEYINPUT24), .ZN(new_n235_));
  NOR2_X1   g034(.A1(G169gat), .A2(G176gat), .ZN(new_n236_));
  OAI21_X1  g035(.A(new_n234_), .B1(new_n235_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n202_), .A2(new_n207_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n238_), .A2(KEYINPUT80), .A3(KEYINPUT24), .A4(new_n209_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NOR2_X1   g039(.A1(new_n233_), .A2(new_n240_), .ZN(new_n241_));
  OAI21_X1  g040(.A(KEYINPUT83), .B1(new_n223_), .B2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n209_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n204_), .A2(G169gat), .ZN(new_n244_));
  AOI21_X1  g043(.A(G176gat), .B1(new_n244_), .B2(KEYINPUT22), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n245_), .B2(new_n206_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n217_), .B1(G183gat), .B2(G190gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n229_), .A2(KEYINPUT82), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n247_), .B1(new_n248_), .B2(new_n218_), .ZN(new_n249_));
  OAI21_X1  g048(.A(new_n246_), .B1(new_n249_), .B2(new_n221_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT25), .B(G183gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(KEYINPUT26), .B(G190gat), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n231_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n253_), .A2(new_n230_), .A3(new_n239_), .A4(new_n237_), .ZN(new_n254_));
  INV_X1    g053(.A(KEYINPUT83), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n250_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n242_), .A2(new_n256_), .ZN(new_n257_));
  XNOR2_X1  g056(.A(G71gat), .B(G99gat), .ZN(new_n258_));
  INV_X1    g057(.A(G43gat), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n257_), .B(new_n260_), .ZN(new_n261_));
  OR2_X1    g060(.A1(G113gat), .A2(G120gat), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT84), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G113gat), .A2(G120gat), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n262_), .A2(new_n263_), .A3(new_n264_), .ZN(new_n265_));
  AND2_X1   g064(.A1(G113gat), .A2(G120gat), .ZN(new_n266_));
  NOR2_X1   g065(.A1(G113gat), .A2(G120gat), .ZN(new_n267_));
  OAI21_X1  g066(.A(KEYINPUT84), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n265_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G127gat), .B(G134gat), .ZN(new_n270_));
  INV_X1    g069(.A(new_n270_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n265_), .A2(new_n268_), .A3(new_n270_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n272_), .A2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(G227gat), .A2(G233gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT30), .B(G15gat), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n277_), .B(KEYINPUT31), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n276_), .B(new_n278_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n261_), .A2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n261_), .A2(new_n279_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n282_), .ZN(new_n283_));
  XNOR2_X1  g082(.A(G197gat), .B(G204gat), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT21), .ZN(new_n285_));
  NOR2_X1   g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(G211gat), .B(G218gat), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n286_), .A2(new_n288_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n284_), .A2(new_n285_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n287_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n289_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT85), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT85), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n296_), .A2(G155gat), .A3(G162gat), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n295_), .A2(new_n297_), .ZN(new_n298_));
  NOR2_X1   g097(.A1(G155gat), .A2(G162gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n298_), .A2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT86), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  AOI21_X1  g102(.A(new_n299_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT86), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT3), .ZN(new_n306_));
  INV_X1    g105(.A(G141gat), .ZN(new_n307_));
  INV_X1    g106(.A(G148gat), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n306_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  NAND2_X1  g108(.A1(G141gat), .A2(G148gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT2), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n310_), .A2(new_n311_), .ZN(new_n312_));
  OAI21_X1  g111(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n314_));
  NAND4_X1  g113(.A1(new_n309_), .A2(new_n312_), .A3(new_n313_), .A4(new_n314_), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n303_), .A2(new_n305_), .A3(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n298_), .A2(KEYINPUT1), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT1), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n295_), .A2(new_n297_), .A3(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n317_), .A2(new_n300_), .A3(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n310_), .ZN(new_n321_));
  NOR2_X1   g120(.A1(G141gat), .A2(G148gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n320_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n316_), .A2(new_n324_), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n293_), .B1(new_n325_), .B2(KEYINPUT29), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G228gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT28), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G22gat), .B(G50gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n326_), .B(new_n330_), .ZN(new_n331_));
  NOR2_X1   g130(.A1(new_n325_), .A2(KEYINPUT29), .ZN(new_n332_));
  XOR2_X1   g131(.A(G78gat), .B(G106gat), .Z(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  OR2_X1    g133(.A1(new_n331_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n331_), .A2(new_n334_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G8gat), .B(G36gat), .ZN(new_n339_));
  INV_X1    g138(.A(G92gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT18), .B(G64gat), .ZN(new_n342_));
  XOR2_X1   g141(.A(new_n341_), .B(new_n342_), .Z(new_n343_));
  NAND2_X1  g142(.A1(G226gat), .A2(G233gat), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT19), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT20), .ZN(new_n346_));
  NOR2_X1   g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n230_), .A2(new_n222_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n205_), .A2(G169gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n202_), .A2(KEYINPUT22), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n349_), .A2(new_n350_), .A3(new_n207_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n209_), .A2(KEYINPUT88), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT88), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n354_), .A2(G169gat), .A3(G176gat), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n352_), .A2(KEYINPUT89), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT89), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n353_), .A2(new_n355_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n358_), .B1(new_n359_), .B2(new_n351_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n348_), .B1(new_n357_), .B2(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n238_), .A2(KEYINPUT24), .A3(new_n209_), .ZN(new_n362_));
  AND3_X1   g161(.A1(new_n228_), .A2(new_n232_), .A3(new_n362_), .ZN(new_n363_));
  AOI21_X1  g162(.A(KEYINPUT87), .B1(new_n363_), .B2(new_n220_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n228_), .A2(new_n232_), .A3(new_n362_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT87), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n365_), .A2(new_n249_), .A3(new_n366_), .ZN(new_n367_));
  OAI21_X1  g166(.A(new_n361_), .B1(new_n364_), .B2(new_n367_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n347_), .B1(new_n368_), .B2(new_n292_), .ZN(new_n369_));
  AND3_X1   g168(.A1(new_n250_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n255_), .B1(new_n250_), .B2(new_n254_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n292_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT90), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n257_), .A2(KEYINPUT90), .A3(new_n292_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n369_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n345_), .ZN(new_n377_));
  AOI21_X1  g176(.A(new_n346_), .B1(new_n368_), .B2(new_n292_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n242_), .A2(new_n293_), .A3(new_n256_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n377_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n343_), .B1(new_n376_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n369_), .ZN(new_n382_));
  AOI21_X1  g181(.A(KEYINPUT90), .B1(new_n257_), .B2(new_n292_), .ZN(new_n383_));
  AOI211_X1 g182(.A(new_n373_), .B(new_n293_), .C1(new_n242_), .C2(new_n256_), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n382_), .B1(new_n383_), .B2(new_n384_), .ZN(new_n385_));
  INV_X1    g184(.A(new_n343_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n379_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n366_), .B1(new_n365_), .B2(new_n249_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n363_), .A2(KEYINPUT87), .A3(new_n220_), .ZN(new_n389_));
  OAI21_X1  g188(.A(KEYINPUT89), .B1(new_n352_), .B2(new_n356_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n359_), .A2(new_n358_), .A3(new_n351_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n390_), .A2(new_n391_), .ZN(new_n392_));
  AOI22_X1  g191(.A1(new_n388_), .A2(new_n389_), .B1(new_n392_), .B2(new_n348_), .ZN(new_n393_));
  OAI21_X1  g192(.A(KEYINPUT20), .B1(new_n393_), .B2(new_n293_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n345_), .B1(new_n387_), .B2(new_n394_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n385_), .A2(new_n386_), .A3(new_n395_), .ZN(new_n396_));
  AND2_X1   g195(.A1(new_n381_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT91), .ZN(new_n398_));
  INV_X1    g197(.A(new_n273_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n270_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n315_), .B1(new_n304_), .B2(KEYINPUT86), .ZN(new_n402_));
  AOI211_X1 g201(.A(new_n302_), .B(new_n299_), .C1(new_n295_), .C2(new_n297_), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(new_n323_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n299_), .B1(new_n298_), .B2(KEYINPUT1), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n405_), .B1(new_n406_), .B2(new_n319_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n401_), .B1(new_n404_), .B2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n316_), .A2(new_n324_), .A3(new_n274_), .ZN(new_n409_));
  AND3_X1   g208(.A1(new_n408_), .A2(new_n409_), .A3(KEYINPUT4), .ZN(new_n410_));
  NAND2_X1  g209(.A1(G225gat), .A2(G233gat), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n412_), .B1(new_n408_), .B2(KEYINPUT4), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n398_), .B1(new_n410_), .B2(new_n413_), .ZN(new_n414_));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415_));
  INV_X1    g214(.A(G85gat), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n415_), .B(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT0), .B(G57gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n417_), .B(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n408_), .A2(new_n409_), .A3(KEYINPUT4), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT4), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n325_), .A2(new_n421_), .A3(new_n401_), .ZN(new_n422_));
  NAND4_X1  g221(.A1(new_n420_), .A2(KEYINPUT91), .A3(new_n412_), .A4(new_n422_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n408_), .A2(new_n409_), .A3(new_n411_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n414_), .A2(new_n419_), .A3(new_n423_), .A4(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n425_), .A2(KEYINPUT92), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n426_), .A2(KEYINPUT33), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT33), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n425_), .A2(KEYINPUT92), .A3(new_n428_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n420_), .A2(new_n411_), .A3(new_n422_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n419_), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n408_), .A2(new_n409_), .A3(new_n412_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n397_), .A2(new_n427_), .A3(new_n429_), .A4(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n414_), .A2(new_n423_), .A3(new_n424_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n435_), .A2(new_n431_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n425_), .ZN(new_n437_));
  NOR2_X1   g236(.A1(new_n376_), .A2(new_n380_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n386_), .A2(KEYINPUT32), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n378_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT95), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT95), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n378_), .A2(new_n443_), .A3(new_n377_), .A4(new_n379_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n442_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n374_), .A2(new_n375_), .ZN(new_n446_));
  XNOR2_X1  g245(.A(KEYINPUT93), .B(KEYINPUT20), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n363_), .A2(new_n220_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n361_), .A2(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n292_), .B1(new_n449_), .B2(KEYINPUT94), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT94), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n361_), .A2(new_n451_), .A3(new_n448_), .ZN(new_n452_));
  AOI21_X1  g251(.A(new_n447_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n377_), .B1(new_n446_), .B2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n445_), .A2(new_n454_), .ZN(new_n455_));
  OAI211_X1 g254(.A(new_n437_), .B(new_n440_), .C1(new_n455_), .C2(new_n439_), .ZN(new_n456_));
  AOI21_X1  g255(.A(new_n338_), .B1(new_n434_), .B2(new_n456_), .ZN(new_n457_));
  NOR2_X1   g256(.A1(new_n437_), .A2(new_n337_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n343_), .B1(new_n445_), .B2(new_n454_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT27), .ZN(new_n460_));
  AOI21_X1  g259(.A(new_n460_), .B1(new_n438_), .B2(new_n386_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n459_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n381_), .A2(new_n396_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n460_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n458_), .A2(new_n462_), .A3(new_n464_), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n283_), .B1(new_n457_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n462_), .A2(new_n464_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n282_), .A2(new_n337_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(new_n437_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n466_), .A2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G230gat), .A2(G233gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n473_), .B(KEYINPUT64), .ZN(new_n474_));
  INV_X1    g273(.A(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT7), .ZN(new_n476_));
  INV_X1    g275(.A(G99gat), .ZN(new_n477_));
  INV_X1    g276(.A(G106gat), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n476_), .A2(new_n477_), .A3(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n484_));
  NAND4_X1  g283(.A1(new_n479_), .A2(new_n482_), .A3(new_n483_), .A4(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n340_), .A2(G85gat), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n416_), .A2(G92gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n485_), .A2(new_n488_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT8), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n485_), .A2(KEYINPUT8), .A3(new_n488_), .ZN(new_n492_));
  AND2_X1   g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n482_), .A2(new_n483_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n494_), .B1(KEYINPUT9), .B2(new_n488_), .ZN(new_n495_));
  NOR2_X1   g294(.A1(new_n416_), .A2(KEYINPUT9), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n340_), .A2(KEYINPUT66), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT66), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(G92gat), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(KEYINPUT10), .B(G99gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT65), .B1(new_n501_), .B2(G106gat), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT65), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n477_), .A2(KEYINPUT10), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n477_), .A2(KEYINPUT10), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n503_), .B(new_n478_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n495_), .A2(new_n500_), .A3(new_n502_), .A4(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(G71gat), .B(G78gat), .Z(new_n508_));
  INV_X1    g307(.A(G57gat), .ZN(new_n509_));
  INV_X1    g308(.A(G64gat), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT11), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G57gat), .A2(G64gat), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n508_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT67), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n511_), .A2(new_n513_), .ZN(new_n517_));
  INV_X1    g316(.A(KEYINPUT67), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n508_), .A2(new_n514_), .A3(new_n518_), .ZN(new_n519_));
  NAND4_X1  g318(.A1(new_n516_), .A2(KEYINPUT11), .A3(new_n517_), .A4(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(KEYINPUT11), .ZN(new_n521_));
  AND3_X1   g320(.A1(new_n508_), .A2(new_n514_), .A3(new_n518_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n518_), .B1(new_n508_), .B2(new_n514_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n521_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  NAND4_X1  g323(.A1(new_n493_), .A2(new_n507_), .A3(new_n520_), .A4(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n520_), .A2(new_n524_), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n507_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n525_), .A2(new_n528_), .A3(KEYINPUT12), .ZN(new_n529_));
  INV_X1    g328(.A(KEYINPUT12), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n526_), .A2(new_n527_), .A3(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n475_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT68), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n525_), .A2(new_n528_), .A3(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n526_), .A2(new_n527_), .A3(KEYINPUT68), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n535_), .A2(new_n475_), .A3(new_n536_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n533_), .A2(new_n537_), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G120gat), .B(G148gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT70), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(KEYINPUT69), .ZN(new_n541_));
  XOR2_X1   g340(.A(G176gat), .B(G204gat), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n542_), .B(KEYINPUT5), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n541_), .B(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n538_), .A2(new_n545_), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n533_), .A2(new_n537_), .A3(new_n544_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT13), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n546_), .A2(KEYINPUT13), .A3(new_n547_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n550_), .A2(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G15gat), .B(G22gat), .ZN(new_n553_));
  INV_X1    g352(.A(G1gat), .ZN(new_n554_));
  INV_X1    g353(.A(G8gat), .ZN(new_n555_));
  OAI21_X1  g354(.A(KEYINPUT14), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n553_), .A2(new_n556_), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G1gat), .B(G8gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n557_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(G36gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(G29gat), .ZN(new_n561_));
  INV_X1    g360(.A(G29gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(G36gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n561_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(G50gat), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(G43gat), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n259_), .A2(G50gat), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT71), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n568_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n564_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n259_), .A2(G50gat), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n565_), .A2(G43gat), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT71), .B1(new_n572_), .B2(new_n573_), .ZN(new_n574_));
  NAND3_X1  g373(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n575_));
  AND2_X1   g374(.A1(new_n561_), .A2(new_n563_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n571_), .A2(new_n577_), .ZN(new_n578_));
  AND2_X1   g377(.A1(new_n559_), .A2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n559_), .A2(new_n578_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G229gat), .A2(G233gat), .ZN(new_n582_));
  NOR2_X1   g381(.A1(new_n581_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(KEYINPUT72), .B(KEYINPUT15), .Z(new_n585_));
  NAND3_X1  g384(.A1(new_n571_), .A2(new_n577_), .A3(new_n585_), .ZN(new_n586_));
  OAI211_X1 g385(.A(new_n586_), .B(new_n582_), .C1(new_n581_), .C2(new_n585_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n584_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(G113gat), .B(G141gat), .ZN(new_n589_));
  XNOR2_X1  g388(.A(G169gat), .B(G197gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n589_), .B(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n591_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n588_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n584_), .A2(new_n587_), .A3(new_n591_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n593_), .A2(new_n594_), .A3(KEYINPUT79), .ZN(new_n595_));
  OR3_X1    g394(.A1(new_n588_), .A2(KEYINPUT79), .A3(new_n592_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n552_), .A2(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(new_n472_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n585_), .ZN(new_n600_));
  NOR3_X1   g399(.A1(new_n569_), .A2(new_n570_), .A3(new_n564_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n576_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n600_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n491_), .A2(new_n492_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n502_), .A2(new_n506_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n488_), .A2(KEYINPUT9), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n482_), .A2(new_n483_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n606_), .A2(new_n607_), .A3(new_n500_), .ZN(new_n608_));
  NOR2_X1   g407(.A1(new_n605_), .A2(new_n608_), .ZN(new_n609_));
  OAI211_X1 g408(.A(new_n603_), .B(new_n586_), .C1(new_n604_), .C2(new_n609_), .ZN(new_n610_));
  NAND4_X1  g409(.A1(new_n507_), .A2(new_n578_), .A3(new_n491_), .A4(new_n492_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n612_), .A2(KEYINPUT35), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n610_), .A2(KEYINPUT73), .A3(new_n611_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT34), .ZN(new_n615_));
  INV_X1    g414(.A(G232gat), .ZN(new_n616_));
  INV_X1    g415(.A(G233gat), .ZN(new_n617_));
  NOR2_X1   g416(.A1(new_n616_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT34), .ZN(new_n620_));
  NAND4_X1  g419(.A1(new_n610_), .A2(KEYINPUT73), .A3(new_n620_), .A4(new_n611_), .ZN(new_n621_));
  AND3_X1   g420(.A1(new_n615_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n619_), .B1(new_n615_), .B2(new_n621_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n613_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n615_), .A2(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n625_), .A2(new_n618_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n615_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n627_));
  NAND3_X1  g426(.A1(new_n626_), .A2(KEYINPUT35), .A3(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n624_), .A2(new_n628_), .A3(KEYINPUT75), .ZN(new_n629_));
  XOR2_X1   g428(.A(G134gat), .B(G162gat), .Z(new_n630_));
  XNOR2_X1  g429(.A(new_n630_), .B(KEYINPUT74), .ZN(new_n631_));
  XOR2_X1   g430(.A(G190gat), .B(G218gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(new_n631_), .B(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT36), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n633_), .A2(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n624_), .A2(new_n628_), .ZN(new_n637_));
  NOR2_X1   g436(.A1(new_n633_), .A2(new_n634_), .ZN(new_n638_));
  AOI22_X1  g437(.A1(new_n629_), .A2(new_n636_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n624_), .A2(new_n628_), .A3(KEYINPUT75), .A4(new_n635_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT37), .B1(new_n639_), .B2(new_n640_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n629_), .A2(new_n636_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n637_), .A2(new_n638_), .ZN(new_n643_));
  AND4_X1   g442(.A1(KEYINPUT37), .A2(new_n642_), .A3(new_n640_), .A4(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n641_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(G231gat), .A2(G233gat), .ZN(new_n646_));
  XNOR2_X1  g445(.A(new_n559_), .B(new_n646_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(new_n526_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(G127gat), .B(G155gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(G211gat), .ZN(new_n650_));
  XNOR2_X1  g449(.A(KEYINPUT16), .B(G183gat), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n650_), .B(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(KEYINPUT78), .B(KEYINPUT17), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n652_), .B(new_n653_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n648_), .A2(new_n654_), .ZN(new_n655_));
  XOR2_X1   g454(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n656_));
  NAND2_X1  g455(.A1(new_n652_), .A2(new_n656_), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT77), .Z(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(new_n648_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n655_), .A2(new_n659_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n645_), .A2(new_n660_), .ZN(new_n661_));
  AND2_X1   g460(.A1(new_n599_), .A2(new_n661_), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n554_), .A3(new_n437_), .ZN(new_n663_));
  XNOR2_X1  g462(.A(new_n663_), .B(KEYINPUT38), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n642_), .A2(new_n640_), .A3(new_n643_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n472_), .A2(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n660_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n598_), .A2(new_n670_), .ZN(new_n671_));
  XNOR2_X1  g470(.A(new_n671_), .B(KEYINPUT96), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n669_), .A2(new_n672_), .ZN(new_n673_));
  OAI21_X1  g472(.A(G1gat), .B1(new_n673_), .B2(new_n470_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n664_), .A2(new_n674_), .ZN(G1324gat));
  NAND3_X1  g474(.A1(new_n662_), .A2(new_n555_), .A3(new_n467_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT98), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n667_), .A2(new_n668_), .ZN(new_n678_));
  AOI21_X1  g477(.A(KEYINPUT97), .B1(new_n472_), .B2(new_n666_), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n467_), .B(new_n672_), .C1(new_n678_), .C2(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT99), .ZN(new_n681_));
  OR2_X1    g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT39), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n555_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n684_));
  AND3_X1   g483(.A1(new_n682_), .A2(new_n683_), .A3(new_n684_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n683_), .B1(new_n682_), .B2(new_n684_), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n677_), .B1(new_n685_), .B2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT40), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT40), .B(new_n677_), .C1(new_n685_), .C2(new_n686_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(G1325gat));
  OAI21_X1  g490(.A(G15gat), .B1(new_n673_), .B2(new_n283_), .ZN(new_n692_));
  XOR2_X1   g491(.A(KEYINPUT100), .B(KEYINPUT41), .Z(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(new_n662_), .ZN(new_n695_));
  OR2_X1    g494(.A1(new_n283_), .A2(G15gat), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(G1326gat));
  OAI21_X1  g496(.A(G22gat), .B1(new_n673_), .B2(new_n337_), .ZN(new_n698_));
  XOR2_X1   g497(.A(KEYINPUT101), .B(KEYINPUT42), .Z(new_n699_));
  OR2_X1    g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n698_), .A2(new_n699_), .ZN(new_n701_));
  OR3_X1    g500(.A1(new_n695_), .A2(G22gat), .A3(new_n337_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n700_), .A2(new_n701_), .A3(new_n702_), .ZN(G1327gat));
  NOR2_X1   g502(.A1(new_n666_), .A2(new_n670_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n599_), .A2(new_n704_), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n705_), .B(KEYINPUT104), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(new_n562_), .A3(new_n437_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT37), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n665_), .A2(new_n709_), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n639_), .A2(KEYINPUT37), .A3(new_n640_), .ZN(new_n711_));
  NAND2_X1  g510(.A1(new_n710_), .A2(new_n711_), .ZN(new_n712_));
  AOI21_X1  g511(.A(new_n712_), .B1(new_n466_), .B2(new_n471_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT102), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n708_), .B1(new_n713_), .B2(new_n714_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n472_), .A2(new_n645_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n716_), .A2(KEYINPUT102), .A3(KEYINPUT43), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n715_), .A2(new_n717_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n552_), .A2(new_n597_), .A3(new_n670_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT44), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(KEYINPUT103), .A3(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n721_), .A2(KEYINPUT103), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n718_), .A2(new_n723_), .A3(new_n719_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n722_), .A2(new_n437_), .A3(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n707_), .B1(new_n725_), .B2(new_n562_), .ZN(G1328gat));
  INV_X1    g525(.A(new_n467_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n727_), .A2(G36gat), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n706_), .A2(new_n728_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(KEYINPUT45), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n731_));
  NAND3_X1  g530(.A1(new_n706_), .A2(new_n731_), .A3(new_n728_), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n730_), .A2(new_n732_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n722_), .A2(new_n467_), .A3(new_n724_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n734_), .A2(G36gat), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n733_), .A2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT46), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  NAND3_X1  g537(.A1(new_n733_), .A2(new_n735_), .A3(KEYINPUT46), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(G1329gat));
  NAND3_X1  g539(.A1(new_n722_), .A2(new_n282_), .A3(new_n724_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(G43gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n706_), .A2(new_n259_), .A3(new_n282_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n745_));
  INV_X1    g544(.A(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n744_), .A2(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n742_), .A2(new_n743_), .A3(new_n745_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1330gat));
  NAND3_X1  g548(.A1(new_n706_), .A2(new_n565_), .A3(new_n338_), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n722_), .A2(new_n338_), .A3(new_n724_), .ZN(new_n751_));
  OAI21_X1  g550(.A(new_n750_), .B1(new_n751_), .B2(new_n565_), .ZN(G1331gat));
  AND2_X1   g551(.A1(new_n550_), .A2(new_n551_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n597_), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(new_n754_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(new_n756_), .B1(new_n466_), .B2(new_n471_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n757_), .A2(new_n661_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(G57gat), .B1(new_n759_), .B2(new_n437_), .ZN(new_n760_));
  AND3_X1   g559(.A1(new_n669_), .A2(new_n670_), .A3(new_n755_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n470_), .A2(new_n509_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(G1332gat));
  AOI21_X1  g562(.A(new_n510_), .B1(new_n761_), .B2(new_n467_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT48), .Z(new_n765_));
  NAND3_X1  g564(.A1(new_n759_), .A2(new_n510_), .A3(new_n467_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(G1333gat));
  INV_X1    g566(.A(G71gat), .ZN(new_n768_));
  AOI21_X1  g567(.A(new_n768_), .B1(new_n761_), .B2(new_n282_), .ZN(new_n769_));
  XOR2_X1   g568(.A(new_n769_), .B(KEYINPUT49), .Z(new_n770_));
  NAND2_X1  g569(.A1(new_n282_), .A2(new_n768_), .ZN(new_n771_));
  XOR2_X1   g570(.A(new_n771_), .B(KEYINPUT106), .Z(new_n772_));
  OAI21_X1  g571(.A(new_n770_), .B1(new_n758_), .B2(new_n772_), .ZN(G1334gat));
  NAND2_X1  g572(.A1(new_n761_), .A2(new_n338_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n774_), .A2(G78gat), .ZN(new_n775_));
  XNOR2_X1  g574(.A(new_n775_), .B(KEYINPUT50), .ZN(new_n776_));
  OR2_X1    g575(.A1(new_n337_), .A2(G78gat), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n776_), .B1(new_n758_), .B2(new_n777_), .ZN(G1335gat));
  NAND2_X1  g577(.A1(new_n757_), .A2(new_n704_), .ZN(new_n779_));
  INV_X1    g578(.A(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(G85gat), .B1(new_n780_), .B2(new_n437_), .ZN(new_n781_));
  NOR2_X1   g580(.A1(new_n756_), .A2(new_n670_), .ZN(new_n782_));
  AND2_X1   g581(.A1(new_n718_), .A2(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n470_), .A2(new_n416_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n781_), .B1(new_n783_), .B2(new_n784_), .ZN(G1336gat));
  AOI21_X1  g584(.A(G92gat), .B1(new_n780_), .B2(new_n467_), .ZN(new_n786_));
  AND3_X1   g585(.A1(new_n467_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n783_), .B2(new_n787_), .ZN(G1337gat));
  NOR3_X1   g587(.A1(new_n779_), .A2(new_n283_), .A3(new_n501_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n783_), .A2(new_n282_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n789_), .B1(new_n790_), .B2(G99gat), .ZN(new_n791_));
  XOR2_X1   g590(.A(new_n791_), .B(KEYINPUT51), .Z(G1338gat));
  XNOR2_X1  g591(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n793_));
  AOI21_X1  g592(.A(KEYINPUT43), .B1(new_n716_), .B2(KEYINPUT102), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n714_), .B(new_n708_), .C1(new_n472_), .C2(new_n645_), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n338_), .B(new_n782_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n718_), .A2(KEYINPUT108), .A3(new_n338_), .A4(new_n782_), .ZN(new_n799_));
  NAND3_X1  g598(.A1(new_n798_), .A2(G106gat), .A3(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(KEYINPUT52), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  NAND4_X1  g601(.A1(new_n798_), .A2(new_n799_), .A3(new_n802_), .A4(G106gat), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n801_), .A2(new_n803_), .ZN(new_n804_));
  AND4_X1   g603(.A1(new_n478_), .A2(new_n757_), .A3(new_n338_), .A4(new_n704_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n805_), .A2(KEYINPUT107), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(KEYINPUT107), .ZN(new_n807_));
  AND2_X1   g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  INV_X1    g607(.A(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n793_), .B1(new_n804_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(new_n793_), .ZN(new_n811_));
  AOI211_X1 g610(.A(new_n808_), .B(new_n811_), .C1(new_n801_), .C2(new_n803_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n810_), .A2(new_n812_), .ZN(G1339gat));
  INV_X1    g612(.A(G113gat), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n581_), .A2(new_n582_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n815_), .A2(new_n591_), .ZN(new_n816_));
  OR2_X1    g615(.A1(new_n816_), .A2(KEYINPUT111), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n586_), .B1(new_n581_), .B2(new_n585_), .ZN(new_n818_));
  NAND3_X1  g617(.A1(new_n818_), .A2(G229gat), .A3(G233gat), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n816_), .A2(KEYINPUT111), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n817_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n821_));
  AND2_X1   g620(.A1(new_n821_), .A2(new_n593_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n822_), .A2(new_n548_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n529_), .A2(new_n475_), .A3(new_n531_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT110), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT55), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NOR2_X1   g626(.A1(new_n825_), .A2(new_n826_), .ZN(new_n828_));
  OAI211_X1 g627(.A(new_n824_), .B(new_n827_), .C1(new_n532_), .C2(new_n828_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n532_), .A2(new_n828_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n545_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT56), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT56), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n833_), .B(new_n545_), .C1(new_n829_), .C2(new_n830_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n832_), .A2(new_n547_), .A3(new_n834_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n823_), .B1(new_n835_), .B2(new_n597_), .ZN(new_n836_));
  AND3_X1   g635(.A1(new_n836_), .A2(KEYINPUT57), .A3(new_n666_), .ZN(new_n837_));
  AOI21_X1  g636(.A(KEYINPUT57), .B1(new_n836_), .B2(new_n666_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n837_), .A2(new_n838_), .ZN(new_n839_));
  NAND4_X1  g638(.A1(new_n832_), .A2(new_n822_), .A3(new_n547_), .A4(new_n834_), .ZN(new_n840_));
  NOR2_X1   g639(.A1(KEYINPUT112), .A2(KEYINPUT58), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  AND2_X1   g642(.A1(new_n834_), .A2(new_n547_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n844_), .A2(new_n841_), .A3(new_n822_), .A4(new_n832_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n845_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n846_), .A2(new_n710_), .A3(new_n711_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT113), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n645_), .A2(KEYINPUT113), .A3(new_n846_), .ZN(new_n850_));
  NAND3_X1  g649(.A1(new_n839_), .A2(new_n849_), .A3(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT114), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n839_), .A2(new_n849_), .A3(KEYINPUT114), .A4(new_n850_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n853_), .A2(new_n660_), .A3(new_n854_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n712_), .A2(new_n597_), .A3(new_n753_), .A4(new_n670_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT54), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n469_), .A2(new_n437_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n814_), .B1(new_n861_), .B2(new_n597_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(KEYINPUT115), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(KEYINPUT59), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n839_), .A2(new_n847_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(new_n660_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n857_), .A2(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT59), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n867_), .A2(new_n868_), .A3(new_n860_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n864_), .A2(G113gat), .A3(new_n754_), .A4(new_n869_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT115), .ZN(new_n871_));
  OAI211_X1 g670(.A(new_n871_), .B(new_n814_), .C1(new_n861_), .C2(new_n597_), .ZN(new_n872_));
  AND3_X1   g671(.A1(new_n863_), .A2(new_n870_), .A3(new_n872_), .ZN(G1340gat));
  NAND3_X1  g672(.A1(new_n864_), .A2(new_n552_), .A3(new_n869_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT116), .B(G120gat), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n859_), .B1(new_n855_), .B2(new_n857_), .ZN(new_n877_));
  INV_X1    g676(.A(new_n875_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n878_), .A2(KEYINPUT60), .ZN(new_n879_));
  OAI21_X1  g678(.A(new_n878_), .B1(new_n753_), .B2(KEYINPUT60), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(KEYINPUT117), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n877_), .B(new_n881_), .C1(KEYINPUT117), .C2(new_n880_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n876_), .A2(new_n882_), .ZN(G1341gat));
  AOI21_X1  g682(.A(G127gat), .B1(new_n877_), .B2(new_n670_), .ZN(new_n884_));
  AND2_X1   g683(.A1(new_n864_), .A2(new_n869_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n886_), .A2(G127gat), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n670_), .A2(KEYINPUT118), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n887_), .B1(new_n888_), .B2(G127gat), .ZN(new_n889_));
  AOI21_X1  g688(.A(new_n884_), .B1(new_n885_), .B2(new_n889_), .ZN(G1342gat));
  NAND3_X1  g689(.A1(new_n858_), .A2(new_n665_), .A3(new_n860_), .ZN(new_n891_));
  INV_X1    g690(.A(G134gat), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n891_), .A2(new_n892_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(new_n712_), .A2(new_n892_), .ZN(new_n894_));
  OAI211_X1 g693(.A(new_n869_), .B(new_n894_), .C1(new_n877_), .C2(new_n868_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n893_), .A2(new_n895_), .ZN(new_n896_));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n896_), .A2(new_n897_), .ZN(new_n898_));
  NAND3_X1  g697(.A1(new_n893_), .A2(new_n895_), .A3(KEYINPUT119), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(new_n899_), .ZN(G1343gat));
  XOR2_X1   g699(.A(new_n856_), .B(KEYINPUT54), .Z(new_n901_));
  AOI21_X1  g700(.A(new_n670_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n901_), .B1(new_n902_), .B2(new_n854_), .ZN(new_n903_));
  NOR4_X1   g702(.A1(new_n467_), .A2(new_n470_), .A3(new_n337_), .A4(new_n282_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(KEYINPUT120), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n903_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n906_), .A2(new_n754_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n907_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n552_), .ZN(new_n909_));
  XNOR2_X1  g708(.A(new_n909_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g709(.A1(new_n906_), .A2(new_n670_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(KEYINPUT61), .B(G155gat), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n911_), .B(new_n912_), .ZN(G1346gat));
  AOI21_X1  g712(.A(G162gat), .B1(new_n906_), .B2(new_n665_), .ZN(new_n914_));
  AND2_X1   g713(.A1(new_n645_), .A2(G162gat), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n906_), .B2(new_n915_), .ZN(G1347gat));
  INV_X1    g715(.A(KEYINPUT62), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n467_), .A2(new_n470_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n918_), .A2(new_n468_), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n867_), .A2(new_n754_), .A3(new_n919_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT121), .ZN(new_n921_));
  NAND3_X1  g720(.A1(new_n920_), .A2(new_n921_), .A3(G169gat), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n921_), .B1(new_n920_), .B2(G169gat), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n917_), .B1(new_n923_), .B2(new_n924_), .ZN(new_n925_));
  INV_X1    g724(.A(new_n924_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n926_), .A2(KEYINPUT62), .A3(new_n922_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n349_), .A2(new_n350_), .ZN(new_n928_));
  OAI211_X1 g727(.A(new_n925_), .B(new_n927_), .C1(new_n928_), .C2(new_n920_), .ZN(G1348gat));
  NAND2_X1  g728(.A1(new_n867_), .A2(new_n919_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n930_), .ZN(new_n931_));
  AOI21_X1  g730(.A(G176gat), .B1(new_n931_), .B2(new_n552_), .ZN(new_n932_));
  OAI21_X1  g731(.A(KEYINPUT122), .B1(new_n903_), .B2(new_n338_), .ZN(new_n933_));
  INV_X1    g732(.A(KEYINPUT122), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n858_), .A2(new_n934_), .A3(new_n337_), .ZN(new_n935_));
  NOR2_X1   g734(.A1(new_n918_), .A2(new_n283_), .ZN(new_n936_));
  AND3_X1   g735(.A1(new_n933_), .A2(new_n935_), .A3(new_n936_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n753_), .A2(new_n207_), .ZN(new_n938_));
  AOI21_X1  g737(.A(new_n932_), .B1(new_n937_), .B2(new_n938_), .ZN(G1349gat));
  NOR3_X1   g738(.A1(new_n930_), .A2(new_n251_), .A3(new_n660_), .ZN(new_n940_));
  NAND4_X1  g739(.A1(new_n933_), .A2(new_n935_), .A3(new_n670_), .A4(new_n936_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n940_), .B1(new_n941_), .B2(new_n211_), .ZN(G1350gat));
  OAI21_X1  g741(.A(G190gat), .B1(new_n930_), .B2(new_n712_), .ZN(new_n943_));
  NAND2_X1  g742(.A1(new_n665_), .A2(new_n252_), .ZN(new_n944_));
  OAI21_X1  g743(.A(new_n943_), .B1(new_n930_), .B2(new_n944_), .ZN(G1351gat));
  NOR3_X1   g744(.A1(new_n437_), .A2(new_n282_), .A3(new_n337_), .ZN(new_n946_));
  OR2_X1    g745(.A1(new_n946_), .A2(KEYINPUT123), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n946_), .A2(KEYINPUT123), .ZN(new_n948_));
  NAND3_X1  g747(.A1(new_n947_), .A2(new_n467_), .A3(new_n948_), .ZN(new_n949_));
  OAI21_X1  g748(.A(KEYINPUT124), .B1(new_n903_), .B2(new_n949_), .ZN(new_n950_));
  INV_X1    g749(.A(KEYINPUT124), .ZN(new_n951_));
  INV_X1    g750(.A(new_n949_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n858_), .A2(new_n951_), .A3(new_n952_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n950_), .A2(new_n953_), .ZN(new_n954_));
  AOI21_X1  g753(.A(G197gat), .B1(new_n954_), .B2(new_n754_), .ZN(new_n955_));
  INV_X1    g754(.A(G197gat), .ZN(new_n956_));
  AOI211_X1 g755(.A(new_n956_), .B(new_n597_), .C1(new_n950_), .C2(new_n953_), .ZN(new_n957_));
  NOR2_X1   g756(.A1(new_n955_), .A2(new_n957_), .ZN(G1352gat));
  NAND2_X1  g757(.A1(new_n954_), .A2(new_n552_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n959_), .A2(G204gat), .ZN(new_n960_));
  INV_X1    g759(.A(G204gat), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n954_), .A2(new_n961_), .A3(new_n552_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n960_), .A2(new_n962_), .ZN(G1353gat));
  AOI21_X1  g762(.A(new_n660_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n954_), .A2(new_n964_), .ZN(new_n965_));
  NOR2_X1   g764(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n966_));
  XNOR2_X1  g765(.A(new_n966_), .B(KEYINPUT125), .ZN(new_n967_));
  INV_X1    g766(.A(new_n967_), .ZN(new_n968_));
  NAND2_X1  g767(.A1(new_n965_), .A2(new_n968_), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n954_), .A2(new_n964_), .A3(new_n967_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n969_), .A2(new_n970_), .ZN(G1354gat));
  NAND2_X1  g770(.A1(new_n954_), .A2(new_n665_), .ZN(new_n972_));
  INV_X1    g771(.A(G218gat), .ZN(new_n973_));
  NOR2_X1   g772(.A1(new_n712_), .A2(new_n973_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(KEYINPUT126), .ZN(new_n975_));
  AOI22_X1  g774(.A1(new_n972_), .A2(new_n973_), .B1(new_n954_), .B2(new_n975_), .ZN(G1355gat));
endmodule


