//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n685_, new_n686_, new_n687_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n773_, new_n774_, new_n776_, new_n777_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n817_, new_n818_, new_n819_, new_n820_, new_n821_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n883_, new_n885_,
    new_n886_, new_n887_, new_n889_, new_n890_, new_n891_, new_n893_,
    new_n894_, new_n895_, new_n896_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n924_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n937_, new_n938_, new_n940_, new_n941_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n965_, new_n966_, new_n967_, new_n968_;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT82), .ZN(new_n203_));
  OAI21_X1  g002(.A(KEYINPUT81), .B1(G141gat), .B2(G148gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  NOR3_X1   g005(.A1(KEYINPUT81), .A2(G141gat), .A3(G148gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n203_), .B1(new_n206_), .B2(new_n207_), .ZN(new_n208_));
  OR3_X1    g007(.A1(KEYINPUT81), .A2(G141gat), .A3(G148gat), .ZN(new_n209_));
  NAND4_X1  g008(.A1(new_n209_), .A2(KEYINPUT82), .A3(new_n205_), .A4(new_n204_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G141gat), .A2(G148gat), .ZN(new_n211_));
  INV_X1    g010(.A(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(G141gat), .ZN(new_n213_));
  INV_X1    g012(.A(G148gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  AOI22_X1  g014(.A1(new_n212_), .A2(KEYINPUT2), .B1(new_n215_), .B2(KEYINPUT3), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(KEYINPUT79), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT79), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G141gat), .A3(G148gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT2), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND4_X1  g020(.A1(new_n208_), .A2(new_n210_), .A3(new_n216_), .A4(new_n221_), .ZN(new_n222_));
  NOR2_X1   g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT80), .ZN(new_n224_));
  XNOR2_X1  g023(.A(new_n223_), .B(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(G155gat), .A2(G162gat), .ZN(new_n226_));
  AND2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n222_), .A2(new_n227_), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n217_), .A2(new_n219_), .A3(new_n215_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n230_));
  XNOR2_X1  g029(.A(new_n226_), .B(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n225_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n228_), .A2(new_n233_), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G127gat), .B(G134gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(G113gat), .B(G120gat), .ZN(new_n236_));
  AND2_X1   g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NOR2_X1   g036(.A1(new_n235_), .A2(new_n236_), .ZN(new_n238_));
  NOR2_X1   g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n234_), .A2(new_n239_), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n232_), .B1(new_n222_), .B2(new_n227_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n239_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(G225gat), .A2(G233gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n240_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G1gat), .B(G29gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  XNOR2_X1  g047(.A(G57gat), .B(G85gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(new_n250_), .ZN(new_n251_));
  AOI211_X1 g050(.A(new_n232_), .B(new_n239_), .C1(new_n222_), .C2(new_n227_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n242_), .B1(new_n228_), .B2(new_n233_), .ZN(new_n253_));
  INV_X1    g052(.A(KEYINPUT4), .ZN(new_n254_));
  NOR3_X1   g053(.A1(new_n252_), .A2(new_n253_), .A3(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n234_), .A2(new_n254_), .A3(new_n239_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n244_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  OAI211_X1 g057(.A(new_n245_), .B(new_n251_), .C1(new_n255_), .C2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(KEYINPUT33), .B1(new_n259_), .B2(KEYINPUT92), .ZN(new_n260_));
  OAI21_X1  g059(.A(new_n260_), .B1(KEYINPUT92), .B2(new_n259_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n261_), .A2(KEYINPUT93), .ZN(new_n262_));
  INV_X1    g061(.A(KEYINPUT93), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n260_), .B(new_n263_), .C1(KEYINPUT92), .C2(new_n259_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n240_), .A2(KEYINPUT4), .A3(new_n243_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n265_), .A2(new_n244_), .A3(new_n256_), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n240_), .A2(new_n243_), .A3(new_n257_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n266_), .A2(new_n250_), .A3(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n244_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n265_), .A2(new_n269_), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n270_), .A2(KEYINPUT33), .A3(new_n245_), .A4(new_n251_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n272_));
  NAND2_X1  g071(.A1(G226gat), .A2(G233gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT21), .ZN(new_n275_));
  INV_X1    g074(.A(G218gat), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(G211gat), .ZN(new_n277_));
  INV_X1    g076(.A(G211gat), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(G218gat), .ZN(new_n279_));
  AOI21_X1  g078(.A(new_n275_), .B1(new_n277_), .B2(new_n279_), .ZN(new_n280_));
  AND2_X1   g079(.A1(KEYINPUT84), .A2(G197gat), .ZN(new_n281_));
  NOR2_X1   g080(.A1(KEYINPUT84), .A2(G197gat), .ZN(new_n282_));
  OAI21_X1  g081(.A(G204gat), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NOR2_X1   g082(.A1(G197gat), .A2(G204gat), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n280_), .A2(new_n283_), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n277_), .A2(new_n279_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n283_), .A2(new_n285_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n288_), .B1(new_n289_), .B2(new_n275_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT84), .ZN(new_n291_));
  INV_X1    g090(.A(G197gat), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(KEYINPUT84), .A2(G197gat), .ZN(new_n294_));
  AOI21_X1  g093(.A(G204gat), .B1(new_n293_), .B2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT85), .ZN(new_n296_));
  INV_X1    g095(.A(G204gat), .ZN(new_n297_));
  OAI21_X1  g096(.A(new_n296_), .B1(new_n297_), .B2(G197gat), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n292_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n298_), .A2(new_n299_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT21), .B1(new_n295_), .B2(new_n300_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n287_), .B1(new_n290_), .B2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT89), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT22), .ZN(new_n304_));
  NOR2_X1   g103(.A1(new_n304_), .A2(G169gat), .ZN(new_n305_));
  INV_X1    g104(.A(G169gat), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n306_), .A2(KEYINPUT22), .ZN(new_n307_));
  OAI21_X1  g106(.A(new_n303_), .B1(new_n305_), .B2(new_n307_), .ZN(new_n308_));
  XOR2_X1   g107(.A(KEYINPUT78), .B(G176gat), .Z(new_n309_));
  NAND2_X1  g108(.A1(new_n306_), .A2(KEYINPUT22), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n304_), .A2(G169gat), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n310_), .A2(new_n311_), .A3(KEYINPUT89), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n308_), .A2(new_n309_), .A3(new_n312_), .ZN(new_n313_));
  AOI21_X1  g112(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(G183gat), .A2(G190gat), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n316_), .A2(new_n317_), .B1(G169gat), .B2(G176gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT25), .B(G183gat), .ZN(new_n319_));
  XNOR2_X1  g118(.A(KEYINPUT26), .B(G190gat), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n321_), .B1(G169gat), .B2(G176gat), .ZN(new_n322_));
  NOR2_X1   g121(.A1(G169gat), .A2(G176gat), .ZN(new_n323_));
  INV_X1    g122(.A(new_n323_), .ZN(new_n324_));
  AOI22_X1  g123(.A1(new_n319_), .A2(new_n320_), .B1(new_n322_), .B2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(G183gat), .ZN(new_n326_));
  INV_X1    g125(.A(G190gat), .ZN(new_n327_));
  OAI21_X1  g126(.A(KEYINPUT23), .B1(new_n326_), .B2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT23), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(G183gat), .A3(G190gat), .ZN(new_n330_));
  AOI22_X1  g129(.A1(new_n328_), .A2(new_n330_), .B1(new_n321_), .B2(new_n323_), .ZN(new_n331_));
  AOI22_X1  g130(.A1(new_n313_), .A2(new_n318_), .B1(new_n325_), .B2(new_n331_), .ZN(new_n332_));
  OAI21_X1  g131(.A(KEYINPUT20), .B1(new_n302_), .B2(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n297_), .B1(new_n293_), .B2(new_n294_), .ZN(new_n334_));
  OAI21_X1  g133(.A(new_n275_), .B1(new_n334_), .B2(new_n284_), .ZN(new_n335_));
  INV_X1    g134(.A(new_n288_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n301_), .A2(new_n335_), .A3(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n286_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n309_), .A2(new_n310_), .A3(new_n311_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n318_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n325_), .A2(new_n331_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n274_), .B1(new_n333_), .B2(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G8gat), .B(G36gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G64gat), .B(G92gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n345_), .B(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(KEYINPUT90), .B(KEYINPUT18), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n347_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT20), .ZN(new_n350_));
  AOI21_X1  g149(.A(new_n350_), .B1(new_n302_), .B2(new_n332_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n274_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n338_), .A2(new_n342_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n352_), .A3(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n344_), .A2(new_n349_), .A3(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n344_), .A2(new_n354_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n349_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n268_), .A2(new_n271_), .A3(new_n355_), .A4(new_n358_), .ZN(new_n359_));
  INV_X1    g158(.A(new_n359_), .ZN(new_n360_));
  NAND3_X1  g159(.A1(new_n262_), .A2(new_n264_), .A3(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n313_), .A2(new_n318_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n362_), .A2(new_n341_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT20), .B1(new_n338_), .B2(new_n363_), .ZN(new_n364_));
  AOI22_X1  g163(.A1(new_n318_), .A2(new_n339_), .B1(new_n325_), .B2(new_n331_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n302_), .A2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n274_), .B1(new_n364_), .B2(new_n366_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n350_), .B1(new_n338_), .B2(new_n363_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n302_), .A2(new_n365_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n368_), .A2(new_n352_), .A3(new_n369_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n349_), .A2(KEYINPUT32), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n371_), .A2(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n374_), .A2(KEYINPUT94), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT94), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n371_), .A2(new_n376_), .A3(new_n373_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n344_), .A2(new_n354_), .A3(new_n372_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n375_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n259_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n251_), .B1(new_n270_), .B2(new_n245_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NOR2_X1   g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G22gat), .B(G50gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(KEYINPUT28), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT83), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n388_));
  AND3_X1   g187(.A1(new_n241_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n387_), .B1(new_n241_), .B2(new_n388_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n386_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  OAI21_X1  g190(.A(KEYINPUT83), .B1(new_n234_), .B2(KEYINPUT29), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n241_), .A2(new_n387_), .A3(new_n388_), .ZN(new_n393_));
  NAND3_X1  g192(.A1(new_n392_), .A2(new_n393_), .A3(new_n385_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n338_), .B1(new_n241_), .B2(new_n388_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(G228gat), .A2(G233gat), .ZN(new_n397_));
  OR2_X1    g196(.A1(new_n397_), .A2(KEYINPUT86), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(KEYINPUT86), .ZN(new_n399_));
  AND2_X1   g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n338_), .B(new_n398_), .C1(new_n241_), .C2(new_n388_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n402_), .A2(new_n404_), .A3(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT87), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n395_), .A2(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n402_), .A2(new_n405_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n409_), .A2(new_n403_), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(new_n406_), .ZN(new_n411_));
  NOR2_X1   g210(.A1(new_n408_), .A2(new_n411_), .ZN(new_n412_));
  AOI22_X1  g211(.A1(new_n395_), .A2(new_n407_), .B1(new_n410_), .B2(new_n406_), .ZN(new_n413_));
  NOR2_X1   g212(.A1(new_n412_), .A2(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n383_), .A2(new_n414_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n361_), .A2(new_n415_), .ZN(new_n416_));
  XOR2_X1   g215(.A(G71gat), .B(G99gat), .Z(new_n417_));
  XNOR2_X1  g216(.A(new_n417_), .B(G43gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n365_), .B(new_n418_), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(new_n242_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(G227gat), .A2(G233gat), .ZN(new_n421_));
  INV_X1    g220(.A(G15gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n423_), .B(KEYINPUT30), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT31), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n420_), .B(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT27), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n349_), .B(KEYINPUT96), .ZN(new_n430_));
  AOI22_X1  g229(.A1(KEYINPUT97), .A2(new_n355_), .B1(new_n371_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT97), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n344_), .A2(new_n432_), .A3(new_n354_), .A4(new_n349_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n429_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n358_), .A2(new_n429_), .A3(new_n355_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT95), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n380_), .A2(new_n381_), .A3(new_n437_), .ZN(new_n438_));
  OAI21_X1  g237(.A(new_n245_), .B1(new_n255_), .B2(new_n258_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n439_), .A2(new_n250_), .ZN(new_n440_));
  AOI21_X1  g239(.A(KEYINPUT95), .B1(new_n440_), .B2(new_n259_), .ZN(new_n441_));
  OAI22_X1  g240(.A1(new_n434_), .A2(new_n436_), .B1(new_n438_), .B2(new_n441_), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n428_), .B1(new_n442_), .B2(new_n414_), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT98), .B1(new_n434_), .B2(new_n436_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n355_), .A2(KEYINPUT97), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n371_), .A2(new_n430_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n445_), .A2(new_n433_), .A3(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(KEYINPUT27), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT98), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n448_), .A2(new_n449_), .A3(new_n435_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n414_), .B1(new_n444_), .B2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n440_), .A2(KEYINPUT95), .A3(new_n259_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n437_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n427_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  AOI22_X1  g253(.A1(new_n416_), .A2(new_n443_), .B1(new_n451_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G1gat), .B(G8gat), .ZN(new_n456_));
  OR2_X1    g255(.A1(new_n456_), .A2(KEYINPUT74), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(KEYINPUT74), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(G15gat), .B(G22gat), .ZN(new_n460_));
  INV_X1    g259(.A(G1gat), .ZN(new_n461_));
  INV_X1    g260(.A(G8gat), .ZN(new_n462_));
  OAI21_X1  g261(.A(KEYINPUT14), .B1(new_n461_), .B2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n459_), .A2(new_n464_), .ZN(new_n465_));
  NAND4_X1  g264(.A1(new_n457_), .A2(new_n463_), .A3(new_n460_), .A4(new_n458_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G43gat), .B(G50gat), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  INV_X1    g268(.A(G36gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(G29gat), .ZN(new_n471_));
  INV_X1    g270(.A(G29gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n472_), .A2(G36gat), .ZN(new_n473_));
  AND3_X1   g272(.A1(new_n471_), .A2(new_n473_), .A3(KEYINPUT69), .ZN(new_n474_));
  AOI21_X1  g273(.A(KEYINPUT69), .B1(new_n471_), .B2(new_n473_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n469_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT69), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n472_), .A2(G36gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n470_), .A2(G29gat), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n477_), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n471_), .A2(new_n473_), .A3(KEYINPUT69), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n480_), .A2(new_n481_), .A3(new_n468_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n476_), .A2(new_n482_), .ZN(new_n483_));
  XNOR2_X1  g282(.A(new_n467_), .B(new_n483_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(G229gat), .A2(G233gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n476_), .A2(new_n482_), .A3(KEYINPUT15), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  AOI21_X1  g287(.A(KEYINPUT15), .B1(new_n476_), .B2(new_n482_), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n490_), .A2(new_n466_), .A3(new_n465_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n486_), .B1(new_n467_), .B2(new_n483_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n484_), .A2(new_n486_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G113gat), .B(G141gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(G169gat), .B(G197gat), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XOR2_X1   g295(.A(new_n493_), .B(new_n496_), .Z(new_n497_));
  OAI21_X1  g296(.A(new_n202_), .B1(new_n455_), .B2(new_n497_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n408_), .A2(new_n411_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n413_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NOR3_X1   g300(.A1(new_n434_), .A2(KEYINPUT98), .A3(new_n436_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n449_), .B1(new_n448_), .B2(new_n435_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n501_), .B(new_n454_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  OAI22_X1  g303(.A1(new_n379_), .A2(new_n382_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n359_), .B1(new_n261_), .B2(KEYINPUT93), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n505_), .B1(new_n506_), .B2(new_n264_), .ZN(new_n507_));
  AOI22_X1  g306(.A1(new_n448_), .A2(new_n435_), .B1(new_n453_), .B2(new_n452_), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n427_), .B1(new_n508_), .B2(new_n501_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n504_), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n497_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n510_), .A2(KEYINPUT99), .A3(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n498_), .A2(new_n512_), .ZN(new_n513_));
  INV_X1    g312(.A(KEYINPUT13), .ZN(new_n514_));
  NAND2_X1  g313(.A1(G99gat), .A2(G106gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(KEYINPUT6), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT6), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n517_), .A2(G99gat), .A3(G106gat), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n516_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(G99gat), .ZN(new_n520_));
  INV_X1    g319(.A(G106gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n520_), .A2(new_n521_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(KEYINPUT7), .ZN(new_n523_));
  NOR4_X1   g322(.A1(KEYINPUT65), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT65), .ZN(new_n525_));
  NOR2_X1   g324(.A1(G99gat), .A2(G106gat), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT7), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n525_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n519_), .B(new_n523_), .C1(new_n524_), .C2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G85gat), .B(G92gat), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT8), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n533_), .B1(new_n530_), .B2(KEYINPUT66), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n527_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT65), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n526_), .A2(new_n525_), .A3(new_n527_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  AOI22_X1  g339(.A1(new_n516_), .A2(new_n518_), .B1(new_n522_), .B2(KEYINPUT7), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n530_), .B1(new_n540_), .B2(new_n541_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n542_), .A2(new_n534_), .ZN(new_n543_));
  AND2_X1   g342(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n544_));
  NOR2_X1   g343(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n544_), .A2(new_n545_), .ZN(new_n546_));
  AOI22_X1  g345(.A1(new_n546_), .A2(new_n521_), .B1(new_n516_), .B2(new_n518_), .ZN(new_n547_));
  INV_X1    g346(.A(KEYINPUT9), .ZN(new_n548_));
  INV_X1    g347(.A(G92gat), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n548_), .A2(new_n549_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n548_), .A2(KEYINPUT64), .ZN(new_n551_));
  NOR2_X1   g350(.A1(new_n548_), .A2(KEYINPUT64), .ZN(new_n552_));
  OAI211_X1 g351(.A(new_n530_), .B(new_n550_), .C1(new_n551_), .C2(new_n552_), .ZN(new_n553_));
  AND2_X1   g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554_));
  NOR2_X1   g353(.A1(G85gat), .A2(G92gat), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n550_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n547_), .A2(new_n553_), .A3(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n536_), .A2(new_n543_), .A3(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G57gat), .B(G64gat), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT11), .ZN(new_n562_));
  XOR2_X1   g361(.A(G71gat), .B(G78gat), .Z(new_n563_));
  OR2_X1    g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NOR2_X1   g363(.A1(new_n561_), .A2(KEYINPUT11), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n562_), .A2(new_n563_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n567_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n560_), .A2(new_n568_), .A3(KEYINPUT12), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(KEYINPUT67), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT67), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n564_), .B(new_n571_), .C1(new_n565_), .C2(new_n566_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n569_), .B1(new_n573_), .B2(new_n560_), .ZN(new_n574_));
  AOI21_X1  g373(.A(KEYINPUT12), .B1(new_n573_), .B2(new_n560_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(G230gat), .A2(G233gat), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n576_), .A2(new_n577_), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n573_), .B(new_n560_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n577_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n578_), .A2(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G120gat), .B(G148gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT5), .ZN(new_n584_));
  XNOR2_X1  g383(.A(G176gat), .B(G204gat), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n584_), .B(new_n585_), .Z(new_n586_));
  NAND2_X1  g385(.A1(new_n582_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n586_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n578_), .A2(new_n581_), .A3(new_n588_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n587_), .A2(KEYINPUT68), .A3(new_n589_), .ZN(new_n590_));
  NOR3_X1   g389(.A1(new_n574_), .A2(new_n575_), .A3(new_n580_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n591_), .B1(new_n580_), .B2(new_n579_), .ZN(new_n592_));
  NOR3_X1   g391(.A1(new_n592_), .A2(KEYINPUT68), .A3(new_n588_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n514_), .B1(new_n590_), .B2(new_n593_), .ZN(new_n594_));
  INV_X1    g393(.A(new_n593_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n587_), .A2(KEYINPUT68), .A3(new_n589_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n595_), .A2(new_n596_), .A3(KEYINPUT13), .ZN(new_n597_));
  AND2_X1   g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  AND2_X1   g397(.A1(G231gat), .A2(G233gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n467_), .B(new_n599_), .ZN(new_n600_));
  OR2_X1    g399(.A1(new_n600_), .A2(new_n567_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n600_), .A2(new_n567_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(KEYINPUT67), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n601_), .A2(new_n571_), .A3(new_n602_), .ZN(new_n605_));
  XOR2_X1   g404(.A(G127gat), .B(G155gat), .Z(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT16), .ZN(new_n607_));
  XNOR2_X1  g406(.A(G183gat), .B(G211gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n607_), .B(new_n608_), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT17), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n604_), .A2(new_n605_), .A3(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(KEYINPUT75), .B(KEYINPUT17), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n609_), .A2(new_n612_), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n613_), .B(KEYINPUT76), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n614_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n611_), .A2(KEYINPUT77), .A3(new_n615_), .ZN(new_n616_));
  INV_X1    g415(.A(new_n616_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT77), .B1(new_n611_), .B2(new_n615_), .ZN(new_n618_));
  OR2_X1    g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT15), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n483_), .A2(new_n620_), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n559_), .B1(new_n542_), .B2(new_n534_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n529_), .A2(new_n531_), .A3(new_n534_), .ZN(new_n623_));
  OAI211_X1 g422(.A(new_n487_), .B(new_n621_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n624_));
  NAND4_X1  g423(.A1(new_n536_), .A2(new_n543_), .A3(new_n483_), .A4(new_n559_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(G232gat), .A2(G233gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n626_), .B(KEYINPUT34), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  INV_X1    g427(.A(KEYINPUT35), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n628_), .A2(new_n629_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n624_), .A2(new_n625_), .A3(new_n630_), .ZN(new_n631_));
  INV_X1    g430(.A(KEYINPUT70), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n632_), .B1(new_n490_), .B2(new_n560_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n628_), .A2(new_n629_), .ZN(new_n634_));
  INV_X1    g433(.A(new_n634_), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n631_), .B1(new_n633_), .B2(new_n635_), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n624_), .A2(new_n632_), .A3(new_n634_), .A4(new_n625_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(G190gat), .B(G218gat), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT71), .ZN(new_n639_));
  XOR2_X1   g438(.A(G134gat), .B(G162gat), .Z(new_n640_));
  XNOR2_X1  g439(.A(new_n639_), .B(new_n640_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n641_), .A2(KEYINPUT36), .ZN(new_n642_));
  INV_X1    g441(.A(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n641_), .A2(KEYINPUT36), .ZN(new_n644_));
  NAND4_X1  g443(.A1(new_n636_), .A2(new_n637_), .A3(new_n643_), .A4(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT73), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n646_), .A2(KEYINPUT37), .ZN(new_n647_));
  AND3_X1   g446(.A1(new_n624_), .A2(new_n625_), .A3(new_n630_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n635_), .B1(new_n624_), .B2(KEYINPUT70), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n637_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n642_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT72), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n650_), .A2(KEYINPUT72), .A3(new_n642_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n647_), .B1(new_n655_), .B2(new_n645_), .ZN(new_n656_));
  AOI211_X1 g455(.A(new_n652_), .B(new_n643_), .C1(new_n636_), .C2(new_n637_), .ZN(new_n657_));
  AOI21_X1  g456(.A(KEYINPUT72), .B1(new_n650_), .B2(new_n642_), .ZN(new_n658_));
  OAI21_X1  g457(.A(new_n645_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT37), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n660_), .B1(new_n645_), .B2(KEYINPUT73), .ZN(new_n661_));
  NOR2_X1   g460(.A1(new_n659_), .A2(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n656_), .A2(new_n662_), .ZN(new_n663_));
  NOR3_X1   g462(.A1(new_n598_), .A2(new_n619_), .A3(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n513_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n438_), .A2(new_n441_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n666_), .A2(new_n461_), .A3(new_n667_), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT38), .ZN(new_n669_));
  AND2_X1   g468(.A1(new_n668_), .A2(new_n669_), .ZN(new_n670_));
  NOR2_X1   g469(.A1(new_n668_), .A2(new_n669_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n659_), .ZN(new_n672_));
  NOR3_X1   g471(.A1(new_n455_), .A2(new_n619_), .A3(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n598_), .A2(new_n497_), .ZN(new_n674_));
  AND2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(new_n461_), .B1(new_n675_), .B2(new_n667_), .ZN(new_n676_));
  OR3_X1    g475(.A1(new_n670_), .A2(new_n671_), .A3(new_n676_), .ZN(G1324gat));
  NOR2_X1   g476(.A1(new_n502_), .A2(new_n503_), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n462_), .B1(new_n675_), .B2(new_n678_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT39), .Z(new_n680_));
  NAND3_X1  g479(.A1(new_n666_), .A2(new_n462_), .A3(new_n678_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n683_));
  XNOR2_X1  g482(.A(new_n682_), .B(new_n683_), .ZN(G1325gat));
  AOI21_X1  g483(.A(new_n422_), .B1(new_n675_), .B2(new_n428_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n685_), .B(KEYINPUT41), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n666_), .A2(new_n422_), .A3(new_n428_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(new_n687_), .ZN(G1326gat));
  INV_X1    g487(.A(G22gat), .ZN(new_n689_));
  XNOR2_X1  g488(.A(new_n501_), .B(KEYINPUT101), .ZN(new_n690_));
  INV_X1    g489(.A(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n689_), .B1(new_n675_), .B2(new_n691_), .ZN(new_n692_));
  XOR2_X1   g491(.A(new_n692_), .B(KEYINPUT42), .Z(new_n693_));
  NAND3_X1  g492(.A1(new_n666_), .A2(new_n689_), .A3(new_n691_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT102), .Z(G1327gat));
  NAND2_X1  g495(.A1(new_n619_), .A2(new_n672_), .ZN(new_n697_));
  INV_X1    g496(.A(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n594_), .A2(new_n597_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n698_), .A2(new_n699_), .ZN(new_n700_));
  AOI21_X1  g499(.A(new_n700_), .B1(new_n498_), .B2(new_n512_), .ZN(new_n701_));
  AOI21_X1  g500(.A(G29gat), .B1(new_n701_), .B2(new_n667_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n699_), .A2(new_n511_), .A3(new_n619_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n659_), .A2(new_n661_), .ZN(new_n704_));
  OAI221_X1 g503(.A(new_n645_), .B1(KEYINPUT73), .B2(new_n660_), .C1(new_n657_), .C2(new_n658_), .ZN(new_n705_));
  AND3_X1   g504(.A1(new_n704_), .A2(new_n705_), .A3(KEYINPUT103), .ZN(new_n706_));
  AOI21_X1  g505(.A(KEYINPUT103), .B1(new_n704_), .B2(new_n705_), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(KEYINPUT43), .B1(new_n455_), .B2(new_n708_), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n510_), .A2(new_n710_), .A3(new_n663_), .ZN(new_n711_));
  AOI21_X1  g510(.A(new_n703_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n712_), .A2(new_n713_), .A3(KEYINPUT44), .ZN(new_n714_));
  AND3_X1   g513(.A1(new_n699_), .A2(new_n511_), .A3(new_n619_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n716_));
  OAI21_X1  g515(.A(new_n716_), .B1(new_n656_), .B2(new_n662_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n704_), .A2(new_n705_), .A3(KEYINPUT103), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n710_), .B1(new_n510_), .B2(new_n719_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n704_), .A2(new_n705_), .A3(new_n710_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n416_), .A2(new_n443_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n721_), .B1(new_n722_), .B2(new_n504_), .ZN(new_n723_));
  OAI211_X1 g522(.A(KEYINPUT44), .B(new_n715_), .C1(new_n720_), .C2(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT104), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n715_), .B1(new_n720_), .B2(new_n723_), .ZN(new_n727_));
  AOI22_X1  g526(.A1(new_n714_), .A2(new_n725_), .B1(new_n726_), .B2(new_n727_), .ZN(new_n728_));
  INV_X1    g527(.A(new_n667_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n729_), .A2(new_n472_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n702_), .B1(new_n728_), .B2(new_n730_), .ZN(G1328gat));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n732_));
  INV_X1    g531(.A(new_n678_), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n727_), .B2(new_n726_), .ZN(new_n734_));
  AOI21_X1  g533(.A(new_n713_), .B1(new_n712_), .B2(KEYINPUT44), .ZN(new_n735_));
  NOR2_X1   g534(.A1(new_n724_), .A2(KEYINPUT104), .ZN(new_n736_));
  OAI211_X1 g535(.A(new_n732_), .B(new_n734_), .C1(new_n735_), .C2(new_n736_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n737_), .A2(G36gat), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n714_), .A2(new_n725_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n732_), .B1(new_n739_), .B2(new_n734_), .ZN(new_n740_));
  OAI21_X1  g539(.A(KEYINPUT106), .B1(new_n738_), .B2(new_n740_), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n734_), .B1(new_n735_), .B2(new_n736_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT105), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n744_));
  NAND4_X1  g543(.A1(new_n743_), .A2(new_n744_), .A3(G36gat), .A4(new_n737_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT107), .ZN(new_n747_));
  NOR2_X1   g546(.A1(new_n733_), .A2(G36gat), .ZN(new_n748_));
  AND3_X1   g547(.A1(new_n701_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n747_), .B1(new_n701_), .B2(new_n748_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n746_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n701_), .A2(new_n748_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(KEYINPUT107), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n701_), .A2(new_n747_), .A3(new_n748_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n753_), .A2(new_n754_), .A3(KEYINPUT45), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n751_), .A2(new_n755_), .ZN(new_n756_));
  NAND3_X1  g555(.A1(new_n741_), .A2(new_n745_), .A3(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT46), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(KEYINPUT108), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n758_), .A2(KEYINPUT108), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n757_), .A2(new_n759_), .A3(new_n760_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n751_), .A2(new_n755_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n743_), .A2(G36gat), .A3(new_n737_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n762_), .B1(new_n763_), .B2(KEYINPUT106), .ZN(new_n764_));
  NAND4_X1  g563(.A1(new_n764_), .A2(KEYINPUT108), .A3(new_n758_), .A4(new_n745_), .ZN(new_n765_));
  AND2_X1   g564(.A1(new_n761_), .A2(new_n765_), .ZN(G1329gat));
  NAND3_X1  g565(.A1(new_n728_), .A2(G43gat), .A3(new_n428_), .ZN(new_n767_));
  XOR2_X1   g566(.A(KEYINPUT109), .B(G43gat), .Z(new_n768_));
  INV_X1    g567(.A(new_n701_), .ZN(new_n769_));
  OAI21_X1  g568(.A(new_n768_), .B1(new_n769_), .B2(new_n427_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n767_), .A2(new_n770_), .ZN(new_n771_));
  XNOR2_X1  g570(.A(new_n771_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g571(.A(G50gat), .B1(new_n701_), .B2(new_n691_), .ZN(new_n773_));
  AND2_X1   g572(.A1(new_n414_), .A2(G50gat), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n728_), .B2(new_n774_), .ZN(G1331gat));
  NOR2_X1   g574(.A1(new_n699_), .A2(new_n511_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n673_), .A2(new_n776_), .ZN(new_n777_));
  OAI21_X1  g576(.A(G57gat), .B1(new_n777_), .B2(new_n729_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n779_));
  NOR3_X1   g578(.A1(new_n455_), .A2(new_n779_), .A3(new_n511_), .ZN(new_n780_));
  AOI21_X1  g579(.A(KEYINPUT110), .B1(new_n510_), .B2(new_n497_), .ZN(new_n781_));
  NOR3_X1   g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n699_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n619_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n663_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  OR2_X1    g584(.A1(new_n729_), .A2(G57gat), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n778_), .B1(new_n785_), .B2(new_n786_), .ZN(G1332gat));
  OAI21_X1  g586(.A(G64gat), .B1(new_n777_), .B2(new_n733_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT48), .ZN(new_n789_));
  OR2_X1    g588(.A1(new_n733_), .A2(G64gat), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n789_), .B1(new_n785_), .B2(new_n790_), .ZN(G1333gat));
  OAI21_X1  g590(.A(G71gat), .B1(new_n777_), .B2(new_n427_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT49), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n427_), .A2(G71gat), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n785_), .B2(new_n794_), .ZN(G1334gat));
  OAI21_X1  g594(.A(G78gat), .B1(new_n777_), .B2(new_n690_), .ZN(new_n796_));
  XOR2_X1   g595(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n797_));
  XNOR2_X1  g596(.A(new_n796_), .B(new_n797_), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n690_), .A2(G78gat), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n785_), .B2(new_n799_), .ZN(G1335gat));
  NAND2_X1  g599(.A1(new_n776_), .A2(new_n619_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n709_), .B2(new_n711_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n667_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(G85gat), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n782_), .A2(new_n698_), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n729_), .A2(G85gat), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n804_), .B1(new_n805_), .B2(new_n806_), .ZN(G1336gat));
  OAI21_X1  g606(.A(new_n549_), .B1(new_n805_), .B2(new_n733_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT112), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n678_), .A2(G92gat), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT113), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n809_), .B1(new_n802_), .B2(new_n811_), .ZN(G1337gat));
  NOR4_X1   g611(.A1(new_n805_), .A2(new_n427_), .A3(new_n545_), .A4(new_n544_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n520_), .B1(new_n802_), .B2(new_n428_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  XOR2_X1   g614(.A(new_n815_), .B(KEYINPUT51), .Z(G1338gat));
  NOR3_X1   g615(.A1(new_n805_), .A2(G106gat), .A3(new_n501_), .ZN(new_n817_));
  XOR2_X1   g616(.A(new_n817_), .B(KEYINPUT114), .Z(new_n818_));
  AOI21_X1  g617(.A(new_n521_), .B1(new_n802_), .B2(new_n414_), .ZN(new_n819_));
  XOR2_X1   g618(.A(new_n819_), .B(KEYINPUT52), .Z(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT53), .ZN(G1339gat));
  AND2_X1   g621(.A1(new_n451_), .A2(new_n428_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n823_), .A2(new_n667_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT118), .ZN(new_n825_));
  AOI21_X1  g624(.A(KEYINPUT59), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT56), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n580_), .B1(new_n574_), .B2(new_n575_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(KEYINPUT55), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(new_n578_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n576_), .A2(KEYINPUT55), .A3(new_n577_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n588_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n827_), .B1(new_n832_), .B2(KEYINPUT115), .ZN(new_n833_));
  AOI21_X1  g632(.A(new_n591_), .B1(KEYINPUT55), .B2(new_n828_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n831_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n586_), .B1(new_n834_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n836_), .A2(new_n837_), .A3(KEYINPUT56), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n497_), .B1(new_n592_), .B2(new_n588_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n833_), .A2(new_n838_), .A3(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n590_), .A2(new_n593_), .ZN(new_n842_));
  AOI21_X1  g641(.A(new_n496_), .B1(new_n484_), .B2(new_n485_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n485_), .B1(new_n467_), .B2(new_n483_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n491_), .A2(new_n844_), .ZN(new_n845_));
  AOI22_X1  g644(.A1(new_n493_), .A2(new_n496_), .B1(new_n843_), .B2(new_n845_), .ZN(new_n846_));
  AOI22_X1  g645(.A1(new_n840_), .A2(new_n841_), .B1(new_n842_), .B2(new_n846_), .ZN(new_n847_));
  NAND4_X1  g646(.A1(new_n833_), .A2(new_n838_), .A3(KEYINPUT116), .A4(new_n839_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n672_), .B1(new_n847_), .B2(new_n848_), .ZN(new_n849_));
  AND2_X1   g648(.A1(new_n849_), .A2(KEYINPUT57), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n589_), .A2(new_n846_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n851_), .B1(new_n836_), .B2(KEYINPUT56), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n832_), .A2(new_n827_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(KEYINPUT58), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(KEYINPUT117), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n852_), .A2(new_n856_), .A3(KEYINPUT58), .A4(new_n853_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(KEYINPUT58), .B1(new_n852_), .B2(new_n853_), .ZN(new_n859_));
  NOR2_X1   g658(.A1(new_n784_), .A2(new_n859_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n858_), .A2(new_n860_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n849_), .B2(KEYINPUT57), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT119), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n850_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n861_), .B(KEYINPUT119), .C1(new_n849_), .C2(KEYINPUT57), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n783_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n664_), .A2(new_n497_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n867_), .B(new_n868_), .ZN(new_n869_));
  OAI221_X1 g668(.A(new_n826_), .B1(new_n825_), .B2(new_n824_), .C1(new_n866_), .C2(new_n869_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n867_), .B(KEYINPUT54), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n619_), .B1(new_n850_), .B2(new_n862_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n729_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n823_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(KEYINPUT59), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n870_), .A2(new_n875_), .A3(new_n511_), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n876_), .A2(G113gat), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n497_), .A2(G113gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n874_), .B2(new_n878_), .ZN(G1340gat));
  AND3_X1   g678(.A1(new_n870_), .A2(new_n875_), .A3(new_n598_), .ZN(new_n880_));
  INV_X1    g679(.A(G120gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n881_), .B1(new_n699_), .B2(KEYINPUT60), .ZN(new_n882_));
  OAI21_X1  g681(.A(new_n882_), .B1(KEYINPUT60), .B2(new_n881_), .ZN(new_n883_));
  OAI22_X1  g682(.A1(new_n880_), .A2(new_n881_), .B1(new_n874_), .B2(new_n883_), .ZN(G1341gat));
  NAND3_X1  g683(.A1(new_n870_), .A2(new_n875_), .A3(new_n783_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n885_), .A2(G127gat), .ZN(new_n886_));
  OR2_X1    g685(.A1(new_n619_), .A2(G127gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n886_), .B1(new_n874_), .B2(new_n887_), .ZN(G1342gat));
  NAND3_X1  g687(.A1(new_n870_), .A2(new_n875_), .A3(new_n663_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(G134gat), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n659_), .A2(G134gat), .ZN(new_n891_));
  OAI21_X1  g690(.A(new_n890_), .B1(new_n874_), .B2(new_n891_), .ZN(G1343gat));
  NOR3_X1   g691(.A1(new_n678_), .A2(new_n501_), .A3(new_n428_), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n873_), .A2(new_n893_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n497_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(KEYINPUT120), .B(G141gat), .ZN(new_n896_));
  XNOR2_X1  g695(.A(new_n895_), .B(new_n896_), .ZN(G1344gat));
  NOR2_X1   g696(.A1(new_n894_), .A2(new_n699_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(new_n214_), .ZN(G1345gat));
  NOR2_X1   g698(.A1(new_n894_), .A2(new_n619_), .ZN(new_n900_));
  XOR2_X1   g699(.A(KEYINPUT61), .B(G155gat), .Z(new_n901_));
  XNOR2_X1  g700(.A(new_n900_), .B(new_n901_), .ZN(G1346gat));
  INV_X1    g701(.A(new_n894_), .ZN(new_n903_));
  AND3_X1   g702(.A1(new_n903_), .A2(G162gat), .A3(new_n719_), .ZN(new_n904_));
  AOI21_X1  g703(.A(G162gat), .B1(new_n903_), .B2(new_n672_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1347gat));
  NAND2_X1  g705(.A1(new_n862_), .A2(new_n863_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n850_), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n907_), .A2(new_n908_), .A3(new_n865_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n869_), .B1(new_n909_), .B2(new_n619_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n678_), .A2(new_n454_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n691_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n912_), .ZN(new_n913_));
  OAI21_X1  g712(.A(KEYINPUT121), .B1(new_n910_), .B2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT121), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n915_), .B(new_n912_), .C1(new_n866_), .C2(new_n869_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n914_), .A2(new_n916_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n917_), .A2(new_n511_), .A3(new_n308_), .A4(new_n312_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT62), .ZN(new_n919_));
  OAI211_X1 g718(.A(new_n511_), .B(new_n912_), .C1(new_n866_), .C2(new_n869_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n919_), .B1(new_n920_), .B2(G169gat), .ZN(new_n921_));
  AND3_X1   g720(.A1(new_n920_), .A2(new_n919_), .A3(G169gat), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n918_), .B1(new_n921_), .B2(new_n922_), .ZN(G1348gat));
  AOI21_X1  g722(.A(new_n414_), .B1(new_n871_), .B2(new_n872_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n911_), .ZN(new_n925_));
  AND4_X1   g724(.A1(G176gat), .A2(new_n924_), .A3(new_n598_), .A4(new_n925_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n917_), .A2(new_n598_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n926_), .B1(new_n927_), .B2(new_n309_), .ZN(G1349gat));
  NOR2_X1   g727(.A1(new_n619_), .A2(new_n319_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n917_), .A2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(KEYINPUT122), .ZN(new_n931_));
  NOR2_X1   g730(.A1(new_n619_), .A2(new_n911_), .ZN(new_n932_));
  AOI21_X1  g731(.A(G183gat), .B1(new_n924_), .B2(new_n932_), .ZN(new_n933_));
  INV_X1    g732(.A(new_n933_), .ZN(new_n934_));
  NAND3_X1  g733(.A1(new_n930_), .A2(new_n931_), .A3(new_n934_), .ZN(new_n935_));
  INV_X1    g734(.A(new_n929_), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n936_), .B1(new_n914_), .B2(new_n916_), .ZN(new_n937_));
  OAI21_X1  g736(.A(KEYINPUT122), .B1(new_n937_), .B2(new_n933_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n935_), .A2(new_n938_), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n917_), .A2(new_n320_), .A3(new_n672_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n784_), .B1(new_n914_), .B2(new_n916_), .ZN(new_n941_));
  OAI21_X1  g740(.A(new_n940_), .B1(new_n327_), .B2(new_n941_), .ZN(G1351gat));
  NAND2_X1  g741(.A1(new_n871_), .A2(new_n872_), .ZN(new_n943_));
  NOR4_X1   g742(.A1(new_n733_), .A2(new_n501_), .A3(new_n667_), .A4(new_n428_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n943_), .A2(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n945_), .A2(new_n497_), .ZN(new_n946_));
  XNOR2_X1  g745(.A(new_n946_), .B(new_n292_), .ZN(G1352gat));
  NOR2_X1   g746(.A1(new_n945_), .A2(new_n699_), .ZN(new_n948_));
  INV_X1    g747(.A(KEYINPUT123), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n949_), .B2(new_n297_), .ZN(new_n950_));
  XOR2_X1   g749(.A(KEYINPUT123), .B(G204gat), .Z(new_n951_));
  OAI21_X1  g750(.A(new_n950_), .B1(new_n948_), .B2(new_n951_), .ZN(G1353gat));
  NAND3_X1  g751(.A1(new_n943_), .A2(new_n783_), .A3(new_n944_), .ZN(new_n953_));
  XNOR2_X1  g752(.A(KEYINPUT63), .B(G211gat), .ZN(new_n954_));
  OR2_X1    g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n956_));
  NOR2_X1   g755(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n957_));
  AND3_X1   g756(.A1(new_n953_), .A2(new_n956_), .A3(new_n957_), .ZN(new_n958_));
  AOI21_X1  g757(.A(new_n956_), .B1(new_n953_), .B2(new_n957_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n955_), .B1(new_n958_), .B2(new_n959_), .ZN(new_n960_));
  NAND2_X1  g759(.A1(new_n960_), .A2(KEYINPUT125), .ZN(new_n961_));
  INV_X1    g760(.A(KEYINPUT125), .ZN(new_n962_));
  OAI211_X1 g761(.A(new_n955_), .B(new_n962_), .C1(new_n958_), .C2(new_n959_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n961_), .A2(new_n963_), .ZN(G1354gat));
  XOR2_X1   g763(.A(KEYINPUT127), .B(G218gat), .Z(new_n965_));
  NOR3_X1   g764(.A1(new_n945_), .A2(new_n784_), .A3(new_n965_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n945_), .A2(new_n659_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(new_n967_), .B(KEYINPUT126), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n966_), .B1(new_n968_), .B2(new_n965_), .ZN(G1355gat));
endmodule


