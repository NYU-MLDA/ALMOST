//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n797_, new_n798_, new_n799_, new_n800_, new_n802_,
    new_n803_, new_n805_, new_n806_, new_n807_, new_n808_, new_n809_,
    new_n810_, new_n811_, new_n813_, new_n814_, new_n815_, new_n817_,
    new_n818_, new_n819_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n830_, new_n831_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n936_, new_n938_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n946_, new_n947_, new_n948_, new_n949_,
    new_n950_, new_n951_, new_n952_, new_n953_, new_n954_, new_n955_,
    new_n956_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n973_, new_n974_, new_n976_, new_n977_,
    new_n979_, new_n980_, new_n982_, new_n983_, new_n984_, new_n986_,
    new_n987_, new_n988_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_;
  NAND2_X1  g000(.A1(G225gat), .A2(G233gat), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NOR2_X1   g003(.A1(G155gat), .A2(G162gat), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  AOI21_X1  g005(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n207_), .A2(KEYINPUT87), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT3), .ZN(new_n209_));
  NOR3_X1   g008(.A1(new_n209_), .A2(G141gat), .A3(G148gat), .ZN(new_n210_));
  INV_X1    g009(.A(G141gat), .ZN(new_n211_));
  INV_X1    g010(.A(G148gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT3), .B1(new_n211_), .B2(new_n212_), .ZN(new_n213_));
  OAI21_X1  g012(.A(new_n208_), .B1(new_n210_), .B2(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n215_), .B1(new_n207_), .B2(KEYINPUT87), .ZN(new_n216_));
  OAI21_X1  g015(.A(new_n206_), .B1(new_n214_), .B2(new_n216_), .ZN(new_n217_));
  NOR3_X1   g016(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT1), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n211_), .A2(new_n212_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n221_));
  OAI211_X1 g020(.A(new_n219_), .B(new_n220_), .C1(new_n221_), .C2(new_n203_), .ZN(new_n222_));
  OR2_X1    g021(.A1(new_n218_), .A2(new_n222_), .ZN(new_n223_));
  XNOR2_X1  g022(.A(G127gat), .B(G134gat), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(G120gat), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(G113gat), .ZN(new_n227_));
  INV_X1    g026(.A(G113gat), .ZN(new_n228_));
  NAND2_X1  g027(.A1(new_n228_), .A2(G120gat), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT86), .ZN(new_n230_));
  AND3_X1   g029(.A1(new_n227_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n230_), .B1(new_n227_), .B2(new_n229_), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n225_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NOR2_X1   g032(.A1(new_n228_), .A2(G120gat), .ZN(new_n234_));
  NOR2_X1   g033(.A1(new_n226_), .A2(G113gat), .ZN(new_n235_));
  OAI21_X1  g034(.A(KEYINPUT86), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n227_), .A2(new_n229_), .A3(new_n230_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n236_), .A2(new_n224_), .A3(new_n237_), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n217_), .A2(new_n223_), .B1(new_n233_), .B2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n240_));
  AOI21_X1  g039(.A(new_n202_), .B1(new_n239_), .B2(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(new_n238_), .ZN(new_n242_));
  AOI21_X1  g041(.A(new_n224_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n243_));
  OR2_X1    g042(.A1(new_n204_), .A2(new_n205_), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n211_), .A2(new_n212_), .A3(KEYINPUT3), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n209_), .B1(G141gat), .B2(G148gat), .ZN(new_n246_));
  AOI22_X1  g045(.A1(new_n245_), .A2(new_n246_), .B1(new_n207_), .B2(KEYINPUT87), .ZN(new_n247_));
  AND3_X1   g046(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT2), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n220_), .A2(new_n249_), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT87), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n248_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n244_), .B1(new_n247_), .B2(new_n252_), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n218_), .A2(new_n222_), .ZN(new_n254_));
  OAI22_X1  g053(.A1(new_n242_), .A2(new_n243_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  NAND4_X1  g054(.A1(new_n217_), .A2(new_n223_), .A3(new_n238_), .A4(new_n233_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n255_), .A2(new_n256_), .A3(KEYINPUT4), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n241_), .A2(new_n257_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n255_), .A2(new_n256_), .A3(new_n202_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(G57gat), .B(G85gat), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XOR2_X1   g064(.A(KEYINPUT97), .B(KEYINPUT0), .Z(new_n266_));
  NAND2_X1  g065(.A1(new_n266_), .A2(new_n262_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G1gat), .B(G29gat), .ZN(new_n268_));
  INV_X1    g067(.A(new_n268_), .ZN(new_n269_));
  AND3_X1   g068(.A1(new_n265_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n269_), .B1(new_n265_), .B2(new_n267_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n261_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n265_), .A2(new_n267_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(new_n273_), .A2(new_n268_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n265_), .A2(new_n267_), .A3(new_n269_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n274_), .A2(new_n260_), .A3(new_n275_), .ZN(new_n276_));
  AND2_X1   g075(.A1(new_n272_), .A2(new_n276_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n258_), .A2(new_n259_), .A3(new_n277_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n277_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT101), .ZN(new_n280_));
  OAI21_X1  g079(.A(new_n278_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  AND2_X1   g080(.A1(new_n255_), .A2(new_n256_), .ZN(new_n282_));
  AOI22_X1  g081(.A1(new_n282_), .A2(new_n202_), .B1(new_n241_), .B2(new_n257_), .ZN(new_n283_));
  NOR3_X1   g082(.A1(new_n283_), .A2(KEYINPUT101), .A3(new_n277_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT102), .B1(new_n281_), .B2(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(KEYINPUT101), .B1(new_n283_), .B2(new_n277_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(new_n279_), .A2(new_n280_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT102), .ZN(new_n288_));
  NAND4_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .A4(new_n278_), .ZN(new_n289_));
  AND2_X1   g088(.A1(new_n285_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n217_), .A2(new_n223_), .ZN(new_n291_));
  NOR2_X1   g090(.A1(new_n291_), .A2(KEYINPUT29), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G22gat), .B(G50gat), .ZN(new_n293_));
  XOR2_X1   g092(.A(new_n293_), .B(KEYINPUT28), .Z(new_n294_));
  NOR2_X1   g093(.A1(new_n292_), .A2(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n292_), .A2(new_n294_), .ZN(new_n297_));
  AOI21_X1  g096(.A(KEYINPUT93), .B1(new_n296_), .B2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n291_), .A2(KEYINPUT29), .ZN(new_n299_));
  INV_X1    g098(.A(G218gat), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(G211gat), .ZN(new_n301_));
  INV_X1    g100(.A(G211gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G218gat), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n301_), .A2(new_n303_), .A3(KEYINPUT91), .ZN(new_n304_));
  INV_X1    g103(.A(new_n304_), .ZN(new_n305_));
  AOI21_X1  g104(.A(KEYINPUT91), .B1(new_n301_), .B2(new_n303_), .ZN(new_n306_));
  NOR2_X1   g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT92), .ZN(new_n308_));
  INV_X1    g107(.A(G204gat), .ZN(new_n309_));
  OR2_X1    g108(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n311_));
  AOI21_X1  g110(.A(new_n309_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(G197gat), .A2(G204gat), .ZN(new_n313_));
  OAI21_X1  g112(.A(new_n308_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n311_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(KEYINPUT90), .A2(G197gat), .ZN(new_n316_));
  OAI21_X1  g115(.A(G204gat), .B1(new_n315_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(new_n313_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n317_), .A2(KEYINPUT92), .A3(new_n318_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n307_), .A2(new_n314_), .A3(new_n319_), .A4(KEYINPUT21), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n301_), .A2(new_n303_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT91), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n310_), .A2(new_n309_), .A3(new_n311_), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT21), .ZN(new_n325_));
  AOI21_X1  g124(.A(new_n325_), .B1(G197gat), .B2(G204gat), .ZN(new_n326_));
  AOI22_X1  g125(.A1(new_n323_), .A2(new_n304_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  OAI21_X1  g126(.A(new_n325_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n327_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n320_), .A2(new_n329_), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT89), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n299_), .A2(new_n330_), .A3(new_n331_), .ZN(new_n332_));
  XNOR2_X1  g131(.A(KEYINPUT88), .B(G233gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(G228gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G78gat), .B(G106gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n336_), .ZN(new_n338_));
  NAND4_X1  g137(.A1(new_n299_), .A2(new_n330_), .A3(new_n331_), .A4(new_n338_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n298_), .A2(new_n337_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT93), .ZN(new_n341_));
  INV_X1    g140(.A(new_n297_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n341_), .B1(new_n342_), .B2(new_n295_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n296_), .A2(KEYINPUT93), .A3(new_n297_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n337_), .A2(new_n339_), .ZN(new_n345_));
  NAND3_X1  g144(.A1(new_n343_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n340_), .A2(new_n346_), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n290_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT103), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT25), .ZN(new_n350_));
  NOR2_X1   g149(.A1(new_n350_), .A2(G183gat), .ZN(new_n351_));
  INV_X1    g150(.A(G183gat), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n352_), .A2(KEYINPUT25), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT94), .B1(new_n351_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(KEYINPUT26), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n355_), .A2(G190gat), .ZN(new_n356_));
  INV_X1    g155(.A(G190gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n357_), .A2(KEYINPUT26), .ZN(new_n358_));
  OAI21_X1  g157(.A(KEYINPUT95), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n352_), .A2(KEYINPUT25), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n350_), .A2(G183gat), .ZN(new_n361_));
  INV_X1    g160(.A(KEYINPUT94), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n360_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n357_), .A2(KEYINPUT26), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n355_), .A2(G190gat), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT95), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n364_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  NAND4_X1  g166(.A1(new_n354_), .A2(new_n359_), .A3(new_n363_), .A4(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT24), .ZN(new_n369_));
  INV_X1    g168(.A(G169gat), .ZN(new_n370_));
  INV_X1    g169(.A(G176gat), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n369_), .A2(new_n370_), .A3(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G183gat), .A2(G190gat), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT23), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n372_), .A2(new_n375_), .A3(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n370_), .A2(new_n371_), .A3(KEYINPUT81), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT81), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n379_), .B1(G169gat), .B2(G176gat), .ZN(new_n380_));
  AND2_X1   g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n369_), .B1(G169gat), .B2(G176gat), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n377_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n368_), .A2(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT22), .B(G169gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(new_n371_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n352_), .A2(new_n357_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n375_), .A2(new_n387_), .A3(new_n376_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(G169gat), .A2(G176gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n386_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n384_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n330_), .A2(new_n391_), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n375_), .A2(new_n376_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n393_), .B(new_n394_), .C1(new_n381_), .C2(KEYINPUT24), .ZN(new_n395_));
  AOI21_X1  g194(.A(KEYINPUT24), .B1(new_n378_), .B2(new_n380_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n375_), .A2(new_n376_), .ZN(new_n397_));
  OAI21_X1  g196(.A(KEYINPUT82), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NOR2_X1   g197(.A1(new_n351_), .A2(new_n353_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n364_), .A2(KEYINPUT80), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n356_), .A2(new_n358_), .ZN(new_n401_));
  OAI211_X1 g200(.A(new_n399_), .B(new_n400_), .C1(new_n401_), .C2(KEYINPUT80), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n381_), .A2(new_n382_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n395_), .A2(new_n398_), .A3(new_n402_), .A4(new_n403_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n394_), .A2(KEYINPUT84), .A3(new_n387_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT84), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n388_), .A2(new_n406_), .ZN(new_n407_));
  OR3_X1    g206(.A1(new_n370_), .A2(KEYINPUT83), .A3(KEYINPUT22), .ZN(new_n408_));
  OAI21_X1  g207(.A(KEYINPUT22), .B1(new_n370_), .B2(KEYINPUT83), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n408_), .A2(new_n371_), .A3(new_n409_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n405_), .A2(new_n407_), .A3(new_n389_), .A4(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n404_), .A2(new_n329_), .A3(new_n320_), .A4(new_n411_), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n392_), .A2(new_n412_), .A3(KEYINPUT20), .ZN(new_n413_));
  NAND2_X1  g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414_));
  XNOR2_X1  g213(.A(new_n414_), .B(KEYINPUT19), .ZN(new_n415_));
  NOR2_X1   g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(KEYINPUT20), .B1(new_n330_), .B2(new_n391_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT100), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n404_), .A2(new_n411_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(new_n330_), .ZN(new_n421_));
  OAI211_X1 g220(.A(KEYINPUT100), .B(KEYINPUT20), .C1(new_n330_), .C2(new_n391_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n419_), .A2(new_n421_), .A3(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n416_), .B1(new_n423_), .B2(new_n415_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G64gat), .B(G92gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n425_), .B(new_n426_), .ZN(new_n427_));
  XNOR2_X1  g226(.A(KEYINPUT96), .B(KEYINPUT18), .ZN(new_n428_));
  XNOR2_X1  g227(.A(new_n427_), .B(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n349_), .B1(new_n424_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n415_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n404_), .A2(new_n411_), .B1(new_n320_), .B2(new_n329_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT20), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n323_), .A2(KEYINPUT21), .A3(new_n304_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT92), .B1(new_n317_), .B2(new_n318_), .ZN(new_n436_));
  NOR2_X1   g235(.A1(new_n435_), .A2(new_n436_), .ZN(new_n437_));
  AOI22_X1  g236(.A1(new_n437_), .A2(new_n319_), .B1(new_n328_), .B2(new_n327_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n390_), .ZN(new_n439_));
  AOI21_X1  g238(.A(new_n439_), .B1(new_n368_), .B2(new_n383_), .ZN(new_n440_));
  AOI21_X1  g239(.A(new_n434_), .B1(new_n438_), .B2(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n433_), .B1(new_n441_), .B2(KEYINPUT100), .ZN(new_n442_));
  AOI21_X1  g241(.A(new_n432_), .B1(new_n442_), .B2(new_n419_), .ZN(new_n443_));
  OAI211_X1 g242(.A(KEYINPUT103), .B(new_n429_), .C1(new_n443_), .C2(new_n416_), .ZN(new_n444_));
  NOR3_X1   g243(.A1(new_n417_), .A2(new_n433_), .A3(new_n415_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n434_), .B1(new_n330_), .B2(new_n391_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n432_), .B1(new_n446_), .B2(new_n412_), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n445_), .A2(new_n447_), .A3(new_n429_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT27), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n431_), .A2(new_n444_), .A3(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n413_), .A2(new_n415_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n441_), .A2(new_n432_), .A3(new_n421_), .ZN(new_n453_));
  AOI21_X1  g252(.A(new_n430_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n449_), .B1(new_n448_), .B2(new_n454_), .ZN(new_n455_));
  AND2_X1   g254(.A1(new_n451_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n233_), .A2(new_n238_), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n457_), .B(KEYINPUT31), .ZN(new_n458_));
  XOR2_X1   g257(.A(G15gat), .B(G43gat), .Z(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n460_), .ZN(new_n461_));
  AND3_X1   g260(.A1(new_n404_), .A2(KEYINPUT30), .A3(new_n411_), .ZN(new_n462_));
  AOI21_X1  g261(.A(KEYINPUT30), .B1(new_n404_), .B2(new_n411_), .ZN(new_n463_));
  OAI21_X1  g262(.A(KEYINPUT85), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT30), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n420_), .A2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT85), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n404_), .A2(KEYINPUT30), .A3(new_n411_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(G227gat), .A2(G233gat), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  AND3_X1   g270(.A1(new_n464_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n471_), .B1(new_n464_), .B2(new_n469_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G71gat), .B(G99gat), .ZN(new_n474_));
  NOR3_X1   g273(.A1(new_n472_), .A2(new_n473_), .A3(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n474_), .ZN(new_n476_));
  NOR3_X1   g275(.A1(new_n462_), .A2(new_n463_), .A3(KEYINPUT85), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n467_), .B1(new_n466_), .B2(new_n468_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n470_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n464_), .A2(new_n469_), .A3(new_n471_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n476_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n461_), .B1(new_n475_), .B2(new_n481_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n474_), .B1(new_n472_), .B2(new_n473_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n479_), .A2(new_n476_), .A3(new_n480_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n484_), .A3(new_n460_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n482_), .A2(new_n485_), .ZN(new_n486_));
  AND3_X1   g285(.A1(new_n348_), .A2(new_n456_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n347_), .ZN(new_n488_));
  AND4_X1   g287(.A1(new_n488_), .A2(new_n285_), .A3(new_n455_), .A4(new_n289_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT33), .ZN(new_n490_));
  INV_X1    g289(.A(new_n202_), .ZN(new_n491_));
  AOI22_X1  g290(.A1(new_n282_), .A2(new_n491_), .B1(new_n276_), .B2(new_n272_), .ZN(new_n492_));
  OAI211_X1 g291(.A(new_n257_), .B(new_n202_), .C1(KEYINPUT4), .C2(new_n255_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n278_), .A2(new_n490_), .B1(new_n492_), .B2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n429_), .B1(new_n445_), .B2(new_n447_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n452_), .A2(new_n453_), .A3(new_n430_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n283_), .A2(KEYINPUT33), .A3(new_n277_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n494_), .A2(new_n495_), .A3(new_n496_), .A4(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n430_), .A2(KEYINPUT32), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n452_), .A2(new_n453_), .A3(new_n499_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n500_), .B1(new_n281_), .B2(new_n284_), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n423_), .A2(new_n415_), .ZN(new_n502_));
  INV_X1    g301(.A(new_n416_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n499_), .B1(new_n502_), .B2(new_n503_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n498_), .B1(new_n501_), .B2(new_n504_), .ZN(new_n505_));
  AOI22_X1  g304(.A1(new_n489_), .A2(new_n451_), .B1(new_n347_), .B2(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(KEYINPUT104), .B1(new_n506_), .B2(new_n486_), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT27), .B1(new_n495_), .B2(new_n496_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n508_), .A2(new_n347_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n290_), .A2(new_n451_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n505_), .A2(new_n347_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT104), .ZN(new_n513_));
  INV_X1    g312(.A(new_n486_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(new_n513_), .A3(new_n514_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n487_), .B1(new_n507_), .B2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G15gat), .B(G22gat), .ZN(new_n517_));
  INV_X1    g316(.A(G1gat), .ZN(new_n518_));
  INV_X1    g317(.A(G8gat), .ZN(new_n519_));
  OAI21_X1  g318(.A(KEYINPUT14), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  XOR2_X1   g320(.A(G1gat), .B(G8gat), .Z(new_n522_));
  XNOR2_X1  g321(.A(new_n521_), .B(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n523_), .B(KEYINPUT78), .ZN(new_n524_));
  NAND2_X1  g323(.A1(G231gat), .A2(G233gat), .ZN(new_n525_));
  XOR2_X1   g324(.A(new_n525_), .B(KEYINPUT79), .Z(new_n526_));
  XNOR2_X1  g325(.A(new_n524_), .B(new_n526_), .ZN(new_n527_));
  XOR2_X1   g326(.A(G71gat), .B(G78gat), .Z(new_n528_));
  XNOR2_X1  g327(.A(G57gat), .B(G64gat), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n528_), .B1(KEYINPUT11), .B2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n531_));
  XNOR2_X1  g330(.A(new_n530_), .B(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n527_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G127gat), .B(G155gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT16), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(G183gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n537_), .B(new_n302_), .ZN(new_n538_));
  OR3_X1    g337(.A1(new_n533_), .A2(new_n534_), .A3(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n538_), .B(KEYINPUT17), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n533_), .A2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  NOR2_X1   g341(.A1(new_n516_), .A2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT13), .ZN(new_n544_));
  XNOR2_X1  g343(.A(G120gat), .B(G148gat), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n545_), .B(G204gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(KEYINPUT5), .B(G176gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n546_), .B(new_n547_), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n548_), .B(KEYINPUT68), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT64), .B1(G85gat), .B2(G92gat), .ZN(new_n551_));
  INV_X1    g350(.A(KEYINPUT9), .ZN(new_n552_));
  INV_X1    g351(.A(G85gat), .ZN(new_n553_));
  INV_X1    g352(.A(G92gat), .ZN(new_n554_));
  OAI211_X1 g353(.A(new_n551_), .B(new_n552_), .C1(new_n553_), .C2(new_n554_), .ZN(new_n555_));
  AND2_X1   g354(.A1(G85gat), .A2(G92gat), .ZN(new_n556_));
  NOR2_X1   g355(.A1(G85gat), .A2(G92gat), .ZN(new_n557_));
  NOR3_X1   g356(.A1(new_n556_), .A2(new_n557_), .A3(KEYINPUT64), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n555_), .B1(new_n558_), .B2(new_n552_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G99gat), .A2(G106gat), .ZN(new_n560_));
  INV_X1    g359(.A(KEYINPUT6), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND3_X1  g361(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  INV_X1    g363(.A(G106gat), .ZN(new_n565_));
  AND2_X1   g364(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n566_));
  NOR2_X1   g365(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n567_));
  NOR2_X1   g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n564_), .B1(new_n565_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n559_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT7), .ZN(new_n571_));
  INV_X1    g370(.A(G99gat), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(new_n572_), .A3(new_n565_), .ZN(new_n573_));
  OAI21_X1  g372(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n574_));
  NAND4_X1  g373(.A1(new_n573_), .A2(new_n562_), .A3(new_n563_), .A4(new_n574_), .ZN(new_n575_));
  NOR2_X1   g374(.A1(new_n556_), .A2(new_n557_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n575_), .A2(new_n576_), .ZN(new_n577_));
  INV_X1    g376(.A(KEYINPUT8), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n577_), .A2(new_n578_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n575_), .A2(KEYINPUT8), .A3(new_n576_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n570_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n529_), .A2(KEYINPUT11), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n530_), .B(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(KEYINPUT66), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n570_), .A2(new_n579_), .A3(new_n580_), .ZN(new_n586_));
  INV_X1    g385(.A(KEYINPUT65), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n586_), .A2(new_n587_), .A3(new_n532_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT66), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n581_), .A2(new_n583_), .A3(new_n589_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT65), .B1(new_n581_), .B2(new_n583_), .ZN(new_n591_));
  NAND4_X1  g390(.A1(new_n585_), .A2(new_n588_), .A3(new_n590_), .A4(new_n591_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n592_), .A2(G230gat), .A3(G233gat), .ZN(new_n593_));
  OAI21_X1  g392(.A(KEYINPUT12), .B1(new_n581_), .B2(new_n583_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n594_), .A2(new_n584_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT67), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n581_), .A2(new_n596_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n570_), .A2(new_n579_), .A3(KEYINPUT67), .A4(new_n580_), .ZN(new_n598_));
  NAND4_X1  g397(.A1(new_n597_), .A2(KEYINPUT12), .A3(new_n583_), .A4(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G230gat), .A2(G233gat), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n595_), .A2(new_n599_), .A3(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n550_), .B1(new_n593_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT69), .ZN(new_n603_));
  INV_X1    g402(.A(new_n603_), .ZN(new_n604_));
  NAND3_X1  g403(.A1(new_n593_), .A2(new_n601_), .A3(new_n548_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n605_), .B1(new_n602_), .B2(KEYINPUT69), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n544_), .B1(new_n604_), .B2(new_n606_), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n602_), .A2(KEYINPUT69), .ZN(new_n608_));
  NAND4_X1  g407(.A1(new_n608_), .A2(KEYINPUT13), .A3(new_n603_), .A4(new_n605_), .ZN(new_n609_));
  AND2_X1   g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n610_), .A2(KEYINPUT70), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n607_), .A2(new_n609_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT70), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n612_), .A2(new_n613_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(G113gat), .B(G141gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(G169gat), .ZN(new_n617_));
  INV_X1    g416(.A(G197gat), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT15), .ZN(new_n621_));
  XOR2_X1   g420(.A(G29gat), .B(G36gat), .Z(new_n622_));
  XNOR2_X1  g421(.A(G43gat), .B(G50gat), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  XOR2_X1   g423(.A(G43gat), .B(G50gat), .Z(new_n625_));
  XNOR2_X1  g424(.A(G29gat), .B(G36gat), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n625_), .A2(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(KEYINPUT71), .B(KEYINPUT72), .ZN(new_n628_));
  AND3_X1   g427(.A1(new_n624_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n628_), .B1(new_n624_), .B2(new_n627_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n621_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n624_), .A2(new_n627_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n628_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n624_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n634_), .A2(KEYINPUT15), .A3(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n631_), .A2(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n521_), .B(new_n522_), .Z(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(new_n639_));
  NOR2_X1   g438(.A1(new_n629_), .A2(new_n630_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n523_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(G229gat), .A2(G233gat), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n639_), .A2(new_n641_), .A3(new_n642_), .ZN(new_n643_));
  OAI21_X1  g442(.A(new_n638_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n642_), .B1(new_n641_), .B2(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n620_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n646_));
  AND2_X1   g445(.A1(new_n641_), .A2(new_n642_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n645_), .B1(new_n639_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(new_n619_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n646_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n615_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT36), .ZN(new_n653_));
  XNOR2_X1  g452(.A(G134gat), .B(G162gat), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT73), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(new_n357_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n657_), .A2(new_n300_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n656_), .B(G190gat), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n659_), .A2(G218gat), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n653_), .B1(new_n658_), .B2(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n659_), .A2(G218gat), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n657_), .A2(new_n300_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n662_), .A2(new_n663_), .A3(KEYINPUT36), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n661_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT76), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n665_), .A2(new_n666_), .ZN(new_n667_));
  NAND3_X1  g466(.A1(new_n661_), .A2(KEYINPUT76), .A3(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n637_), .A2(new_n597_), .A3(new_n598_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n586_), .A2(new_n640_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(G232gat), .A2(G233gat), .ZN(new_n672_));
  XOR2_X1   g471(.A(new_n672_), .B(KEYINPUT34), .Z(new_n673_));
  INV_X1    g472(.A(KEYINPUT35), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n675_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(KEYINPUT74), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n676_), .A2(KEYINPUT74), .ZN(new_n678_));
  AND2_X1   g477(.A1(new_n673_), .A2(new_n674_), .ZN(new_n679_));
  NOR3_X1   g478(.A1(new_n677_), .A2(new_n678_), .A3(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n670_), .A2(new_n671_), .A3(new_n680_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT75), .ZN(new_n682_));
  OR2_X1    g481(.A1(new_n681_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n670_), .A2(new_n671_), .ZN(new_n684_));
  AOI22_X1  g483(.A1(new_n681_), .A2(new_n682_), .B1(new_n684_), .B2(new_n675_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n669_), .B1(new_n683_), .B2(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(new_n661_), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n685_), .A2(new_n683_), .A3(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT37), .B1(new_n686_), .B2(new_n689_), .ZN(new_n690_));
  INV_X1    g489(.A(KEYINPUT77), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n665_), .B1(new_n685_), .B2(new_n683_), .ZN(new_n692_));
  NOR2_X1   g491(.A1(new_n689_), .A2(new_n692_), .ZN(new_n693_));
  INV_X1    g492(.A(KEYINPUT37), .ZN(new_n694_));
  AOI22_X1  g493(.A1(new_n690_), .A2(new_n691_), .B1(new_n693_), .B2(new_n694_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n685_), .A2(new_n683_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n696_), .A2(new_n667_), .A3(new_n668_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n694_), .B1(new_n697_), .B2(new_n688_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT77), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n695_), .A2(new_n699_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n543_), .A2(new_n652_), .A3(new_n700_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT105), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND4_X1  g502(.A1(new_n543_), .A2(new_n652_), .A3(KEYINPUT105), .A4(new_n700_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT38), .ZN(new_n706_));
  INV_X1    g505(.A(new_n290_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n518_), .ZN(new_n708_));
  OR3_X1    g507(.A1(new_n705_), .A2(new_n706_), .A3(new_n708_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n348_), .A2(new_n456_), .A3(new_n486_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n513_), .B1(new_n512_), .B2(new_n514_), .ZN(new_n711_));
  AOI211_X1 g510(.A(KEYINPUT104), .B(new_n486_), .C1(new_n510_), .C2(new_n511_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n710_), .B1(new_n711_), .B2(new_n712_), .ZN(new_n713_));
  NAND3_X1  g512(.A1(new_n607_), .A2(new_n609_), .A3(new_n650_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT106), .ZN(new_n715_));
  INV_X1    g514(.A(new_n542_), .ZN(new_n716_));
  INV_X1    g515(.A(new_n692_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n688_), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n713_), .A2(new_n715_), .A3(new_n716_), .A4(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G1gat), .B1(new_n719_), .B2(new_n290_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n706_), .B1(new_n705_), .B2(new_n708_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n709_), .A2(new_n720_), .A3(new_n721_), .ZN(G1324gat));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n723_));
  INV_X1    g522(.A(new_n456_), .ZN(new_n724_));
  NAND4_X1  g523(.A1(new_n703_), .A2(new_n704_), .A3(new_n519_), .A4(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G8gat), .B1(new_n719_), .B2(new_n456_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT39), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT39), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n728_), .B(G8gat), .C1(new_n719_), .C2(new_n456_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  AOI21_X1  g529(.A(new_n723_), .B1(new_n725_), .B2(new_n730_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n731_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n725_), .A2(new_n730_), .A3(new_n723_), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n732_), .A2(KEYINPUT40), .A3(new_n733_), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT40), .ZN(new_n735_));
  INV_X1    g534(.A(new_n733_), .ZN(new_n736_));
  OAI21_X1  g535(.A(new_n735_), .B1(new_n736_), .B2(new_n731_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n737_), .ZN(G1325gat));
  NOR3_X1   g537(.A1(new_n516_), .A2(new_n542_), .A3(new_n693_), .ZN(new_n739_));
  NAND3_X1  g538(.A1(new_n739_), .A2(new_n486_), .A3(new_n715_), .ZN(new_n740_));
  NAND3_X1  g539(.A1(new_n740_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n741_));
  INV_X1    g540(.A(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(KEYINPUT41), .B1(new_n740_), .B2(G15gat), .ZN(new_n743_));
  OR2_X1    g542(.A1(new_n514_), .A2(G15gat), .ZN(new_n744_));
  OAI22_X1  g543(.A1(new_n742_), .A2(new_n743_), .B1(new_n705_), .B2(new_n744_), .ZN(new_n745_));
  XOR2_X1   g544(.A(new_n745_), .B(KEYINPUT108), .Z(G1326gat));
  OR3_X1    g545(.A1(new_n705_), .A2(G22gat), .A3(new_n347_), .ZN(new_n747_));
  OAI21_X1  g546(.A(G22gat), .B1(new_n719_), .B2(new_n347_), .ZN(new_n748_));
  OR2_X1    g547(.A1(new_n748_), .A2(KEYINPUT109), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n748_), .A2(KEYINPUT109), .ZN(new_n750_));
  AND3_X1   g549(.A1(new_n749_), .A2(KEYINPUT42), .A3(new_n750_), .ZN(new_n751_));
  AOI21_X1  g550(.A(KEYINPUT42), .B1(new_n749_), .B2(new_n750_), .ZN(new_n752_));
  OAI21_X1  g551(.A(new_n747_), .B1(new_n751_), .B2(new_n752_), .ZN(G1327gat));
  NOR3_X1   g552(.A1(new_n516_), .A2(new_n716_), .A3(new_n718_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n714_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n754_), .A2(new_n755_), .ZN(new_n756_));
  AOI21_X1  g555(.A(G29gat), .B1(new_n756_), .B2(new_n707_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n715_), .A2(new_n542_), .ZN(new_n758_));
  INV_X1    g557(.A(new_n758_), .ZN(new_n759_));
  NOR3_X1   g558(.A1(new_n516_), .A2(KEYINPUT43), .A3(new_n700_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n761_));
  OAI22_X1  g560(.A1(new_n698_), .A2(KEYINPUT77), .B1(new_n718_), .B2(KEYINPUT37), .ZN(new_n762_));
  NOR2_X1   g561(.A1(new_n690_), .A2(new_n691_), .ZN(new_n763_));
  NOR2_X1   g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n761_), .B1(new_n713_), .B2(new_n764_), .ZN(new_n765_));
  OAI211_X1 g564(.A(KEYINPUT44), .B(new_n759_), .C1(new_n760_), .C2(new_n765_), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n766_), .A2(G29gat), .A3(new_n707_), .ZN(new_n767_));
  OAI21_X1  g566(.A(new_n759_), .B1(new_n760_), .B2(new_n765_), .ZN(new_n768_));
  XOR2_X1   g567(.A(KEYINPUT110), .B(KEYINPUT44), .Z(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n757_), .B1(new_n767_), .B2(new_n771_), .ZN(G1328gat));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n766_), .A2(new_n724_), .ZN(new_n774_));
  OAI21_X1  g573(.A(KEYINPUT43), .B1(new_n516_), .B2(new_n700_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n713_), .A2(new_n761_), .A3(new_n764_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n758_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n777_), .A2(new_n769_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n773_), .B1(new_n774_), .B2(new_n778_), .ZN(new_n779_));
  NAND4_X1  g578(.A1(new_n771_), .A2(KEYINPUT111), .A3(new_n724_), .A4(new_n766_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n779_), .A2(G36gat), .A3(new_n780_), .ZN(new_n781_));
  XOR2_X1   g580(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(new_n756_), .ZN(new_n784_));
  INV_X1    g583(.A(G36gat), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n724_), .A2(new_n785_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n783_), .B1(new_n784_), .B2(new_n786_), .ZN(new_n787_));
  NAND4_X1  g586(.A1(new_n756_), .A2(new_n785_), .A3(new_n724_), .A4(new_n782_), .ZN(new_n788_));
  AND2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n781_), .A2(KEYINPUT46), .A3(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n787_), .A2(new_n788_), .ZN(new_n791_));
  OAI211_X1 g590(.A(new_n766_), .B(new_n724_), .C1(new_n777_), .C2(new_n769_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n785_), .B1(new_n792_), .B2(new_n773_), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n791_), .B1(new_n793_), .B2(new_n780_), .ZN(new_n794_));
  XOR2_X1   g593(.A(KEYINPUT113), .B(KEYINPUT46), .Z(new_n795_));
  OAI21_X1  g594(.A(new_n790_), .B1(new_n794_), .B2(new_n795_), .ZN(G1329gat));
  INV_X1    g595(.A(G43gat), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n797_), .B1(new_n784_), .B2(new_n514_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n766_), .A2(G43gat), .A3(new_n486_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n798_), .B1(new_n799_), .B2(new_n778_), .ZN(new_n800_));
  XNOR2_X1  g599(.A(new_n800_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g600(.A(G50gat), .B1(new_n756_), .B2(new_n488_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n766_), .A2(G50gat), .A3(new_n488_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(new_n771_), .ZN(G1331gat));
  INV_X1    g603(.A(new_n615_), .ZN(new_n805_));
  NOR2_X1   g604(.A1(new_n805_), .A2(new_n650_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(new_n739_), .ZN(new_n807_));
  OAI21_X1  g606(.A(G57gat), .B1(new_n807_), .B2(new_n290_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n610_), .A2(new_n650_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n543_), .A2(new_n700_), .A3(new_n809_), .ZN(new_n810_));
  OR2_X1    g609(.A1(new_n290_), .A2(G57gat), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n808_), .B1(new_n810_), .B2(new_n811_), .ZN(G1332gat));
  OAI21_X1  g611(.A(G64gat), .B1(new_n807_), .B2(new_n456_), .ZN(new_n813_));
  XNOR2_X1  g612(.A(new_n813_), .B(KEYINPUT48), .ZN(new_n814_));
  OR2_X1    g613(.A1(new_n456_), .A2(G64gat), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n814_), .B1(new_n810_), .B2(new_n815_), .ZN(G1333gat));
  OAI21_X1  g615(.A(G71gat), .B1(new_n807_), .B2(new_n514_), .ZN(new_n817_));
  XNOR2_X1  g616(.A(new_n817_), .B(KEYINPUT49), .ZN(new_n818_));
  OR2_X1    g617(.A1(new_n514_), .A2(G71gat), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n818_), .B1(new_n810_), .B2(new_n819_), .ZN(G1334gat));
  OAI21_X1  g619(.A(G78gat), .B1(new_n807_), .B2(new_n347_), .ZN(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT50), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n347_), .A2(G78gat), .ZN(new_n823_));
  OAI21_X1  g622(.A(new_n822_), .B1(new_n810_), .B2(new_n823_), .ZN(G1335gat));
  OAI211_X1 g623(.A(new_n542_), .B(new_n809_), .C1(new_n760_), .C2(new_n765_), .ZN(new_n825_));
  OAI21_X1  g624(.A(G85gat), .B1(new_n825_), .B2(new_n290_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n806_), .A2(new_n754_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n827_), .A2(new_n553_), .A3(new_n707_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1336gat));
  OAI21_X1  g628(.A(G92gat), .B1(new_n825_), .B2(new_n456_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(new_n554_), .A3(new_n724_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1337gat));
  OAI21_X1  g631(.A(G99gat), .B1(new_n825_), .B2(new_n514_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT114), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n827_), .A2(new_n486_), .A3(new_n568_), .ZN(new_n835_));
  AND3_X1   g634(.A1(new_n833_), .A2(new_n834_), .A3(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n836_), .B(new_n837_), .ZN(G1338gat));
  NAND3_X1  g637(.A1(new_n827_), .A2(new_n565_), .A3(new_n488_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT52), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n809_), .A2(new_n542_), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n488_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n840_), .B1(new_n843_), .B2(G106gat), .ZN(new_n844_));
  AOI211_X1 g643(.A(KEYINPUT52), .B(new_n565_), .C1(new_n842_), .C2(new_n488_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n839_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  XNOR2_X1  g645(.A(new_n846_), .B(KEYINPUT53), .ZN(G1339gat));
  AOI21_X1  g646(.A(new_n600_), .B1(new_n595_), .B2(new_n599_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n601_), .B1(new_n848_), .B2(new_n849_), .ZN(new_n850_));
  NAND4_X1  g649(.A1(new_n595_), .A2(new_n599_), .A3(KEYINPUT55), .A4(new_n600_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  AOI21_X1  g651(.A(KEYINPUT56), .B1(new_n852_), .B2(new_n549_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854_));
  AOI211_X1 g653(.A(new_n854_), .B(new_n550_), .C1(new_n850_), .C2(new_n851_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n639_), .A2(G229gat), .A3(G233gat), .A4(new_n641_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n641_), .A2(new_n644_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n619_), .B1(new_n857_), .B2(new_n642_), .ZN(new_n858_));
  AOI22_X1  g657(.A1(new_n648_), .A2(new_n619_), .B1(new_n856_), .B2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n605_), .A2(new_n859_), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(new_n860_), .B1(new_n605_), .B2(new_n859_), .ZN(new_n862_));
  OAI22_X1  g661(.A1(new_n853_), .A2(new_n855_), .B1(new_n861_), .B2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT58), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n863_), .A2(new_n864_), .ZN(new_n865_));
  OAI221_X1 g664(.A(KEYINPUT58), .B1(new_n861_), .B2(new_n862_), .C1(new_n853_), .C2(new_n855_), .ZN(new_n866_));
  NAND4_X1  g665(.A1(new_n695_), .A2(new_n699_), .A3(new_n865_), .A4(new_n866_), .ZN(new_n867_));
  AND2_X1   g666(.A1(new_n650_), .A2(new_n605_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n868_), .B1(new_n853_), .B2(new_n855_), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT115), .ZN(new_n870_));
  NAND3_X1  g669(.A1(new_n608_), .A2(new_n603_), .A3(new_n605_), .ZN(new_n871_));
  AOI22_X1  g670(.A1(new_n869_), .A2(new_n870_), .B1(new_n871_), .B2(new_n859_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n868_), .B(KEYINPUT115), .C1(new_n853_), .C2(new_n855_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n693_), .B1(new_n872_), .B2(new_n873_), .ZN(new_n874_));
  OAI21_X1  g673(.A(new_n867_), .B1(new_n874_), .B2(KEYINPUT57), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876_));
  AOI211_X1 g675(.A(new_n876_), .B(new_n693_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n542_), .B1(new_n875_), .B2(new_n877_), .ZN(new_n878_));
  NOR3_X1   g677(.A1(new_n612_), .A2(new_n542_), .A3(new_n650_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n700_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n880_), .A2(KEYINPUT54), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n700_), .A2(new_n879_), .A3(new_n882_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n881_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n878_), .A2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n724_), .A2(new_n290_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n887_), .A2(new_n514_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n885_), .A2(new_n347_), .A3(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(KEYINPUT59), .ZN(new_n890_));
  AOI21_X1  g689(.A(new_n488_), .B1(new_n878_), .B2(new_n884_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n891_), .A2(new_n892_), .A3(new_n888_), .ZN(new_n893_));
  XNOR2_X1  g692(.A(KEYINPUT118), .B(G113gat), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n651_), .A2(new_n894_), .ZN(new_n895_));
  XNOR2_X1  g694(.A(new_n895_), .B(KEYINPUT119), .ZN(new_n896_));
  NAND3_X1  g695(.A1(new_n890_), .A2(new_n893_), .A3(new_n896_), .ZN(new_n897_));
  NAND4_X1  g696(.A1(new_n885_), .A2(new_n347_), .A3(new_n650_), .A4(new_n888_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n899_));
  AND3_X1   g698(.A1(new_n898_), .A2(new_n899_), .A3(new_n228_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(new_n228_), .ZN(new_n901_));
  OAI21_X1  g700(.A(new_n897_), .B1(new_n900_), .B2(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n902_), .A2(new_n903_), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n897_), .B(KEYINPUT120), .C1(new_n900_), .C2(new_n901_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n904_), .A2(new_n905_), .ZN(G1340gat));
  INV_X1    g705(.A(new_n889_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT60), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n610_), .B2(G120gat), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n907_), .A2(new_n908_), .A3(new_n909_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n805_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n911_));
  AND3_X1   g710(.A1(new_n911_), .A2(new_n890_), .A3(new_n893_), .ZN(new_n912_));
  OAI21_X1  g711(.A(new_n910_), .B1(new_n912_), .B2(new_n226_), .ZN(G1341gat));
  NAND3_X1  g712(.A1(new_n890_), .A2(new_n716_), .A3(new_n893_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n914_), .A2(G127gat), .ZN(new_n915_));
  OR2_X1    g714(.A1(new_n542_), .A2(G127gat), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n915_), .B1(new_n889_), .B2(new_n916_), .ZN(G1342gat));
  NAND3_X1  g716(.A1(new_n890_), .A2(new_n764_), .A3(new_n893_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n918_), .A2(G134gat), .ZN(new_n919_));
  OR2_X1    g718(.A1(new_n718_), .A2(G134gat), .ZN(new_n920_));
  OAI21_X1  g719(.A(new_n919_), .B1(new_n889_), .B2(new_n920_), .ZN(G1343gat));
  NOR2_X1   g720(.A1(new_n486_), .A2(new_n347_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n869_), .A2(new_n870_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n871_), .A2(new_n859_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n923_), .A2(new_n873_), .A3(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(new_n718_), .ZN(new_n926_));
  AND2_X1   g725(.A1(new_n865_), .A2(new_n866_), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n926_), .A2(new_n876_), .B1(new_n764_), .B2(new_n927_), .ZN(new_n928_));
  INV_X1    g727(.A(new_n877_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n716_), .B1(new_n928_), .B2(new_n929_), .ZN(new_n930_));
  INV_X1    g729(.A(new_n883_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n882_), .B1(new_n700_), .B2(new_n879_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n931_), .A2(new_n932_), .ZN(new_n933_));
  OAI211_X1 g732(.A(new_n886_), .B(new_n922_), .C1(new_n930_), .C2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n934_), .A2(new_n651_), .ZN(new_n935_));
  XOR2_X1   g734(.A(KEYINPUT121), .B(G141gat), .Z(new_n936_));
  XNOR2_X1  g735(.A(new_n935_), .B(new_n936_), .ZN(G1344gat));
  NOR2_X1   g736(.A1(new_n934_), .A2(new_n805_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(new_n212_), .ZN(G1345gat));
  XNOR2_X1  g738(.A(KEYINPUT61), .B(G155gat), .ZN(new_n940_));
  INV_X1    g739(.A(new_n940_), .ZN(new_n941_));
  OAI21_X1  g740(.A(KEYINPUT122), .B1(new_n934_), .B2(new_n542_), .ZN(new_n942_));
  INV_X1    g741(.A(KEYINPUT123), .ZN(new_n943_));
  INV_X1    g742(.A(new_n922_), .ZN(new_n944_));
  AOI21_X1  g743(.A(new_n944_), .B1(new_n878_), .B2(new_n884_), .ZN(new_n945_));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n945_), .A2(new_n946_), .A3(new_n716_), .A4(new_n886_), .ZN(new_n947_));
  AND3_X1   g746(.A1(new_n942_), .A2(new_n943_), .A3(new_n947_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n943_), .B1(new_n942_), .B2(new_n947_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n941_), .B1(new_n948_), .B2(new_n949_), .ZN(new_n950_));
  AOI211_X1 g749(.A(new_n887_), .B(new_n944_), .C1(new_n878_), .C2(new_n884_), .ZN(new_n951_));
  AOI21_X1  g750(.A(new_n946_), .B1(new_n951_), .B2(new_n716_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n947_), .ZN(new_n953_));
  OAI21_X1  g752(.A(KEYINPUT123), .B1(new_n952_), .B2(new_n953_), .ZN(new_n954_));
  NAND3_X1  g753(.A1(new_n942_), .A2(new_n943_), .A3(new_n947_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n954_), .A2(new_n940_), .A3(new_n955_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n950_), .A2(new_n956_), .ZN(G1346gat));
  INV_X1    g756(.A(G162gat), .ZN(new_n958_));
  NOR3_X1   g757(.A1(new_n934_), .A2(new_n958_), .A3(new_n700_), .ZN(new_n959_));
  OAI21_X1  g758(.A(new_n958_), .B1(new_n934_), .B2(new_n718_), .ZN(new_n960_));
  OR2_X1    g759(.A1(new_n960_), .A2(KEYINPUT124), .ZN(new_n961_));
  NAND2_X1  g760(.A1(new_n960_), .A2(KEYINPUT124), .ZN(new_n962_));
  AOI21_X1  g761(.A(new_n959_), .B1(new_n961_), .B2(new_n962_), .ZN(G1347gat));
  NOR3_X1   g762(.A1(new_n456_), .A2(new_n514_), .A3(new_n707_), .ZN(new_n964_));
  NAND2_X1  g763(.A1(new_n891_), .A2(new_n964_), .ZN(new_n965_));
  OAI21_X1  g764(.A(G169gat), .B1(new_n965_), .B2(new_n651_), .ZN(new_n966_));
  INV_X1    g765(.A(KEYINPUT62), .ZN(new_n967_));
  OR2_X1    g766(.A1(new_n966_), .A2(new_n967_), .ZN(new_n968_));
  INV_X1    g767(.A(new_n965_), .ZN(new_n969_));
  NAND3_X1  g768(.A1(new_n969_), .A2(new_n385_), .A3(new_n650_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(new_n966_), .A2(new_n967_), .ZN(new_n971_));
  NAND3_X1  g770(.A1(new_n968_), .A2(new_n970_), .A3(new_n971_), .ZN(G1348gat));
  NOR3_X1   g771(.A1(new_n965_), .A2(new_n371_), .A3(new_n805_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n969_), .A2(new_n612_), .ZN(new_n974_));
  AOI21_X1  g773(.A(new_n973_), .B1(new_n371_), .B2(new_n974_), .ZN(G1349gat));
  NAND2_X1  g774(.A1(new_n969_), .A2(new_n716_), .ZN(new_n976_));
  AOI21_X1  g775(.A(new_n976_), .B1(new_n354_), .B2(new_n363_), .ZN(new_n977_));
  AOI21_X1  g776(.A(new_n977_), .B1(new_n352_), .B2(new_n976_), .ZN(G1350gat));
  OAI21_X1  g777(.A(G190gat), .B1(new_n965_), .B2(new_n700_), .ZN(new_n979_));
  NAND3_X1  g778(.A1(new_n693_), .A2(new_n359_), .A3(new_n367_), .ZN(new_n980_));
  OAI21_X1  g779(.A(new_n979_), .B1(new_n965_), .B2(new_n980_), .ZN(G1351gat));
  NOR2_X1   g780(.A1(new_n456_), .A2(new_n707_), .ZN(new_n982_));
  AND2_X1   g781(.A1(new_n945_), .A2(new_n982_), .ZN(new_n983_));
  NAND2_X1  g782(.A1(new_n983_), .A2(new_n650_), .ZN(new_n984_));
  XNOR2_X1  g783(.A(new_n984_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g784(.A1(KEYINPUT125), .A2(G204gat), .ZN(new_n986_));
  XNOR2_X1  g785(.A(KEYINPUT125), .B(G204gat), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n983_), .A2(new_n615_), .ZN(new_n988_));
  MUX2_X1   g787(.A(new_n986_), .B(new_n987_), .S(new_n988_), .Z(G1353gat));
  NAND2_X1  g788(.A1(new_n983_), .A2(new_n716_), .ZN(new_n990_));
  NOR2_X1   g789(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n991_));
  AND2_X1   g790(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n992_));
  NOR3_X1   g791(.A1(new_n990_), .A2(new_n991_), .A3(new_n992_), .ZN(new_n993_));
  AOI21_X1  g792(.A(new_n993_), .B1(new_n990_), .B2(new_n991_), .ZN(G1354gat));
  NAND4_X1  g793(.A1(new_n885_), .A2(new_n693_), .A3(new_n922_), .A4(new_n982_), .ZN(new_n995_));
  NAND2_X1  g794(.A1(new_n995_), .A2(KEYINPUT126), .ZN(new_n996_));
  INV_X1    g795(.A(KEYINPUT126), .ZN(new_n997_));
  NAND4_X1  g796(.A1(new_n945_), .A2(new_n997_), .A3(new_n693_), .A4(new_n982_), .ZN(new_n998_));
  NAND3_X1  g797(.A1(new_n996_), .A2(new_n300_), .A3(new_n998_), .ZN(new_n999_));
  NAND3_X1  g798(.A1(new_n983_), .A2(G218gat), .A3(new_n764_), .ZN(new_n1000_));
  NAND2_X1  g799(.A1(new_n999_), .A2(new_n1000_), .ZN(new_n1001_));
  NAND2_X1  g800(.A1(new_n1001_), .A2(KEYINPUT127), .ZN(new_n1002_));
  INV_X1    g801(.A(KEYINPUT127), .ZN(new_n1003_));
  NAND3_X1  g802(.A1(new_n999_), .A2(new_n1003_), .A3(new_n1000_), .ZN(new_n1004_));
  NAND2_X1  g803(.A1(new_n1002_), .A2(new_n1004_), .ZN(G1355gat));
endmodule


