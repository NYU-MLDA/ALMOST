//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n801_,
    new_n802_, new_n803_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n846_, new_n847_, new_n849_, new_n850_, new_n851_,
    new_n853_, new_n854_, new_n855_, new_n856_, new_n857_, new_n858_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n938_, new_n939_, new_n940_,
    new_n942_, new_n943_, new_n944_, new_n945_, new_n946_, new_n947_,
    new_n948_, new_n949_, new_n950_, new_n952_, new_n953_, new_n955_,
    new_n956_, new_n957_, new_n958_, new_n960_, new_n961_, new_n962_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n995_,
    new_n996_, new_n998_, new_n999_, new_n1000_, new_n1002_, new_n1003_,
    new_n1004_, new_n1005_, new_n1006_, new_n1007_, new_n1009_, new_n1011_,
    new_n1012_, new_n1013_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_;
  XOR2_X1   g000(.A(KEYINPUT86), .B(KEYINPUT31), .Z(new_n202_));
  NAND2_X1  g001(.A1(G227gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G15gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT84), .ZN(new_n205_));
  INV_X1    g004(.A(G15gat), .ZN(new_n206_));
  XNOR2_X1  g005(.A(new_n203_), .B(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT84), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n205_), .A2(new_n209_), .ZN(new_n210_));
  XNOR2_X1  g009(.A(G71gat), .B(G99gat), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(G43gat), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G43gat), .ZN(new_n214_));
  XNOR2_X1  g013(.A(new_n211_), .B(new_n214_), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n215_), .A2(new_n205_), .A3(new_n209_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219_));
  INV_X1    g018(.A(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G169gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n221_), .A2(KEYINPUT22), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT22), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(G169gat), .ZN(new_n224_));
  INV_X1    g023(.A(G176gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n222_), .A2(new_n224_), .A3(new_n225_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT82), .ZN(new_n227_));
  XNOR2_X1  g026(.A(KEYINPUT22), .B(G169gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT82), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(new_n229_), .A3(new_n225_), .ZN(new_n230_));
  AOI21_X1  g029(.A(new_n220_), .B1(new_n227_), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT23), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(G183gat), .A3(G190gat), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT83), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT23), .ZN(new_n237_));
  NAND4_X1  g036(.A1(new_n232_), .A2(KEYINPUT83), .A3(G183gat), .A4(G190gat), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n235_), .A2(new_n237_), .A3(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(G183gat), .ZN(new_n240_));
  INV_X1    g039(.A(G190gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n239_), .A2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n231_), .A2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n240_), .A2(KEYINPUT25), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(G183gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n241_), .A2(KEYINPUT26), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT26), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(G190gat), .ZN(new_n250_));
  AND4_X1   g049(.A1(new_n245_), .A2(new_n247_), .A3(new_n248_), .A4(new_n250_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(G169gat), .A2(G176gat), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT24), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n252_), .A2(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n219_), .A2(KEYINPUT24), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n254_), .B1(new_n255_), .B2(new_n252_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n251_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT81), .ZN(new_n258_));
  AOI22_X1  g057(.A1(new_n233_), .A2(new_n258_), .B1(KEYINPUT23), .B2(new_n236_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n240_), .A2(KEYINPUT23), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n260_), .A2(KEYINPUT81), .A3(G190gat), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n259_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n257_), .A2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n244_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT30), .ZN(new_n265_));
  NOR2_X1   g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  AOI22_X1  g065(.A1(new_n231_), .A2(new_n243_), .B1(new_n257_), .B2(new_n262_), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n267_), .A2(KEYINPUT30), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n218_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G127gat), .B(G134gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(G113gat), .B(G120gat), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT85), .ZN(new_n272_));
  OR3_X1    g071(.A1(new_n270_), .A2(new_n271_), .A3(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n272_), .B1(new_n270_), .B2(new_n271_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n270_), .A2(new_n271_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n273_), .A2(new_n274_), .A3(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n264_), .A2(new_n265_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n267_), .A2(KEYINPUT30), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n277_), .A2(new_n278_), .A3(new_n217_), .ZN(new_n279_));
  AND3_X1   g078(.A1(new_n269_), .A2(new_n276_), .A3(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n276_), .B1(new_n269_), .B2(new_n279_), .ZN(new_n281_));
  OAI21_X1  g080(.A(new_n202_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n276_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n279_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n217_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n283_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n269_), .A2(new_n276_), .A3(new_n279_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n202_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n286_), .A2(new_n287_), .A3(new_n288_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n282_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(G155gat), .A2(G162gat), .ZN(new_n293_));
  NOR2_X1   g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n294_), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT87), .ZN(new_n296_));
  INV_X1    g095(.A(KEYINPUT3), .ZN(new_n297_));
  INV_X1    g096(.A(G141gat), .ZN(new_n298_));
  INV_X1    g097(.A(G148gat), .ZN(new_n299_));
  NAND4_X1  g098(.A1(new_n296_), .A2(new_n297_), .A3(new_n298_), .A4(new_n299_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(KEYINPUT87), .A2(KEYINPUT3), .ZN(new_n301_));
  OAI22_X1  g100(.A1(KEYINPUT87), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G141gat), .A2(G148gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT2), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  AND4_X1   g104(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .A4(new_n305_), .ZN(new_n306_));
  NAND3_X1  g105(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT88), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  AOI21_X1  g108(.A(new_n295_), .B1(new_n306_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n298_), .A2(new_n299_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n311_), .A2(new_n303_), .ZN(new_n312_));
  INV_X1    g111(.A(KEYINPUT1), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n292_), .A2(new_n313_), .ZN(new_n314_));
  OAI21_X1  g113(.A(new_n291_), .B1(new_n293_), .B2(KEYINPUT1), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n312_), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  OAI21_X1  g115(.A(KEYINPUT29), .B1(new_n310_), .B2(new_n316_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT92), .ZN(new_n318_));
  INV_X1    g117(.A(G218gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n319_), .A2(G211gat), .ZN(new_n320_));
  INV_X1    g119(.A(G211gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n321_), .A2(G218gat), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(G197gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n324_), .A2(KEYINPUT90), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT90), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n326_), .A2(G197gat), .ZN(new_n327_));
  INV_X1    g126(.A(G204gat), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n325_), .A2(new_n327_), .A3(new_n328_), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT21), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n330_), .B1(G197gat), .B2(G204gat), .ZN(new_n331_));
  AOI21_X1  g130(.A(new_n323_), .B1(new_n329_), .B2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n325_), .A2(new_n327_), .A3(G204gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n328_), .A2(G197gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(KEYINPUT91), .B(KEYINPUT21), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n333_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n332_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n333_), .A2(new_n334_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n330_), .B1(new_n320_), .B2(new_n322_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n337_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(KEYINPUT89), .A2(G228gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(G233gat), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND4_X1  g145(.A1(new_n317_), .A2(new_n318_), .A3(new_n341_), .A4(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n345_), .A2(KEYINPUT92), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n318_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT29), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n300_), .A2(new_n301_), .A3(new_n302_), .A4(new_n305_), .ZN(new_n351_));
  XNOR2_X1  g150(.A(new_n307_), .B(KEYINPUT88), .ZN(new_n352_));
  OAI21_X1  g151(.A(new_n294_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n316_), .ZN(new_n354_));
  AOI21_X1  g153(.A(new_n350_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  AOI22_X1  g154(.A1(new_n332_), .A2(new_n336_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n356_));
  OAI211_X1 g155(.A(new_n348_), .B(new_n349_), .C1(new_n355_), .C2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n347_), .A2(new_n357_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n358_), .A2(KEYINPUT93), .ZN(new_n359_));
  XNOR2_X1  g158(.A(G78gat), .B(G106gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n359_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT94), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n358_), .A2(KEYINPUT93), .A3(new_n360_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n362_), .A2(new_n363_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n360_), .B1(new_n358_), .B2(KEYINPUT93), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT93), .ZN(new_n367_));
  AOI211_X1 g166(.A(new_n367_), .B(new_n361_), .C1(new_n347_), .C2(new_n357_), .ZN(new_n368_));
  OAI21_X1  g167(.A(KEYINPUT94), .B1(new_n366_), .B2(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT28), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n306_), .A2(new_n309_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n316_), .B1(new_n371_), .B2(new_n294_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n370_), .B1(new_n372_), .B2(new_n350_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n353_), .A2(new_n354_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n375_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  XOR2_X1   g176(.A(G22gat), .B(G50gat), .Z(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n374_), .A2(new_n377_), .A3(new_n379_), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n378_), .B1(new_n373_), .B2(new_n376_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n347_), .A2(new_n357_), .A3(new_n367_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n382_), .A2(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n365_), .A2(new_n369_), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(new_n384_), .B1(new_n365_), .B2(new_n369_), .ZN(new_n386_));
  OAI21_X1  g185(.A(new_n290_), .B1(new_n385_), .B2(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n384_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n363_), .B1(new_n362_), .B2(new_n364_), .ZN(new_n389_));
  NOR3_X1   g188(.A1(new_n366_), .A2(new_n368_), .A3(KEYINPUT94), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n388_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NOR3_X1   g190(.A1(new_n280_), .A2(new_n281_), .A3(new_n202_), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n288_), .B1(new_n286_), .B2(new_n287_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n365_), .A2(new_n369_), .A3(new_n384_), .ZN(new_n395_));
  NAND3_X1  g194(.A1(new_n391_), .A2(new_n394_), .A3(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n387_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT20), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n398_), .B1(new_n267_), .B2(new_n356_), .ZN(new_n399_));
  AOI22_X1  g198(.A1(new_n259_), .A2(new_n261_), .B1(new_n240_), .B2(new_n241_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n226_), .A2(new_n219_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n221_), .A2(new_n225_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n402_), .A2(KEYINPUT24), .A3(new_n219_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n245_), .A2(new_n247_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n248_), .A2(new_n250_), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n403_), .B(new_n254_), .C1(new_n404_), .C2(new_n405_), .ZN(new_n406_));
  AOI21_X1  g205(.A(KEYINPUT83), .B1(new_n260_), .B2(G190gat), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n238_), .A2(new_n237_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  OAI22_X1  g208(.A1(new_n400_), .A2(new_n401_), .B1(new_n406_), .B2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT95), .ZN(new_n411_));
  AND3_X1   g210(.A1(new_n410_), .A2(new_n411_), .A3(new_n341_), .ZN(new_n412_));
  AOI21_X1  g211(.A(new_n411_), .B1(new_n410_), .B2(new_n341_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n399_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G226gat), .A2(G233gat), .ZN(new_n415_));
  XNOR2_X1  g214(.A(new_n415_), .B(KEYINPUT19), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n264_), .A2(new_n341_), .ZN(new_n418_));
  OR2_X1    g217(.A1(new_n410_), .A2(new_n341_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n416_), .A2(new_n398_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n418_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  XOR2_X1   g220(.A(G8gat), .B(G36gat), .Z(new_n422_));
  XNOR2_X1  g221(.A(new_n422_), .B(KEYINPUT18), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G64gat), .B(G92gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n423_), .B(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n417_), .A2(new_n421_), .A3(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n425_), .B1(new_n417_), .B2(new_n421_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n426_), .B1(new_n427_), .B2(KEYINPUT96), .ZN(new_n428_));
  AND2_X1   g227(.A1(new_n418_), .A2(new_n420_), .ZN(new_n429_));
  AOI22_X1  g228(.A1(new_n419_), .A2(new_n429_), .B1(new_n414_), .B2(new_n416_), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT96), .ZN(new_n431_));
  NAND3_X1  g230(.A1(new_n430_), .A2(new_n431_), .A3(new_n425_), .ZN(new_n432_));
  AOI21_X1  g231(.A(KEYINPUT27), .B1(new_n428_), .B2(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(new_n270_), .B(new_n271_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n353_), .A2(new_n434_), .A3(new_n354_), .ZN(new_n435_));
  OAI211_X1 g234(.A(KEYINPUT4), .B(new_n435_), .C1(new_n372_), .C2(new_n276_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n283_), .A2(new_n437_), .A3(new_n375_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G225gat), .A2(G233gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n439_), .B(KEYINPUT97), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n436_), .A2(new_n438_), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT98), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  NAND4_X1  g242(.A1(new_n436_), .A2(new_n438_), .A3(KEYINPUT98), .A4(new_n440_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n283_), .A2(new_n375_), .ZN(new_n446_));
  AND2_X1   g245(.A1(new_n446_), .A2(new_n435_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n439_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n445_), .A2(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(G1gat), .B(G29gat), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n450_), .B(KEYINPUT0), .ZN(new_n451_));
  OR2_X1    g250(.A1(new_n451_), .A2(G57gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(G57gat), .ZN(new_n453_));
  AND3_X1   g252(.A1(new_n452_), .A2(G85gat), .A3(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(G85gat), .B1(new_n452_), .B2(new_n453_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n449_), .A2(new_n456_), .ZN(new_n457_));
  AOI22_X1  g256(.A1(new_n443_), .A2(new_n444_), .B1(new_n447_), .B2(new_n439_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n456_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n458_), .A2(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n457_), .A2(new_n460_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(KEYINPUT100), .B(KEYINPUT20), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n418_), .A2(new_n419_), .A3(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(new_n416_), .ZN(new_n464_));
  INV_X1    g263(.A(new_n416_), .ZN(new_n465_));
  OAI211_X1 g264(.A(new_n399_), .B(new_n465_), .C1(new_n412_), .C2(new_n413_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n464_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n425_), .ZN(new_n468_));
  NAND2_X1  g267(.A1(new_n467_), .A2(new_n468_), .ZN(new_n469_));
  NAND3_X1  g268(.A1(new_n469_), .A2(KEYINPUT27), .A3(new_n426_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  NOR3_X1   g270(.A1(new_n433_), .A2(new_n461_), .A3(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n425_), .A2(KEYINPUT32), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n473_), .B1(new_n464_), .B2(new_n466_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n474_), .B1(new_n430_), .B2(new_n473_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n458_), .A2(new_n459_), .ZN(new_n476_));
  AND3_X1   g275(.A1(new_n445_), .A2(new_n448_), .A3(new_n459_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n476_), .B2(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT33), .ZN(new_n479_));
  AND4_X1   g278(.A1(new_n479_), .A2(new_n445_), .A3(new_n448_), .A4(new_n459_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n479_), .B1(new_n458_), .B2(new_n459_), .ZN(new_n481_));
  NOR2_X1   g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n436_), .A2(new_n439_), .A3(new_n438_), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n446_), .A2(new_n435_), .A3(new_n440_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n456_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n485_), .A2(KEYINPUT99), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT99), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n456_), .A2(new_n483_), .A3(new_n487_), .A4(new_n484_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n428_), .A2(new_n432_), .A3(new_n489_), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n478_), .B1(new_n482_), .B2(new_n490_), .ZN(new_n491_));
  AOI21_X1  g290(.A(new_n290_), .B1(new_n391_), .B2(new_n395_), .ZN(new_n492_));
  AOI22_X1  g291(.A1(new_n397_), .A2(new_n472_), .B1(new_n491_), .B2(new_n492_), .ZN(new_n493_));
  XOR2_X1   g292(.A(G113gat), .B(G141gat), .Z(new_n494_));
  XNOR2_X1  g293(.A(new_n494_), .B(KEYINPUT79), .ZN(new_n495_));
  XOR2_X1   g294(.A(G169gat), .B(G197gat), .Z(new_n496_));
  XNOR2_X1  g295(.A(new_n495_), .B(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(G229gat), .A2(G233gat), .ZN(new_n499_));
  XNOR2_X1  g298(.A(G1gat), .B(G8gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n500_), .B(KEYINPUT76), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G15gat), .B(G22gat), .ZN(new_n502_));
  INV_X1    g301(.A(G1gat), .ZN(new_n503_));
  INV_X1    g302(.A(G8gat), .ZN(new_n504_));
  OAI21_X1  g303(.A(KEYINPUT14), .B1(new_n503_), .B2(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n501_), .A2(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G29gat), .B(G36gat), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n511_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(new_n509_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n512_), .A2(new_n514_), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n500_), .A2(KEYINPUT76), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n500_), .A2(KEYINPUT76), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n516_), .A2(new_n506_), .A3(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n508_), .A2(new_n515_), .A3(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n512_), .A2(new_n514_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT15), .ZN(new_n521_));
  INV_X1    g320(.A(new_n518_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n506_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n522_), .A2(new_n523_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n499_), .B(new_n519_), .C1(new_n521_), .C2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n499_), .ZN(new_n526_));
  NOR3_X1   g325(.A1(new_n522_), .A2(new_n523_), .A3(new_n520_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n515_), .B1(new_n508_), .B2(new_n518_), .ZN(new_n528_));
  OAI211_X1 g327(.A(KEYINPUT78), .B(new_n526_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n525_), .A2(new_n529_), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n520_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n531_), .A2(new_n519_), .ZN(new_n532_));
  AOI21_X1  g331(.A(KEYINPUT78), .B1(new_n532_), .B2(new_n526_), .ZN(new_n533_));
  OAI21_X1  g332(.A(new_n498_), .B1(new_n530_), .B2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT78), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n527_), .A2(new_n528_), .ZN(new_n536_));
  OAI21_X1  g335(.A(new_n535_), .B1(new_n536_), .B2(new_n499_), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n537_), .A2(new_n529_), .A3(new_n525_), .A4(new_n497_), .ZN(new_n538_));
  AND3_X1   g337(.A1(new_n534_), .A2(new_n538_), .A3(KEYINPUT80), .ZN(new_n539_));
  AOI21_X1  g338(.A(KEYINPUT80), .B1(new_n534_), .B2(new_n538_), .ZN(new_n540_));
  NOR2_X1   g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI21_X1  g340(.A(KEYINPUT101), .B1(new_n493_), .B2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT101), .ZN(new_n543_));
  INV_X1    g342(.A(new_n541_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n476_), .A2(new_n477_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n426_), .A2(KEYINPUT96), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n431_), .B1(new_n430_), .B2(new_n425_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n546_), .B1(new_n426_), .B2(new_n547_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n545_), .B(new_n470_), .C1(new_n548_), .C2(KEYINPUT27), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n549_), .B1(new_n396_), .B2(new_n387_), .ZN(new_n550_));
  AND2_X1   g349(.A1(new_n491_), .A2(new_n492_), .ZN(new_n551_));
  OAI211_X1 g350(.A(new_n543_), .B(new_n544_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT71), .ZN(new_n553_));
  OR2_X1    g352(.A1(new_n553_), .A2(KEYINPUT13), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n553_), .A2(KEYINPUT13), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT67), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G57gat), .B(G64gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(G71gat), .B(G78gat), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n557_), .A2(new_n558_), .A3(KEYINPUT11), .ZN(new_n559_));
  INV_X1    g358(.A(G64gat), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n560_), .A2(G57gat), .ZN(new_n561_));
  INV_X1    g360(.A(G57gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(G64gat), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n561_), .A2(new_n563_), .A3(KEYINPUT11), .ZN(new_n564_));
  AND2_X1   g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565_));
  NOR2_X1   g364(.A1(G71gat), .A2(G78gat), .ZN(new_n566_));
  NOR2_X1   g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n564_), .A2(new_n567_), .ZN(new_n568_));
  NOR2_X1   g367(.A1(new_n557_), .A2(KEYINPUT11), .ZN(new_n569_));
  OAI211_X1 g368(.A(new_n556_), .B(new_n559_), .C1(new_n568_), .C2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT11), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n562_), .A2(G64gat), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n560_), .A2(G57gat), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n572_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n575_), .A2(new_n564_), .A3(new_n567_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n556_), .B1(new_n576_), .B2(new_n559_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n571_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT65), .ZN(new_n579_));
  INV_X1    g378(.A(KEYINPUT7), .ZN(new_n580_));
  INV_X1    g379(.A(G99gat), .ZN(new_n581_));
  INV_X1    g380(.A(G106gat), .ZN(new_n582_));
  NAND4_X1  g381(.A1(new_n579_), .A2(new_n580_), .A3(new_n581_), .A4(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(G99gat), .A2(G106gat), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT6), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n587_));
  OAI22_X1  g386(.A1(KEYINPUT65), .A2(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n588_));
  NAND4_X1  g387(.A1(new_n583_), .A2(new_n586_), .A3(new_n587_), .A4(new_n588_), .ZN(new_n589_));
  XOR2_X1   g388(.A(G85gat), .B(G92gat), .Z(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(KEYINPUT66), .A2(KEYINPUT8), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n589_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n595_));
  OR2_X1    g394(.A1(G85gat), .A2(G92gat), .ZN(new_n596_));
  NAND3_X1  g395(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n596_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(G92gat), .ZN(new_n600_));
  OR2_X1    g399(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n601_));
  NAND2_X1  g400(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n602_));
  AOI21_X1  g401(.A(new_n600_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  OAI21_X1  g402(.A(new_n599_), .B1(new_n603_), .B2(KEYINPUT9), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n586_), .A2(new_n587_), .ZN(new_n605_));
  XOR2_X1   g404(.A(KEYINPUT10), .B(G99gat), .Z(new_n606_));
  AOI21_X1  g405(.A(new_n605_), .B1(new_n606_), .B2(new_n582_), .ZN(new_n607_));
  AOI22_X1  g406(.A1(new_n594_), .A2(new_n595_), .B1(new_n604_), .B2(new_n607_), .ZN(new_n608_));
  OAI21_X1  g407(.A(KEYINPUT68), .B1(new_n578_), .B2(new_n608_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n594_), .A2(new_n595_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n604_), .A2(new_n607_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(KEYINPUT68), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n559_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT67), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(new_n570_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n612_), .A2(new_n613_), .A3(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n608_), .A2(new_n615_), .A3(new_n570_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n609_), .A2(new_n617_), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(G230gat), .A2(G233gat), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n619_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT12), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n623_), .B1(new_n578_), .B2(new_n608_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n604_), .A2(new_n607_), .A3(KEYINPUT69), .ZN(new_n625_));
  INV_X1    g424(.A(KEYINPUT69), .ZN(new_n626_));
  AND2_X1   g425(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n627_));
  NOR2_X1   g426(.A1(KEYINPUT64), .A2(G85gat), .ZN(new_n628_));
  OAI21_X1  g427(.A(G92gat), .B1(new_n627_), .B2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT9), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n598_), .B1(new_n629_), .B2(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(KEYINPUT10), .B(G99gat), .ZN(new_n632_));
  OAI211_X1 g431(.A(new_n586_), .B(new_n587_), .C1(new_n632_), .C2(G106gat), .ZN(new_n633_));
  OAI21_X1  g432(.A(new_n626_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n592_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n589_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n625_), .B(new_n634_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n576_), .A2(KEYINPUT12), .A3(new_n559_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n624_), .A2(new_n620_), .A3(new_n618_), .A4(new_n640_), .ZN(new_n641_));
  XNOR2_X1  g440(.A(G120gat), .B(G148gat), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT5), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT70), .ZN(new_n644_));
  XNOR2_X1  g443(.A(G176gat), .B(G204gat), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n644_), .B(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n622_), .A2(new_n641_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n647_), .B1(new_n622_), .B2(new_n641_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n554_), .B(new_n555_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n650_), .ZN(new_n652_));
  NAND4_X1  g451(.A1(new_n652_), .A2(new_n553_), .A3(KEYINPUT13), .A4(new_n648_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n651_), .A2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n542_), .A2(new_n552_), .A3(new_n655_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(G232gat), .A2(G233gat), .ZN(new_n657_));
  XOR2_X1   g456(.A(new_n657_), .B(KEYINPUT34), .Z(new_n658_));
  INV_X1    g457(.A(KEYINPUT35), .ZN(new_n659_));
  NOR2_X1   g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n610_), .A2(new_n515_), .A3(new_n611_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT72), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n658_), .A2(new_n659_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n661_), .A2(new_n662_), .A3(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT15), .ZN(new_n665_));
  XNOR2_X1  g464(.A(new_n520_), .B(new_n665_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n666_), .A2(new_n637_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n664_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n662_), .B1(new_n661_), .B2(new_n663_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n660_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  XNOR2_X1  g469(.A(new_n660_), .B(KEYINPUT74), .ZN(new_n671_));
  NAND4_X1  g470(.A1(new_n667_), .A2(new_n663_), .A3(new_n661_), .A4(new_n671_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(G190gat), .B(G218gat), .ZN(new_n673_));
  XNOR2_X1  g472(.A(G134gat), .B(G162gat), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n673_), .B(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT36), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT73), .ZN(new_n677_));
  OR2_X1    g476(.A1(new_n676_), .A2(KEYINPUT73), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n675_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n670_), .A2(new_n672_), .A3(new_n679_), .ZN(new_n680_));
  INV_X1    g479(.A(new_n672_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n661_), .A2(new_n663_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n682_), .A2(KEYINPUT72), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(new_n664_), .A3(new_n667_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n681_), .B1(new_n684_), .B2(new_n660_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n675_), .B(KEYINPUT36), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n680_), .B(KEYINPUT75), .C1(new_n685_), .C2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT37), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  AND2_X1   g488(.A1(G231gat), .A2(G233gat), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n524_), .B(new_n690_), .ZN(new_n691_));
  XOR2_X1   g490(.A(new_n691_), .B(new_n614_), .Z(new_n692_));
  XNOR2_X1  g491(.A(G127gat), .B(G155gat), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT16), .ZN(new_n694_));
  XNOR2_X1  g493(.A(G183gat), .B(G211gat), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n694_), .B(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT17), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(KEYINPUT77), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT67), .B1(new_n696_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n692_), .A2(new_n699_), .ZN(new_n700_));
  XNOR2_X1  g499(.A(new_n691_), .B(new_n614_), .ZN(new_n701_));
  INV_X1    g500(.A(new_n696_), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n556_), .B1(new_n702_), .B2(new_n697_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n696_), .A2(KEYINPUT17), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n697_), .A2(KEYINPUT77), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n705_), .B1(new_n696_), .B2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n700_), .A2(new_n704_), .A3(new_n707_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n670_), .A2(new_n672_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n686_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n711_), .A2(KEYINPUT75), .A3(KEYINPUT37), .A4(new_n680_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n689_), .A2(new_n708_), .A3(new_n712_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n656_), .A2(new_n713_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(new_n503_), .A3(new_n461_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(KEYINPUT38), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(KEYINPUT38), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n544_), .A2(new_n653_), .A3(new_n651_), .ZN(new_n718_));
  OR2_X1    g517(.A1(new_n718_), .A2(KEYINPUT102), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n718_), .A2(KEYINPUT102), .ZN(new_n720_));
  AND3_X1   g519(.A1(new_n719_), .A2(new_n720_), .A3(new_n708_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n711_), .A2(new_n680_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n722_), .ZN(new_n723_));
  NOR2_X1   g522(.A1(new_n493_), .A2(new_n723_), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n721_), .A2(new_n461_), .A3(new_n724_), .ZN(new_n725_));
  OAI22_X1  g524(.A1(new_n716_), .A2(new_n717_), .B1(new_n503_), .B2(new_n725_), .ZN(G1324gat));
  INV_X1    g525(.A(new_n433_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n727_), .A2(new_n470_), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n714_), .A2(new_n504_), .A3(new_n728_), .ZN(new_n729_));
  NAND3_X1  g528(.A1(new_n721_), .A2(new_n728_), .A3(new_n724_), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT39), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n730_), .A2(new_n731_), .A3(G8gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n731_), .B1(new_n730_), .B2(G8gat), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n729_), .B1(new_n732_), .B2(new_n733_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT40), .Z(G1325gat));
  NAND3_X1  g534(.A1(new_n714_), .A2(new_n206_), .A3(new_n290_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n721_), .A2(new_n290_), .A3(new_n724_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n738_));
  AND3_X1   g537(.A1(new_n737_), .A2(G15gat), .A3(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n738_), .B1(new_n737_), .B2(G15gat), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(G1326gat));
  INV_X1    g540(.A(G22gat), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n385_), .A2(new_n386_), .ZN(new_n743_));
  NAND3_X1  g542(.A1(new_n714_), .A2(new_n742_), .A3(new_n743_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n721_), .A2(new_n743_), .A3(new_n724_), .ZN(new_n745_));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(new_n746_), .A3(G22gat), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(G22gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n744_), .B1(new_n747_), .B2(new_n748_), .ZN(G1327gat));
  NOR2_X1   g548(.A1(new_n708_), .A2(new_n722_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n542_), .A2(new_n552_), .A3(new_n655_), .A4(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  AOI21_X1  g551(.A(G29gat), .B1(new_n752_), .B2(new_n461_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n689_), .A2(new_n712_), .ZN(new_n754_));
  INV_X1    g553(.A(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(KEYINPUT43), .B1(new_n493_), .B2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT43), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(new_n754_), .C1(new_n550_), .C2(new_n551_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n708_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n719_), .A2(new_n720_), .A3(new_n760_), .ZN(new_n761_));
  INV_X1    g560(.A(new_n761_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n759_), .A2(KEYINPUT44), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT105), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n761_), .B1(new_n756_), .B2(new_n758_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n766_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n765_), .A2(new_n767_), .ZN(new_n768_));
  AND3_X1   g567(.A1(new_n768_), .A2(G29gat), .A3(new_n461_), .ZN(new_n769_));
  NOR3_X1   g568(.A1(new_n385_), .A2(new_n386_), .A3(new_n290_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n394_), .B1(new_n391_), .B2(new_n395_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n472_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n491_), .A2(new_n492_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n757_), .B1(new_n774_), .B2(new_n754_), .ZN(new_n775_));
  AOI211_X1 g574(.A(KEYINPUT43), .B(new_n755_), .C1(new_n772_), .C2(new_n773_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n762_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT104), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n777_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(KEYINPUT104), .B1(new_n766_), .B2(KEYINPUT44), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(new_n753_), .B1(new_n769_), .B2(new_n782_), .ZN(G1328gat));
  NAND2_X1  g582(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n784_));
  INV_X1    g583(.A(new_n784_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(KEYINPUT106), .A2(KEYINPUT46), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n788_));
  INV_X1    g587(.A(new_n728_), .ZN(new_n789_));
  NOR2_X1   g588(.A1(new_n789_), .A2(G36gat), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n788_), .B1(new_n752_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n790_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n751_), .A2(KEYINPUT45), .A3(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n787_), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n768_), .A2(new_n782_), .A3(new_n728_), .ZN(new_n795_));
  AOI211_X1 g594(.A(new_n785_), .B(new_n794_), .C1(G36gat), .C2(new_n795_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(G36gat), .ZN(new_n797_));
  INV_X1    g596(.A(new_n794_), .ZN(new_n798_));
  AOI21_X1  g597(.A(new_n784_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n796_), .A2(new_n799_), .ZN(G1329gat));
  NAND4_X1  g599(.A1(new_n768_), .A2(new_n782_), .A3(G43gat), .A4(new_n290_), .ZN(new_n801_));
  OAI21_X1  g600(.A(new_n214_), .B1(new_n751_), .B2(new_n394_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n801_), .A2(new_n802_), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n803_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g603(.A1(new_n768_), .A2(new_n782_), .A3(new_n743_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT107), .ZN(new_n806_));
  AND3_X1   g605(.A1(new_n805_), .A2(new_n806_), .A3(G50gat), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n805_), .B2(G50gat), .ZN(new_n808_));
  INV_X1    g607(.A(new_n743_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n809_), .A2(G50gat), .ZN(new_n810_));
  XNOR2_X1  g609(.A(new_n810_), .B(KEYINPUT108), .ZN(new_n811_));
  OAI22_X1  g610(.A1(new_n807_), .A2(new_n808_), .B1(new_n751_), .B2(new_n811_), .ZN(G1331gat));
  NOR3_X1   g611(.A1(new_n655_), .A2(new_n544_), .A3(new_n760_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n724_), .A2(new_n813_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n814_), .A2(new_n562_), .A3(new_n545_), .ZN(new_n815_));
  NOR2_X1   g614(.A1(new_n655_), .A2(new_n544_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n774_), .A2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n817_), .A2(new_n713_), .ZN(new_n818_));
  INV_X1    g617(.A(new_n818_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n545_), .B1(new_n819_), .B2(KEYINPUT109), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n820_), .B1(KEYINPUT109), .B2(new_n819_), .ZN(new_n821_));
  AOI21_X1  g620(.A(new_n815_), .B1(new_n821_), .B2(new_n562_), .ZN(G1332gat));
  OAI21_X1  g621(.A(G64gat), .B1(new_n814_), .B2(new_n789_), .ZN(new_n823_));
  XOR2_X1   g622(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n824_));
  OR2_X1    g623(.A1(new_n823_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n823_), .A2(new_n824_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n818_), .A2(new_n560_), .A3(new_n728_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n825_), .A2(new_n826_), .A3(new_n827_), .ZN(G1333gat));
  OAI21_X1  g627(.A(G71gat), .B1(new_n814_), .B2(new_n394_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n829_), .A2(KEYINPUT49), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n829_), .A2(KEYINPUT49), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n394_), .A2(G71gat), .ZN(new_n832_));
  XOR2_X1   g631(.A(new_n832_), .B(KEYINPUT111), .Z(new_n833_));
  OAI22_X1  g632(.A1(new_n830_), .A2(new_n831_), .B1(new_n819_), .B2(new_n833_), .ZN(G1334gat));
  OAI21_X1  g633(.A(G78gat), .B1(new_n814_), .B2(new_n809_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n835_), .A2(KEYINPUT50), .ZN(new_n836_));
  NOR2_X1   g635(.A1(new_n835_), .A2(KEYINPUT50), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n809_), .A2(G78gat), .ZN(new_n838_));
  OAI22_X1  g637(.A1(new_n836_), .A2(new_n837_), .B1(new_n819_), .B2(new_n838_), .ZN(G1335gat));
  NOR3_X1   g638(.A1(new_n817_), .A2(new_n722_), .A3(new_n708_), .ZN(new_n840_));
  AOI21_X1  g639(.A(G85gat), .B1(new_n840_), .B2(new_n461_), .ZN(new_n841_));
  AND3_X1   g640(.A1(new_n759_), .A2(new_n760_), .A3(new_n816_), .ZN(new_n842_));
  XNOR2_X1  g641(.A(new_n842_), .B(KEYINPUT112), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n545_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n841_), .B1(new_n843_), .B2(new_n844_), .ZN(G1336gat));
  NAND3_X1  g644(.A1(new_n840_), .A2(new_n600_), .A3(new_n728_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n843_), .A2(new_n728_), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n600_), .ZN(G1337gat));
  AOI21_X1  g647(.A(new_n581_), .B1(new_n842_), .B2(new_n290_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n394_), .A2(new_n632_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n849_), .B1(new_n840_), .B2(new_n850_), .ZN(new_n851_));
  XOR2_X1   g650(.A(new_n851_), .B(KEYINPUT51), .Z(G1338gat));
  NAND3_X1  g651(.A1(new_n840_), .A2(new_n582_), .A3(new_n743_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n842_), .A2(new_n743_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n854_), .B1(new_n855_), .B2(G106gat), .ZN(new_n856_));
  AOI211_X1 g655(.A(KEYINPUT52), .B(new_n582_), .C1(new_n842_), .C2(new_n743_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n853_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT53), .ZN(G1339gat));
  OAI21_X1  g658(.A(new_n648_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n860_));
  AOI22_X1  g659(.A1(new_n610_), .A2(new_n611_), .B1(new_n615_), .B2(new_n570_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n640_), .B(new_n618_), .C1(new_n861_), .C2(KEYINPUT12), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n862_), .A2(new_n621_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n863_), .A2(KEYINPUT116), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT115), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT55), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n641_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n862_), .A2(new_n868_), .A3(new_n621_), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n864_), .A2(new_n867_), .A3(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n866_), .B1(new_n641_), .B2(new_n865_), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n646_), .B1(new_n870_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT56), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n641_), .A2(new_n865_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n875_), .A2(KEYINPUT55), .ZN(new_n876_));
  NAND4_X1  g675(.A1(new_n876_), .A2(new_n867_), .A3(new_n864_), .A4(new_n869_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n877_), .A2(KEYINPUT56), .A3(new_n646_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n860_), .B1(new_n874_), .B2(new_n878_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n526_), .B(new_n519_), .C1(new_n521_), .C2(new_n524_), .ZN(new_n880_));
  OAI211_X1 g679(.A(new_n880_), .B(new_n498_), .C1(new_n536_), .C2(new_n526_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n538_), .A2(new_n881_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n882_), .B1(new_n652_), .B2(new_n648_), .ZN(new_n883_));
  OAI211_X1 g682(.A(KEYINPUT57), .B(new_n722_), .C1(new_n879_), .C2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(KEYINPUT117), .ZN(new_n885_));
  INV_X1    g684(.A(new_n883_), .ZN(new_n886_));
  AND3_X1   g685(.A1(new_n877_), .A2(KEYINPUT56), .A3(new_n646_), .ZN(new_n887_));
  AOI21_X1  g686(.A(KEYINPUT56), .B1(new_n877_), .B2(new_n646_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n887_), .A2(new_n888_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n886_), .B1(new_n889_), .B2(new_n860_), .ZN(new_n890_));
  INV_X1    g689(.A(KEYINPUT117), .ZN(new_n891_));
  NAND4_X1  g690(.A1(new_n890_), .A2(new_n891_), .A3(KEYINPUT57), .A4(new_n722_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n885_), .A2(new_n892_), .ZN(new_n893_));
  NAND3_X1  g692(.A1(new_n648_), .A2(new_n538_), .A3(new_n881_), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n894_), .B1(new_n874_), .B2(new_n878_), .ZN(new_n895_));
  OR2_X1    g694(.A1(new_n895_), .A2(KEYINPUT58), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n755_), .B1(new_n895_), .B2(KEYINPUT58), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n722_), .B1(new_n879_), .B2(new_n883_), .ZN(new_n898_));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n899_));
  AOI22_X1  g698(.A1(new_n896_), .A2(new_n897_), .B1(new_n898_), .B2(new_n899_), .ZN(new_n900_));
  AOI21_X1  g699(.A(new_n708_), .B1(new_n893_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT54), .ZN(new_n902_));
  NAND2_X1  g701(.A1(new_n902_), .A2(KEYINPUT113), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n541_), .A2(new_n651_), .A3(new_n653_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n713_), .B2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(KEYINPUT114), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT114), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n907_), .B(new_n903_), .C1(new_n713_), .C2(new_n904_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n906_), .A2(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n902_), .A2(KEYINPUT113), .ZN(new_n910_));
  INV_X1    g709(.A(new_n910_), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n906_), .A2(new_n910_), .A3(new_n908_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n912_), .A2(new_n913_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n901_), .A2(new_n914_), .ZN(new_n915_));
  NOR2_X1   g714(.A1(new_n387_), .A2(new_n545_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n915_), .A2(new_n789_), .A3(new_n916_), .ZN(new_n917_));
  INV_X1    g716(.A(new_n917_), .ZN(new_n918_));
  INV_X1    g717(.A(G113gat), .ZN(new_n919_));
  NAND3_X1  g718(.A1(new_n918_), .A2(new_n919_), .A3(new_n544_), .ZN(new_n920_));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n917_), .A2(new_n921_), .ZN(new_n922_));
  NAND4_X1  g721(.A1(new_n915_), .A2(KEYINPUT59), .A3(new_n789_), .A4(new_n916_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n541_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n920_), .B1(new_n924_), .B2(new_n919_), .ZN(G1340gat));
  INV_X1    g724(.A(KEYINPUT60), .ZN(new_n926_));
  INV_X1    g725(.A(G120gat), .ZN(new_n927_));
  NAND3_X1  g726(.A1(new_n654_), .A2(new_n926_), .A3(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n928_), .B1(new_n926_), .B2(new_n927_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n918_), .A2(new_n929_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n655_), .B1(new_n922_), .B2(new_n923_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n931_), .B2(new_n927_), .ZN(G1341gat));
  AOI21_X1  g731(.A(G127gat), .B1(new_n918_), .B2(new_n708_), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n922_), .A2(new_n923_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n708_), .A2(G127gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT118), .ZN(new_n936_));
  AOI21_X1  g735(.A(new_n933_), .B1(new_n934_), .B2(new_n936_), .ZN(G1342gat));
  AOI21_X1  g736(.A(G134gat), .B1(new_n918_), .B2(new_n723_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n754_), .A2(G134gat), .ZN(new_n939_));
  XOR2_X1   g738(.A(new_n939_), .B(KEYINPUT119), .Z(new_n940_));
  AOI21_X1  g739(.A(new_n938_), .B1(new_n934_), .B2(new_n940_), .ZN(G1343gat));
  NOR2_X1   g740(.A1(new_n396_), .A2(new_n545_), .ZN(new_n942_));
  OAI211_X1 g741(.A(new_n942_), .B(new_n789_), .C1(new_n901_), .C2(new_n914_), .ZN(new_n943_));
  INV_X1    g742(.A(KEYINPUT120), .ZN(new_n944_));
  XNOR2_X1  g743(.A(new_n943_), .B(new_n944_), .ZN(new_n945_));
  OAI21_X1  g744(.A(G141gat), .B1(new_n945_), .B2(new_n541_), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n915_), .A2(new_n944_), .A3(new_n789_), .A4(new_n942_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n943_), .A2(KEYINPUT120), .ZN(new_n948_));
  NAND2_X1  g747(.A1(new_n947_), .A2(new_n948_), .ZN(new_n949_));
  NAND3_X1  g748(.A1(new_n949_), .A2(new_n298_), .A3(new_n544_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n946_), .A2(new_n950_), .ZN(G1344gat));
  OAI21_X1  g750(.A(G148gat), .B1(new_n945_), .B2(new_n655_), .ZN(new_n952_));
  NAND3_X1  g751(.A1(new_n949_), .A2(new_n299_), .A3(new_n654_), .ZN(new_n953_));
  NAND2_X1  g752(.A1(new_n952_), .A2(new_n953_), .ZN(G1345gat));
  XNOR2_X1  g753(.A(KEYINPUT61), .B(G155gat), .ZN(new_n955_));
  AOI21_X1  g754(.A(new_n955_), .B1(new_n949_), .B2(new_n708_), .ZN(new_n956_));
  INV_X1    g755(.A(new_n955_), .ZN(new_n957_));
  AOI211_X1 g756(.A(new_n760_), .B(new_n957_), .C1(new_n947_), .C2(new_n948_), .ZN(new_n958_));
  NOR2_X1   g757(.A1(new_n956_), .A2(new_n958_), .ZN(G1346gat));
  OAI21_X1  g758(.A(G162gat), .B1(new_n945_), .B2(new_n755_), .ZN(new_n960_));
  INV_X1    g759(.A(G162gat), .ZN(new_n961_));
  NAND3_X1  g760(.A1(new_n949_), .A2(new_n961_), .A3(new_n723_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n960_), .A2(new_n962_), .ZN(G1347gat));
  NAND3_X1  g762(.A1(new_n728_), .A2(new_n545_), .A3(new_n290_), .ZN(new_n964_));
  INV_X1    g763(.A(KEYINPUT121), .ZN(new_n965_));
  OR2_X1    g764(.A1(new_n964_), .A2(new_n965_), .ZN(new_n966_));
  NAND2_X1  g765(.A1(new_n964_), .A2(new_n965_), .ZN(new_n967_));
  AOI21_X1  g766(.A(new_n743_), .B1(new_n966_), .B2(new_n967_), .ZN(new_n968_));
  OAI211_X1 g767(.A(new_n544_), .B(new_n968_), .C1(new_n901_), .C2(new_n914_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n969_), .A2(G169gat), .ZN(new_n970_));
  XOR2_X1   g769(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n971_));
  NAND2_X1  g770(.A1(new_n970_), .A2(new_n971_), .ZN(new_n972_));
  INV_X1    g771(.A(new_n971_), .ZN(new_n973_));
  NAND3_X1  g772(.A1(new_n969_), .A2(G169gat), .A3(new_n973_), .ZN(new_n974_));
  NAND2_X1  g773(.A1(new_n972_), .A2(new_n974_), .ZN(new_n975_));
  NAND2_X1  g774(.A1(new_n544_), .A2(new_n228_), .ZN(new_n976_));
  OAI21_X1  g775(.A(new_n968_), .B1(new_n901_), .B2(new_n914_), .ZN(new_n977_));
  NAND2_X1  g776(.A1(new_n977_), .A2(KEYINPUT123), .ZN(new_n978_));
  INV_X1    g777(.A(KEYINPUT123), .ZN(new_n979_));
  OAI211_X1 g778(.A(new_n979_), .B(new_n968_), .C1(new_n901_), .C2(new_n914_), .ZN(new_n980_));
  AOI21_X1  g779(.A(new_n976_), .B1(new_n978_), .B2(new_n980_), .ZN(new_n981_));
  OAI21_X1  g780(.A(KEYINPUT124), .B1(new_n975_), .B2(new_n981_), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n978_), .A2(new_n980_), .ZN(new_n983_));
  INV_X1    g782(.A(new_n976_), .ZN(new_n984_));
  NAND2_X1  g783(.A1(new_n983_), .A2(new_n984_), .ZN(new_n985_));
  INV_X1    g784(.A(KEYINPUT124), .ZN(new_n986_));
  NAND4_X1  g785(.A1(new_n985_), .A2(new_n986_), .A3(new_n974_), .A4(new_n972_), .ZN(new_n987_));
  NAND2_X1  g786(.A1(new_n982_), .A2(new_n987_), .ZN(G1348gat));
  AOI21_X1  g787(.A(G176gat), .B1(new_n983_), .B2(new_n654_), .ZN(new_n989_));
  INV_X1    g788(.A(new_n977_), .ZN(new_n990_));
  NOR2_X1   g789(.A1(new_n655_), .A2(new_n225_), .ZN(new_n991_));
  AOI21_X1  g790(.A(KEYINPUT125), .B1(new_n990_), .B2(new_n991_), .ZN(new_n992_));
  AND3_X1   g791(.A1(new_n990_), .A2(KEYINPUT125), .A3(new_n991_), .ZN(new_n993_));
  NOR3_X1   g792(.A1(new_n989_), .A2(new_n992_), .A3(new_n993_), .ZN(G1349gat));
  AOI21_X1  g793(.A(G183gat), .B1(new_n990_), .B2(new_n708_), .ZN(new_n995_));
  AND2_X1   g794(.A1(new_n708_), .A2(new_n404_), .ZN(new_n996_));
  AOI21_X1  g795(.A(new_n995_), .B1(new_n983_), .B2(new_n996_), .ZN(G1350gat));
  INV_X1    g796(.A(new_n983_), .ZN(new_n998_));
  OR2_X1    g797(.A1(new_n722_), .A2(new_n405_), .ZN(new_n999_));
  AOI21_X1  g798(.A(new_n755_), .B1(new_n978_), .B2(new_n980_), .ZN(new_n1000_));
  OAI22_X1  g799(.A1(new_n998_), .A2(new_n999_), .B1(new_n1000_), .B2(new_n241_), .ZN(G1351gat));
  NOR2_X1   g800(.A1(new_n901_), .A2(new_n914_), .ZN(new_n1002_));
  NAND2_X1  g801(.A1(new_n728_), .A2(new_n545_), .ZN(new_n1003_));
  NOR2_X1   g802(.A1(new_n1003_), .A2(new_n396_), .ZN(new_n1004_));
  INV_X1    g803(.A(new_n1004_), .ZN(new_n1005_));
  NOR2_X1   g804(.A1(new_n1002_), .A2(new_n1005_), .ZN(new_n1006_));
  NAND2_X1  g805(.A1(new_n1006_), .A2(new_n544_), .ZN(new_n1007_));
  XNOR2_X1  g806(.A(new_n1007_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g807(.A1(new_n1006_), .A2(new_n654_), .ZN(new_n1009_));
  XNOR2_X1  g808(.A(new_n1009_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g809(.A1(new_n1006_), .A2(new_n708_), .ZN(new_n1011_));
  OAI21_X1  g810(.A(new_n1011_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n1012_));
  XOR2_X1   g811(.A(KEYINPUT63), .B(G211gat), .Z(new_n1013_));
  OAI21_X1  g812(.A(new_n1012_), .B1(new_n1011_), .B2(new_n1013_), .ZN(G1354gat));
  NAND3_X1  g813(.A1(new_n915_), .A2(new_n723_), .A3(new_n1004_), .ZN(new_n1015_));
  XOR2_X1   g814(.A(KEYINPUT126), .B(G218gat), .Z(new_n1016_));
  NAND2_X1  g815(.A1(new_n1015_), .A2(new_n1016_), .ZN(new_n1017_));
  NOR2_X1   g816(.A1(new_n755_), .A2(new_n1016_), .ZN(new_n1018_));
  NAND2_X1  g817(.A1(new_n1006_), .A2(new_n1018_), .ZN(new_n1019_));
  NAND2_X1  g818(.A1(new_n1017_), .A2(new_n1019_), .ZN(new_n1020_));
  INV_X1    g819(.A(KEYINPUT127), .ZN(new_n1021_));
  NAND2_X1  g820(.A1(new_n1020_), .A2(new_n1021_), .ZN(new_n1022_));
  NAND3_X1  g821(.A1(new_n1017_), .A2(KEYINPUT127), .A3(new_n1019_), .ZN(new_n1023_));
  NAND2_X1  g822(.A1(new_n1022_), .A2(new_n1023_), .ZN(G1355gat));
endmodule


