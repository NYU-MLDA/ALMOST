//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n759_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n793_, new_n794_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n800_, new_n801_, new_n802_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n879_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n886_, new_n887_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n902_,
    new_n903_, new_n904_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_, new_n920_, new_n921_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n930_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n940_, new_n941_, new_n942_, new_n943_,
    new_n944_, new_n945_, new_n947_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n955_, new_n956_, new_n957_;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT7), .ZN(new_n203_));
  INV_X1    g002(.A(G99gat), .ZN(new_n204_));
  INV_X1    g003(.A(G106gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n203_), .A2(new_n204_), .A3(new_n205_), .ZN(new_n206_));
  OAI21_X1  g005(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G99gat), .A2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(G99gat), .A3(G106gat), .ZN(new_n212_));
  AND3_X1   g011(.A1(new_n210_), .A2(new_n212_), .A3(KEYINPUT66), .ZN(new_n213_));
  AOI21_X1  g012(.A(KEYINPUT66), .B1(new_n210_), .B2(new_n212_), .ZN(new_n214_));
  OAI21_X1  g013(.A(new_n208_), .B1(new_n213_), .B2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT8), .ZN(new_n216_));
  INV_X1    g015(.A(KEYINPUT67), .ZN(new_n217_));
  AND2_X1   g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(G85gat), .A2(G92gat), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n217_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(G85gat), .ZN(new_n221_));
  INV_X1    g020(.A(G92gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G85gat), .A2(G92gat), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(KEYINPUT67), .A3(new_n224_), .ZN(new_n225_));
  AND2_X1   g024(.A1(new_n220_), .A2(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n215_), .A2(new_n216_), .A3(new_n226_), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n210_), .A2(new_n212_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n228_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n220_), .A2(new_n225_), .ZN(new_n230_));
  OAI21_X1  g029(.A(KEYINPUT8), .B1(new_n229_), .B2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(new_n231_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n221_), .A2(KEYINPUT65), .ZN(new_n233_));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(G85gat), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  NOR2_X1   g035(.A1(new_n222_), .A2(KEYINPUT9), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n223_), .A2(KEYINPUT9), .A3(new_n224_), .ZN(new_n239_));
  OAI211_X1 g038(.A(new_n238_), .B(new_n239_), .C1(new_n213_), .C2(new_n214_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n240_), .ZN(new_n241_));
  INV_X1    g040(.A(KEYINPUT10), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(new_n204_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n244_));
  NAND3_X1  g043(.A1(new_n243_), .A2(KEYINPUT64), .A3(new_n244_), .ZN(new_n245_));
  INV_X1    g044(.A(new_n245_), .ZN(new_n246_));
  AOI21_X1  g045(.A(KEYINPUT64), .B1(new_n243_), .B2(new_n244_), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n205_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n241_), .A2(new_n248_), .ZN(new_n249_));
  XNOR2_X1  g048(.A(G57gat), .B(G64gat), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n252_));
  XOR2_X1   g051(.A(G71gat), .B(G78gat), .Z(new_n253_));
  NAND3_X1  g052(.A1(new_n251_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  OR2_X1    g053(.A1(new_n252_), .A2(new_n253_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n254_), .A2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n232_), .A2(new_n249_), .A3(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT12), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n232_), .A2(new_n249_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n256_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n258_), .B1(new_n259_), .B2(new_n262_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(G230gat), .A2(G233gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n243_), .A2(new_n244_), .ZN(new_n265_));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  AOI21_X1  g066(.A(G106gat), .B1(new_n267_), .B2(new_n245_), .ZN(new_n268_));
  OAI21_X1  g067(.A(KEYINPUT69), .B1(new_n240_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n211_), .B1(G99gat), .B2(G106gat), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n209_), .A2(KEYINPUT6), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n270_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n210_), .A2(new_n212_), .A3(KEYINPUT66), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT69), .ZN(new_n276_));
  NOR2_X1   g075(.A1(new_n218_), .A2(new_n219_), .ZN(new_n277_));
  AOI22_X1  g076(.A1(new_n236_), .A2(new_n237_), .B1(new_n277_), .B2(KEYINPUT9), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n248_), .A2(new_n275_), .A3(new_n276_), .A4(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n269_), .A2(new_n279_), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n220_), .A2(new_n225_), .A3(new_n216_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(new_n275_), .B2(new_n208_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n228_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n216_), .B1(new_n226_), .B2(new_n283_), .ZN(new_n284_));
  OAI21_X1  g083(.A(KEYINPUT68), .B1(new_n282_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n227_), .A2(new_n286_), .A3(new_n231_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n280_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n288_), .A2(KEYINPUT12), .A3(new_n261_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n263_), .A2(new_n264_), .A3(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n262_), .A2(new_n257_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n291_), .A2(G230gat), .A3(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G120gat), .B(G148gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n293_), .B(KEYINPUT5), .ZN(new_n294_));
  XNOR2_X1  g093(.A(G176gat), .B(G204gat), .ZN(new_n295_));
  XOR2_X1   g094(.A(new_n294_), .B(new_n295_), .Z(new_n296_));
  INV_X1    g095(.A(new_n296_), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n290_), .A2(new_n292_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n297_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n202_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n300_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n302_), .A2(KEYINPUT70), .A3(new_n298_), .ZN(new_n303_));
  AND3_X1   g102(.A1(new_n301_), .A2(new_n303_), .A3(KEYINPUT13), .ZN(new_n304_));
  AOI21_X1  g103(.A(KEYINPUT13), .B1(new_n301_), .B2(new_n303_), .ZN(new_n305_));
  NOR2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(new_n306_), .B(KEYINPUT71), .Z(new_n307_));
  XOR2_X1   g106(.A(G1gat), .B(G29gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G57gat), .B(G85gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  NAND2_X1  g111(.A1(G225gat), .A2(G233gat), .ZN(new_n313_));
  INV_X1    g112(.A(KEYINPUT3), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n314_), .A2(KEYINPUT85), .ZN(new_n315_));
  INV_X1    g114(.A(G141gat), .ZN(new_n316_));
  INV_X1    g115(.A(G148gat), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT85), .ZN(new_n318_));
  OAI211_X1 g117(.A(new_n316_), .B(new_n317_), .C1(new_n318_), .C2(KEYINPUT3), .ZN(new_n319_));
  OAI211_X1 g118(.A(new_n314_), .B(KEYINPUT85), .C1(G141gat), .C2(G148gat), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n315_), .B1(new_n319_), .B2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT87), .ZN(new_n322_));
  NAND2_X1  g121(.A1(G141gat), .A2(G148gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(new_n323_), .B1(KEYINPUT86), .B2(KEYINPUT2), .ZN(new_n324_));
  NAND2_X1  g123(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n322_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT88), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  NAND4_X1  g129(.A1(KEYINPUT88), .A2(KEYINPUT2), .A3(G141gat), .A4(G148gat), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  OR2_X1    g131(.A1(KEYINPUT86), .A2(KEYINPUT2), .ZN(new_n333_));
  NAND4_X1  g132(.A1(new_n333_), .A2(KEYINPUT87), .A3(new_n325_), .A4(new_n323_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n321_), .A2(new_n327_), .A3(new_n332_), .A4(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(G155gat), .A2(G162gat), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(G155gat), .A2(G162gat), .ZN(new_n338_));
  NOR2_X1   g137(.A1(new_n337_), .A2(new_n338_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n339_), .ZN(new_n340_));
  NOR3_X1   g139(.A1(new_n337_), .A2(new_n338_), .A3(KEYINPUT1), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n316_), .A2(new_n317_), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT1), .ZN(new_n343_));
  OAI211_X1 g142(.A(new_n342_), .B(new_n323_), .C1(new_n343_), .C2(new_n336_), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n341_), .A2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n340_), .A2(new_n346_), .ZN(new_n347_));
  XOR2_X1   g146(.A(G127gat), .B(G134gat), .Z(new_n348_));
  XOR2_X1   g147(.A(G113gat), .B(G120gat), .Z(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  OAI21_X1  g149(.A(KEYINPUT96), .B1(new_n347_), .B2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT89), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n352_), .B1(new_n340_), .B2(new_n346_), .ZN(new_n353_));
  AOI211_X1 g152(.A(KEYINPUT89), .B(new_n345_), .C1(new_n335_), .C2(new_n339_), .ZN(new_n354_));
  NOR2_X1   g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n351_), .B1(new_n355_), .B2(new_n350_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n350_), .ZN(new_n357_));
  NOR4_X1   g156(.A1(new_n353_), .A2(new_n354_), .A3(KEYINPUT96), .A4(new_n357_), .ZN(new_n358_));
  OAI21_X1  g157(.A(new_n313_), .B1(new_n356_), .B2(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n359_), .A2(KEYINPUT98), .ZN(new_n360_));
  INV_X1    g159(.A(new_n339_), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n327_), .A2(new_n334_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n319_), .A2(new_n320_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n315_), .ZN(new_n364_));
  AND3_X1   g163(.A1(new_n363_), .A2(new_n332_), .A3(new_n364_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n361_), .B1(new_n362_), .B2(new_n365_), .ZN(new_n366_));
  OAI21_X1  g165(.A(KEYINPUT89), .B1(new_n366_), .B2(new_n345_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT96), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n345_), .B1(new_n335_), .B2(new_n339_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n369_), .A2(new_n352_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n367_), .A2(new_n368_), .A3(new_n350_), .A4(new_n370_), .ZN(new_n371_));
  NOR3_X1   g170(.A1(new_n353_), .A2(new_n354_), .A3(new_n357_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n371_), .B1(new_n372_), .B2(new_n351_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT98), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n313_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n360_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n373_), .A2(KEYINPUT4), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT4), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n313_), .B1(new_n372_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n377_), .A2(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n312_), .B1(new_n376_), .B2(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n313_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n367_), .A2(new_n350_), .A3(new_n370_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n368_), .B1(new_n357_), .B2(new_n369_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  AOI211_X1 g184(.A(KEYINPUT98), .B(new_n382_), .C1(new_n385_), .C2(new_n371_), .ZN(new_n386_));
  AOI21_X1  g185(.A(new_n374_), .B1(new_n373_), .B2(new_n313_), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n378_), .B1(new_n385_), .B2(new_n371_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n379_), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n312_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NOR2_X1   g190(.A1(new_n388_), .A2(new_n391_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n381_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(G169gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(KEYINPUT84), .B(G190gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n396_), .A2(G183gat), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G183gat), .A2(G190gat), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT23), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n395_), .B1(new_n397_), .B2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(KEYINPUT25), .B(G183gat), .ZN(new_n404_));
  INV_X1    g203(.A(new_n404_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n396_), .A2(KEYINPUT26), .ZN(new_n406_));
  OR2_X1    g205(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n407_));
  AOI21_X1  g206(.A(new_n405_), .B1(new_n406_), .B2(new_n407_), .ZN(new_n408_));
  INV_X1    g207(.A(new_n402_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(G169gat), .ZN(new_n412_));
  INV_X1    g211(.A(G176gat), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n411_), .B1(new_n412_), .B2(new_n413_), .ZN(new_n414_));
  OR3_X1    g213(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n409_), .A2(new_n414_), .A3(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n403_), .B1(new_n408_), .B2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(G71gat), .B(G99gat), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n418_), .B(G43gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n417_), .B(new_n419_), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(new_n357_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(G227gat), .A2(G233gat), .ZN(new_n422_));
  INV_X1    g221(.A(G15gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT30), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n425_), .B(KEYINPUT31), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n421_), .B(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n393_), .A2(new_n427_), .ZN(new_n428_));
  AND2_X1   g227(.A1(G228gat), .A2(G233gat), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT91), .ZN(new_n430_));
  INV_X1    g229(.A(KEYINPUT29), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n430_), .B1(new_n369_), .B2(new_n431_), .ZN(new_n432_));
  XNOR2_X1  g231(.A(G211gat), .B(G218gat), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n433_), .A2(KEYINPUT21), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G197gat), .B(G204gat), .ZN(new_n435_));
  NOR2_X1   g234(.A1(new_n434_), .A2(new_n435_), .ZN(new_n436_));
  OAI21_X1  g235(.A(KEYINPUT21), .B1(new_n433_), .B2(KEYINPUT90), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  OAI211_X1 g237(.A(KEYINPUT21), .B(new_n435_), .C1(new_n433_), .C2(KEYINPUT90), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n438_), .A2(new_n439_), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n432_), .A2(new_n440_), .ZN(new_n441_));
  NOR3_X1   g240(.A1(new_n369_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n429_), .B1(new_n441_), .B2(new_n442_), .ZN(new_n443_));
  AOI21_X1  g242(.A(new_n429_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n367_), .A2(new_n370_), .ZN(new_n445_));
  OAI21_X1  g244(.A(new_n444_), .B1(new_n445_), .B2(new_n431_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n443_), .A2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n431_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n449_), .A2(KEYINPUT28), .ZN(new_n450_));
  INV_X1    g249(.A(KEYINPUT28), .ZN(new_n451_));
  OAI211_X1 g250(.A(new_n451_), .B(new_n431_), .C1(new_n353_), .C2(new_n354_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(G22gat), .B(G50gat), .ZN(new_n453_));
  INV_X1    g252(.A(new_n453_), .ZN(new_n454_));
  AND3_X1   g253(.A1(new_n450_), .A2(new_n452_), .A3(new_n454_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n454_), .B1(new_n450_), .B2(new_n452_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G78gat), .B(G106gat), .ZN(new_n457_));
  NOR3_X1   g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(KEYINPUT92), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n451_), .B1(new_n445_), .B2(new_n431_), .ZN(new_n460_));
  INV_X1    g259(.A(new_n452_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n453_), .B1(new_n460_), .B2(new_n461_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n450_), .A2(new_n452_), .A3(new_n454_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n459_), .B1(new_n462_), .B2(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(new_n448_), .B1(new_n458_), .B2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n440_), .A2(new_n417_), .ZN(new_n466_));
  OR2_X1    g265(.A1(G183gat), .A2(G190gat), .ZN(new_n467_));
  NAND3_X1  g266(.A1(new_n400_), .A2(new_n467_), .A3(new_n401_), .ZN(new_n468_));
  OR2_X1    g267(.A1(new_n468_), .A2(KEYINPUT94), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n468_), .A2(KEYINPUT94), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n395_), .A3(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT26), .B(G190gat), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n404_), .A2(new_n472_), .ZN(new_n473_));
  NAND4_X1  g272(.A1(new_n409_), .A2(new_n473_), .A3(new_n414_), .A4(new_n415_), .ZN(new_n474_));
  NAND4_X1  g273(.A1(new_n471_), .A2(new_n438_), .A3(new_n439_), .A4(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(G226gat), .A2(G233gat), .ZN(new_n476_));
  XOR2_X1   g275(.A(new_n476_), .B(KEYINPUT19), .Z(new_n477_));
  NAND4_X1  g276(.A1(new_n466_), .A2(new_n475_), .A3(KEYINPUT20), .A4(new_n477_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT95), .ZN(new_n479_));
  XOR2_X1   g278(.A(new_n477_), .B(KEYINPUT93), .Z(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT20), .B1(new_n440_), .B2(new_n417_), .ZN(new_n481_));
  AOI22_X1  g280(.A1(new_n471_), .A2(new_n474_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n480_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(KEYINPUT20), .ZN(new_n484_));
  AOI21_X1  g283(.A(new_n484_), .B1(new_n440_), .B2(new_n417_), .ZN(new_n485_));
  INV_X1    g284(.A(KEYINPUT95), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(new_n477_), .A4(new_n475_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n479_), .A2(new_n483_), .A3(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G8gat), .B(G36gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT18), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G64gat), .B(G92gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n488_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n492_), .ZN(new_n494_));
  NAND4_X1  g293(.A1(new_n479_), .A2(new_n494_), .A3(new_n483_), .A4(new_n487_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n493_), .A2(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT27), .ZN(new_n497_));
  INV_X1    g296(.A(new_n482_), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n440_), .A2(new_n417_), .ZN(new_n499_));
  INV_X1    g298(.A(new_n480_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n498_), .A2(new_n499_), .A3(KEYINPUT20), .A4(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n485_), .A2(new_n475_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(new_n477_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n497_), .B1(new_n503_), .B2(new_n492_), .ZN(new_n504_));
  AOI22_X1  g303(.A1(new_n496_), .A2(new_n497_), .B1(new_n504_), .B2(new_n495_), .ZN(new_n505_));
  INV_X1    g304(.A(new_n457_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n462_), .A2(new_n506_), .A3(new_n463_), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n455_), .A2(new_n456_), .ZN(new_n508_));
  OAI211_X1 g307(.A(new_n447_), .B(new_n507_), .C1(new_n508_), .C2(new_n459_), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n465_), .A2(new_n505_), .A3(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n510_), .A2(KEYINPUT101), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT101), .ZN(new_n512_));
  NAND4_X1  g311(.A1(new_n465_), .A2(new_n505_), .A3(new_n509_), .A4(new_n512_), .ZN(new_n513_));
  AOI21_X1  g312(.A(new_n428_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n514_));
  AND2_X1   g313(.A1(new_n465_), .A2(new_n509_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT99), .ZN(new_n516_));
  NOR2_X1   g315(.A1(new_n516_), .A2(KEYINPUT33), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n517_), .B1(new_n388_), .B2(new_n391_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n312_), .ZN(new_n519_));
  AOI21_X1  g318(.A(new_n519_), .B1(new_n377_), .B2(new_n379_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n517_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n376_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n382_), .B1(new_n372_), .B2(new_n378_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n312_), .B1(new_n377_), .B2(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n373_), .A2(KEYINPUT100), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT100), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n385_), .A2(new_n526_), .A3(new_n371_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n527_), .A3(new_n382_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n496_), .B1(new_n524_), .B2(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n518_), .A2(new_n522_), .A3(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n494_), .A2(KEYINPUT32), .ZN(new_n531_));
  NOR2_X1   g330(.A1(new_n488_), .A2(new_n531_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n532_), .B1(new_n503_), .B2(new_n531_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n389_), .A2(new_n390_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n519_), .B1(new_n388_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n376_), .A2(new_n520_), .ZN(new_n537_));
  AOI21_X1  g336(.A(new_n534_), .B1(new_n536_), .B2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n515_), .B1(new_n530_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n465_), .A2(new_n509_), .ZN(new_n540_));
  NAND3_X1  g339(.A1(new_n393_), .A2(new_n540_), .A3(new_n505_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(new_n541_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n427_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n514_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT74), .ZN(new_n545_));
  INV_X1    g344(.A(G29gat), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n546_), .A2(G36gat), .ZN(new_n547_));
  INV_X1    g346(.A(G36gat), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n548_), .A2(G29gat), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n545_), .B1(new_n547_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(G29gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n546_), .A2(G36gat), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n551_), .A2(new_n552_), .A3(KEYINPUT74), .ZN(new_n553_));
  XNOR2_X1  g352(.A(G43gat), .B(G50gat), .ZN(new_n554_));
  AND3_X1   g353(.A1(new_n550_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n550_), .B2(new_n553_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G15gat), .B(G22gat), .ZN(new_n559_));
  INV_X1    g358(.A(G1gat), .ZN(new_n560_));
  INV_X1    g359(.A(G8gat), .ZN(new_n561_));
  OAI21_X1  g360(.A(KEYINPUT14), .B1(new_n560_), .B2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n559_), .A2(new_n562_), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G1gat), .B(G8gat), .ZN(new_n564_));
  XNOR2_X1  g363(.A(new_n563_), .B(new_n564_), .ZN(new_n565_));
  OR2_X1    g364(.A1(new_n558_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT81), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n566_), .A2(new_n567_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n566_), .A2(new_n567_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(G229gat), .A2(G233gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n557_), .B(KEYINPUT15), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n572_), .A2(new_n565_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n570_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n558_), .A2(new_n565_), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n575_), .B(KEYINPUT82), .Z(new_n576_));
  AOI21_X1  g375(.A(new_n576_), .B1(new_n569_), .B2(new_n568_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n574_), .B1(new_n577_), .B2(new_n571_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G113gat), .B(G141gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n579_), .B(KEYINPUT83), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G169gat), .B(G197gat), .ZN(new_n581_));
  XOR2_X1   g380(.A(new_n580_), .B(new_n581_), .Z(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n578_), .A2(new_n583_), .ZN(new_n584_));
  OAI211_X1 g383(.A(new_n574_), .B(new_n582_), .C1(new_n577_), .C2(new_n571_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT80), .ZN(new_n588_));
  XOR2_X1   g387(.A(G127gat), .B(G155gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT16), .ZN(new_n590_));
  XNOR2_X1  g389(.A(G183gat), .B(G211gat), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n590_), .B(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n588_), .B1(new_n592_), .B2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(new_n594_), .B(new_n565_), .ZN(new_n595_));
  AND2_X1   g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596_));
  OR2_X1    g395(.A1(new_n595_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n596_), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n256_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n593_), .B2(new_n592_), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n597_), .A2(new_n256_), .A3(new_n598_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT78), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT77), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n288_), .A2(new_n572_), .ZN(new_n606_));
  AOI22_X1  g405(.A1(new_n227_), .A2(new_n231_), .B1(new_n241_), .B2(new_n248_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G232gat), .A2(G233gat), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n608_), .B(KEYINPUT34), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(KEYINPUT72), .B(KEYINPUT35), .Z(new_n611_));
  AOI22_X1  g410(.A1(new_n607_), .A2(new_n557_), .B1(new_n610_), .B2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n606_), .A2(new_n612_), .ZN(new_n613_));
  OR2_X1    g412(.A1(new_n610_), .A2(new_n611_), .ZN(new_n614_));
  XOR2_X1   g413(.A(new_n614_), .B(KEYINPUT73), .Z(new_n615_));
  INV_X1    g414(.A(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n613_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n606_), .A2(new_n612_), .A3(new_n615_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT75), .ZN(new_n621_));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n621_), .B(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT36), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n623_), .A2(new_n624_), .ZN(new_n625_));
  XOR2_X1   g424(.A(new_n625_), .B(KEYINPUT76), .Z(new_n626_));
  AOI21_X1  g425(.A(new_n605_), .B1(new_n619_), .B2(new_n626_), .ZN(new_n627_));
  AND3_X1   g426(.A1(new_n606_), .A2(new_n612_), .A3(new_n615_), .ZN(new_n628_));
  AOI21_X1  g427(.A(new_n615_), .B1(new_n606_), .B2(new_n612_), .ZN(new_n629_));
  OAI211_X1 g428(.A(new_n605_), .B(new_n626_), .C1(new_n628_), .C2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n604_), .B1(new_n627_), .B2(new_n631_), .ZN(new_n632_));
  OAI21_X1  g431(.A(new_n626_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n633_), .A2(KEYINPUT77), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(KEYINPUT78), .A3(new_n630_), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n623_), .B(new_n624_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT79), .Z(new_n637_));
  NAND3_X1  g436(.A1(new_n637_), .A2(new_n618_), .A3(new_n617_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n632_), .A2(new_n635_), .A3(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n639_), .A2(KEYINPUT37), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n619_), .A2(new_n636_), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n641_), .B1(new_n627_), .B2(new_n631_), .ZN(new_n642_));
  OR2_X1    g441(.A1(new_n642_), .A2(KEYINPUT37), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n640_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n603_), .A2(new_n644_), .ZN(new_n645_));
  NOR4_X1   g444(.A1(new_n307_), .A2(new_n544_), .A3(new_n587_), .A4(new_n645_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n393_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n646_), .A2(new_n560_), .A3(new_n647_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT38), .ZN(new_n649_));
  OR2_X1    g448(.A1(new_n648_), .A2(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(new_n642_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n544_), .A2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n306_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n653_), .A2(new_n587_), .A3(new_n602_), .ZN(new_n654_));
  AND2_X1   g453(.A1(new_n652_), .A2(new_n654_), .ZN(new_n655_));
  INV_X1    g454(.A(new_n655_), .ZN(new_n656_));
  OAI21_X1  g455(.A(G1gat), .B1(new_n656_), .B2(new_n393_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n648_), .A2(new_n649_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n650_), .A2(new_n657_), .A3(new_n658_), .ZN(G1324gat));
  OAI21_X1  g458(.A(G8gat), .B1(new_n656_), .B2(new_n505_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n660_), .A2(KEYINPUT102), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT39), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n660_), .A2(KEYINPUT102), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n662_), .A2(new_n663_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT40), .ZN(new_n665_));
  INV_X1    g464(.A(new_n505_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n646_), .A2(new_n561_), .A3(new_n666_), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n667_), .B1(new_n661_), .B2(KEYINPUT39), .ZN(new_n668_));
  OR3_X1    g467(.A1(new_n664_), .A2(new_n665_), .A3(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(new_n665_), .B1(new_n664_), .B2(new_n668_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(G1325gat));
  OAI21_X1  g470(.A(G15gat), .B1(new_n656_), .B2(new_n543_), .ZN(new_n672_));
  XNOR2_X1  g471(.A(KEYINPUT103), .B(KEYINPUT41), .ZN(new_n673_));
  OR2_X1    g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n672_), .A2(new_n673_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n646_), .A2(new_n423_), .A3(new_n427_), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n674_), .A2(new_n675_), .A3(new_n676_), .ZN(G1326gat));
  INV_X1    g476(.A(G22gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n678_), .B1(new_n655_), .B2(new_n540_), .ZN(new_n679_));
  XOR2_X1   g478(.A(new_n679_), .B(KEYINPUT42), .Z(new_n680_));
  NAND2_X1  g479(.A1(new_n540_), .A2(new_n678_), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n681_), .B(KEYINPUT104), .Z(new_n682_));
  NAND2_X1  g481(.A1(new_n646_), .A2(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n680_), .A2(new_n683_), .ZN(G1327gat));
  NOR2_X1   g483(.A1(new_n544_), .A2(new_n587_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n602_), .A2(new_n651_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n653_), .A2(new_n686_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n685_), .A2(new_n687_), .ZN(new_n688_));
  AOI21_X1  g487(.A(G29gat), .B1(new_n688_), .B2(new_n647_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n653_), .A2(new_n603_), .A3(new_n587_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  OAI21_X1  g491(.A(KEYINPUT43), .B1(new_n544_), .B2(new_n644_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n533_), .B1(new_n381_), .B2(new_n392_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n518_), .A2(new_n529_), .A3(new_n522_), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n540_), .B1(new_n694_), .B2(new_n695_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n536_), .A2(new_n537_), .A3(new_n505_), .ZN(new_n697_));
  NOR2_X1   g496(.A1(new_n515_), .A2(new_n697_), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n543_), .B1(new_n696_), .B2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n511_), .A2(new_n513_), .ZN(new_n700_));
  INV_X1    g499(.A(new_n428_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n699_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n704_));
  INV_X1    g503(.A(new_n644_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n703_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n692_), .B1(new_n693_), .B2(new_n706_), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n690_), .B1(new_n707_), .B2(KEYINPUT44), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n704_), .B1(new_n703_), .B2(new_n705_), .ZN(new_n709_));
  AOI211_X1 g508(.A(KEYINPUT43), .B(new_n644_), .C1(new_n699_), .C2(new_n702_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n691_), .B1(new_n709_), .B2(new_n710_), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT44), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(KEYINPUT105), .A3(new_n712_), .ZN(new_n713_));
  AOI22_X1  g512(.A1(new_n708_), .A2(new_n713_), .B1(KEYINPUT44), .B2(new_n707_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n393_), .A2(new_n546_), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n689_), .B1(new_n714_), .B2(new_n715_), .ZN(G1328gat));
  INV_X1    g515(.A(KEYINPUT45), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n505_), .A2(G36gat), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n685_), .A2(new_n687_), .A3(new_n718_), .ZN(new_n719_));
  AND2_X1   g518(.A1(new_n719_), .A2(KEYINPUT107), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n719_), .A2(KEYINPUT107), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n719_), .A2(KEYINPUT107), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n719_), .A2(KEYINPUT107), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n723_), .A2(KEYINPUT45), .A3(new_n724_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n722_), .A2(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n505_), .B1(new_n707_), .B2(KEYINPUT44), .ZN(new_n727_));
  AND3_X1   g526(.A1(new_n711_), .A2(KEYINPUT105), .A3(new_n712_), .ZN(new_n728_));
  AOI21_X1  g527(.A(KEYINPUT105), .B1(new_n711_), .B2(new_n712_), .ZN(new_n729_));
  OAI21_X1  g528(.A(new_n727_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n730_), .A2(G36gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n726_), .B1(new_n731_), .B2(KEYINPUT106), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT108), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT46), .ZN(new_n734_));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n730_), .A2(new_n735_), .A3(G36gat), .ZN(new_n736_));
  NAND4_X1  g535(.A1(new_n732_), .A2(new_n733_), .A3(new_n734_), .A4(new_n736_), .ZN(new_n737_));
  OAI211_X1 g536(.A(KEYINPUT44), .B(new_n691_), .C1(new_n709_), .C2(new_n710_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n738_), .A2(new_n666_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n708_), .B2(new_n713_), .ZN(new_n740_));
  OAI21_X1  g539(.A(KEYINPUT106), .B1(new_n740_), .B2(new_n548_), .ZN(new_n741_));
  AND2_X1   g540(.A1(new_n722_), .A2(new_n725_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n736_), .A3(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n733_), .A2(new_n734_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(KEYINPUT108), .A2(KEYINPUT46), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n743_), .A2(new_n744_), .A3(new_n745_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n737_), .A2(new_n746_), .ZN(G1329gat));
  AOI21_X1  g546(.A(G43gat), .B1(new_n688_), .B2(new_n427_), .ZN(new_n748_));
  INV_X1    g547(.A(G43gat), .ZN(new_n749_));
  NOR2_X1   g548(.A1(new_n543_), .A2(new_n749_), .ZN(new_n750_));
  AOI21_X1  g549(.A(new_n748_), .B1(new_n714_), .B2(new_n750_), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n751_), .B(KEYINPUT47), .Z(G1330gat));
  NAND2_X1  g551(.A1(new_n714_), .A2(new_n540_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(G50gat), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n515_), .A2(G50gat), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT109), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n688_), .A2(new_n756_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n754_), .A2(new_n757_), .ZN(G1331gat));
  NOR4_X1   g557(.A1(new_n544_), .A2(new_n645_), .A3(new_n586_), .A4(new_n306_), .ZN(new_n759_));
  INV_X1    g558(.A(G57gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(new_n647_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n602_), .A2(new_n586_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n652_), .A2(new_n307_), .A3(new_n762_), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n763_), .A2(new_n647_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n761_), .B1(new_n764_), .B2(new_n760_), .ZN(G1332gat));
  INV_X1    g564(.A(G64gat), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n763_), .B2(new_n666_), .ZN(new_n767_));
  XOR2_X1   g566(.A(new_n767_), .B(KEYINPUT48), .Z(new_n768_));
  NAND3_X1  g567(.A1(new_n759_), .A2(new_n766_), .A3(new_n666_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n768_), .A2(new_n769_), .ZN(G1333gat));
  INV_X1    g569(.A(G71gat), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n759_), .A2(new_n771_), .A3(new_n427_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n763_), .A2(new_n427_), .ZN(new_n773_));
  XOR2_X1   g572(.A(KEYINPUT110), .B(KEYINPUT49), .Z(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(G71gat), .A3(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(G71gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(G1334gat));
  INV_X1    g576(.A(G78gat), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n778_), .B1(new_n763_), .B2(new_n540_), .ZN(new_n779_));
  XOR2_X1   g578(.A(new_n779_), .B(KEYINPUT50), .Z(new_n780_));
  NAND3_X1  g579(.A1(new_n759_), .A2(new_n778_), .A3(new_n540_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(G1335gat));
  INV_X1    g581(.A(new_n307_), .ZN(new_n783_));
  NOR4_X1   g582(.A1(new_n783_), .A2(new_n544_), .A3(new_n586_), .A4(new_n686_), .ZN(new_n784_));
  AOI21_X1  g583(.A(G85gat), .B1(new_n784_), .B2(new_n647_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n693_), .A2(new_n706_), .ZN(new_n786_));
  NOR3_X1   g585(.A1(new_n603_), .A2(new_n306_), .A3(new_n586_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  XNOR2_X1  g587(.A(new_n788_), .B(KEYINPUT111), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n647_), .A2(new_n236_), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n790_), .B(KEYINPUT112), .Z(new_n791_));
  AOI21_X1  g590(.A(new_n785_), .B1(new_n789_), .B2(new_n791_), .ZN(G1336gat));
  NAND3_X1  g591(.A1(new_n784_), .A2(new_n222_), .A3(new_n666_), .ZN(new_n793_));
  AND2_X1   g592(.A1(new_n789_), .A2(new_n666_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n793_), .B1(new_n794_), .B2(new_n222_), .ZN(G1337gat));
  OAI211_X1 g594(.A(new_n784_), .B(new_n427_), .C1(new_n246_), .C2(new_n247_), .ZN(new_n796_));
  XOR2_X1   g595(.A(new_n796_), .B(KEYINPUT113), .Z(new_n797_));
  OAI21_X1  g596(.A(G99gat), .B1(new_n788_), .B2(new_n543_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT51), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT51), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n797_), .A2(new_n801_), .A3(new_n798_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n800_), .A2(new_n802_), .ZN(G1338gat));
  NAND3_X1  g602(.A1(new_n784_), .A2(new_n205_), .A3(new_n540_), .ZN(new_n804_));
  OAI21_X1  g603(.A(G106gat), .B1(new_n788_), .B2(new_n515_), .ZN(new_n805_));
  AND2_X1   g604(.A1(new_n805_), .A2(KEYINPUT52), .ZN(new_n806_));
  NOR2_X1   g605(.A1(new_n805_), .A2(KEYINPUT52), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n804_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n808_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g608(.A1(new_n762_), .A2(new_n306_), .A3(new_n644_), .ZN(new_n810_));
  XNOR2_X1  g609(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  OR2_X1    g611(.A1(new_n810_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n810_), .A2(new_n812_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n301_), .A2(new_n303_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n571_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n570_), .A2(new_n817_), .A3(new_n573_), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n818_), .B(new_n583_), .C1(new_n577_), .C2(new_n817_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n585_), .A2(new_n819_), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n816_), .A2(KEYINPUT117), .A3(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT117), .B1(new_n816_), .B2(new_n820_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824_));
  NAND2_X1  g623(.A1(new_n290_), .A2(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(KEYINPUT115), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT115), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n290_), .A2(new_n827_), .A3(new_n824_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n263_), .A2(new_n289_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(G230gat), .A3(G233gat), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n826_), .A2(new_n828_), .A3(new_n830_), .ZN(new_n831_));
  NAND4_X1  g630(.A1(new_n263_), .A2(KEYINPUT55), .A3(new_n264_), .A4(new_n289_), .ZN(new_n832_));
  XNOR2_X1  g631(.A(new_n832_), .B(KEYINPUT116), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n296_), .B1(new_n831_), .B2(new_n833_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n299_), .B1(new_n834_), .B2(KEYINPUT56), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT56), .ZN(new_n836_));
  OAI211_X1 g635(.A(new_n836_), .B(new_n296_), .C1(new_n831_), .C2(new_n833_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n835_), .A2(new_n586_), .A3(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n651_), .B1(new_n823_), .B2(new_n838_), .ZN(new_n839_));
  OR2_X1    g638(.A1(new_n839_), .A2(KEYINPUT57), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n835_), .A2(new_n837_), .A3(new_n820_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n841_), .A2(new_n842_), .ZN(new_n843_));
  NAND4_X1  g642(.A1(new_n835_), .A2(KEYINPUT58), .A3(new_n837_), .A4(new_n820_), .ZN(new_n844_));
  NAND3_X1  g643(.A1(new_n843_), .A2(new_n705_), .A3(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n839_), .A2(KEYINPUT57), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n840_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n815_), .B1(new_n847_), .B2(new_n602_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n700_), .A2(new_n427_), .A3(new_n647_), .ZN(new_n849_));
  NOR3_X1   g648(.A1(new_n848_), .A2(KEYINPUT59), .A3(new_n849_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n845_), .A2(new_n851_), .ZN(new_n852_));
  NAND4_X1  g651(.A1(new_n843_), .A2(KEYINPUT118), .A3(new_n705_), .A4(new_n844_), .ZN(new_n853_));
  NAND4_X1  g652(.A1(new_n840_), .A2(new_n852_), .A3(new_n853_), .A4(new_n846_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n815_), .B1(new_n854_), .B2(new_n602_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n855_), .A2(new_n849_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n850_), .B1(new_n856_), .B2(KEYINPUT59), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n586_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G113gat), .ZN(new_n859_));
  OR2_X1    g658(.A1(new_n856_), .A2(KEYINPUT119), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n856_), .A2(KEYINPUT119), .ZN(new_n861_));
  NOR2_X1   g660(.A1(new_n587_), .A2(G113gat), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n860_), .A2(new_n861_), .A3(new_n862_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n859_), .A2(new_n863_), .ZN(G1340gat));
  NAND2_X1  g663(.A1(new_n857_), .A2(new_n307_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(G120gat), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n306_), .A2(KEYINPUT60), .ZN(new_n867_));
  MUX2_X1   g666(.A(new_n867_), .B(KEYINPUT60), .S(G120gat), .Z(new_n868_));
  NAND3_X1  g667(.A1(new_n860_), .A2(new_n861_), .A3(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n866_), .A2(new_n869_), .ZN(G1341gat));
  NAND2_X1  g669(.A1(new_n857_), .A2(new_n603_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(G127gat), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n602_), .A2(G127gat), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n860_), .A2(new_n861_), .A3(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n874_), .ZN(G1342gat));
  NAND3_X1  g674(.A1(new_n860_), .A2(new_n651_), .A3(new_n861_), .ZN(new_n876_));
  INV_X1    g675(.A(G134gat), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT120), .B(G134gat), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n644_), .A2(new_n878_), .ZN(new_n879_));
  AOI22_X1  g678(.A1(new_n876_), .A2(new_n877_), .B1(new_n857_), .B2(new_n879_), .ZN(G1343gat));
  NOR2_X1   g679(.A1(new_n515_), .A2(new_n427_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n854_), .A2(new_n602_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n815_), .ZN(new_n884_));
  AOI21_X1  g683(.A(new_n882_), .B1(new_n883_), .B2(new_n884_), .ZN(new_n885_));
  NOR2_X1   g684(.A1(new_n393_), .A2(new_n666_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n885_), .A2(new_n886_), .ZN(new_n887_));
  AND2_X1   g686(.A1(new_n887_), .A2(new_n586_), .ZN(new_n888_));
  XNOR2_X1  g687(.A(KEYINPUT121), .B(G141gat), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n888_), .B(new_n889_), .ZN(G1344gat));
  AND2_X1   g689(.A1(new_n887_), .A2(new_n307_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(KEYINPUT122), .B(G148gat), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n891_), .B(new_n892_), .ZN(G1345gat));
  NAND3_X1  g692(.A1(new_n885_), .A2(new_n603_), .A3(new_n886_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n894_), .A2(new_n895_), .ZN(new_n896_));
  NAND4_X1  g695(.A1(new_n885_), .A2(KEYINPUT123), .A3(new_n603_), .A4(new_n886_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(KEYINPUT61), .B(G155gat), .ZN(new_n898_));
  AND3_X1   g697(.A1(new_n896_), .A2(new_n897_), .A3(new_n898_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n898_), .B1(new_n896_), .B2(new_n897_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n899_), .A2(new_n900_), .ZN(G1346gat));
  INV_X1    g700(.A(G162gat), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n887_), .A2(new_n902_), .A3(new_n651_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n887_), .A2(new_n705_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n903_), .B1(new_n904_), .B2(new_n902_), .ZN(G1347gat));
  XNOR2_X1  g704(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n906_));
  INV_X1    g705(.A(new_n906_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n848_), .A2(new_n540_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n393_), .A2(new_n666_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n909_), .A2(new_n543_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n908_), .A2(new_n586_), .A3(new_n910_), .ZN(new_n911_));
  OAI211_X1 g710(.A(G169gat), .B(new_n907_), .C1(new_n911_), .C2(KEYINPUT22), .ZN(new_n912_));
  INV_X1    g711(.A(new_n911_), .ZN(new_n913_));
  INV_X1    g712(.A(KEYINPUT22), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n906_), .B1(new_n913_), .B2(new_n914_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n412_), .B1(new_n913_), .B2(new_n906_), .ZN(new_n916_));
  OAI21_X1  g715(.A(new_n912_), .B1(new_n915_), .B2(new_n916_), .ZN(G1348gat));
  NAND3_X1  g716(.A1(new_n908_), .A2(new_n653_), .A3(new_n910_), .ZN(new_n918_));
  NOR2_X1   g717(.A1(new_n855_), .A2(new_n540_), .ZN(new_n919_));
  INV_X1    g718(.A(new_n910_), .ZN(new_n920_));
  NOR3_X1   g719(.A1(new_n783_), .A2(new_n413_), .A3(new_n920_), .ZN(new_n921_));
  AOI22_X1  g720(.A1(new_n918_), .A2(new_n413_), .B1(new_n919_), .B2(new_n921_), .ZN(G1349gat));
  NOR2_X1   g721(.A1(new_n920_), .A2(new_n602_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n405_), .ZN(new_n924_));
  INV_X1    g723(.A(new_n924_), .ZN(new_n925_));
  AND3_X1   g724(.A1(new_n908_), .A2(KEYINPUT125), .A3(new_n925_), .ZN(new_n926_));
  AOI21_X1  g725(.A(G183gat), .B1(new_n919_), .B2(new_n923_), .ZN(new_n927_));
  AOI21_X1  g726(.A(KEYINPUT125), .B1(new_n908_), .B2(new_n925_), .ZN(new_n928_));
  NOR3_X1   g727(.A1(new_n926_), .A2(new_n927_), .A3(new_n928_), .ZN(G1350gat));
  NAND2_X1  g728(.A1(new_n908_), .A2(new_n910_), .ZN(new_n930_));
  OAI21_X1  g729(.A(G190gat), .B1(new_n930_), .B2(new_n644_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n651_), .A2(new_n472_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n930_), .B2(new_n932_), .ZN(G1351gat));
  XNOR2_X1  g732(.A(KEYINPUT127), .B(G197gat), .ZN(new_n934_));
  INV_X1    g733(.A(new_n909_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n885_), .A2(new_n935_), .ZN(new_n936_));
  NAND2_X1  g735(.A1(new_n936_), .A2(KEYINPUT126), .ZN(new_n937_));
  INV_X1    g736(.A(KEYINPUT126), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n885_), .A2(new_n938_), .A3(new_n935_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n937_), .A2(new_n939_), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n934_), .B1(new_n940_), .B2(new_n586_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n938_), .B1(new_n885_), .B2(new_n935_), .ZN(new_n942_));
  NOR4_X1   g741(.A1(new_n855_), .A2(KEYINPUT126), .A3(new_n882_), .A4(new_n909_), .ZN(new_n943_));
  OAI211_X1 g742(.A(new_n586_), .B(new_n934_), .C1(new_n942_), .C2(new_n943_), .ZN(new_n944_));
  INV_X1    g743(.A(new_n944_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n941_), .A2(new_n945_), .ZN(G1352gat));
  OAI21_X1  g745(.A(new_n307_), .B1(new_n942_), .B2(new_n943_), .ZN(new_n947_));
  XNOR2_X1  g746(.A(new_n947_), .B(G204gat), .ZN(G1353gat));
  OR2_X1    g747(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n949_), .B1(new_n940_), .B2(new_n603_), .ZN(new_n950_));
  XOR2_X1   g749(.A(KEYINPUT63), .B(G211gat), .Z(new_n951_));
  OAI211_X1 g750(.A(new_n603_), .B(new_n951_), .C1(new_n942_), .C2(new_n943_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(new_n953_));
  NOR2_X1   g752(.A1(new_n950_), .A2(new_n953_), .ZN(G1354gat));
  INV_X1    g753(.A(G218gat), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n940_), .A2(new_n955_), .A3(new_n651_), .ZN(new_n956_));
  AOI21_X1  g755(.A(new_n644_), .B1(new_n937_), .B2(new_n939_), .ZN(new_n957_));
  OAI21_X1  g756(.A(new_n956_), .B1(new_n955_), .B2(new_n957_), .ZN(G1355gat));
endmodule


