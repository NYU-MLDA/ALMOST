//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:42 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n699_, new_n700_,
    new_n701_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n745_, new_n746_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n864_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n872_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n893_, new_n894_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n920_, new_n921_, new_n922_, new_n923_,
    new_n924_, new_n925_, new_n926_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n944_, new_n945_;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G169gat), .ZN(new_n202_));
  INV_X1    g001(.A(G176gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n204_), .A2(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(G183gat), .ZN(new_n207_));
  INV_X1    g006(.A(G190gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT23), .B1(new_n207_), .B2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT81), .ZN(new_n210_));
  OR3_X1    g009(.A1(new_n207_), .A2(new_n208_), .A3(KEYINPUT23), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n210_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n207_), .A2(new_n208_), .ZN(new_n213_));
  AOI21_X1  g012(.A(new_n206_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n214_));
  XNOR2_X1  g013(.A(KEYINPUT25), .B(G183gat), .ZN(new_n215_));
  XNOR2_X1  g014(.A(KEYINPUT26), .B(G190gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  OR2_X1    g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(KEYINPUT24), .A3(new_n205_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n218_), .A2(KEYINPUT24), .ZN(new_n220_));
  AND3_X1   g019(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n211_), .A2(new_n209_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n214_), .A2(new_n223_), .ZN(new_n224_));
  XOR2_X1   g023(.A(G197gat), .B(G204gat), .Z(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT21), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G211gat), .B(G218gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(G197gat), .B(G204gat), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT21), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n226_), .A2(new_n227_), .A3(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT89), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OR3_X1    g032(.A1(new_n228_), .A2(new_n227_), .A3(new_n229_), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n232_), .B1(new_n231_), .B2(new_n234_), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n233_), .A2(new_n235_), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT20), .B1(new_n224_), .B2(new_n236_), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT92), .ZN(new_n238_));
  AOI22_X1  g037(.A1(new_n206_), .A2(KEYINPUT82), .B1(new_n222_), .B2(new_n213_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n239_), .B1(KEYINPUT82), .B2(new_n206_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n212_), .A2(new_n221_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(new_n233_), .A2(new_n235_), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n238_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n236_), .A2(new_n242_), .A3(KEYINPUT92), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n237_), .B1(new_n245_), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G226gat), .A2(G233gat), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  OR2_X1    g049(.A1(new_n247_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT95), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n251_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n224_), .A2(KEYINPUT91), .A3(new_n236_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n243_), .A2(new_n244_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT91), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n214_), .A2(new_n223_), .ZN(new_n257_));
  OAI21_X1  g056(.A(new_n256_), .B1(new_n257_), .B2(new_n244_), .ZN(new_n258_));
  NAND4_X1  g057(.A1(new_n254_), .A2(new_n255_), .A3(new_n258_), .A4(KEYINPUT20), .ZN(new_n259_));
  INV_X1    g058(.A(new_n250_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  NOR2_X1   g060(.A1(new_n247_), .A2(new_n250_), .ZN(new_n262_));
  AOI21_X1  g061(.A(new_n261_), .B1(new_n262_), .B2(KEYINPUT95), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n253_), .A2(new_n263_), .ZN(new_n264_));
  XNOR2_X1  g063(.A(G8gat), .B(G36gat), .ZN(new_n265_));
  INV_X1    g064(.A(G92gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n265_), .B(new_n266_), .ZN(new_n267_));
  XNOR2_X1  g066(.A(KEYINPUT18), .B(G64gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(new_n268_), .Z(new_n269_));
  NAND2_X1  g068(.A1(new_n264_), .A2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n247_), .A2(new_n250_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n269_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n259_), .A2(new_n260_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n271_), .A2(new_n272_), .A3(new_n273_), .ZN(new_n274_));
  AND2_X1   g073(.A1(new_n274_), .A2(KEYINPUT27), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT27), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n271_), .A2(new_n273_), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n277_), .A2(new_n269_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n278_), .A2(new_n274_), .ZN(new_n279_));
  AOI22_X1  g078(.A1(new_n270_), .A2(new_n275_), .B1(new_n276_), .B2(new_n279_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G225gat), .A2(G233gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G113gat), .B(G120gat), .ZN(new_n283_));
  XNOR2_X1  g082(.A(new_n283_), .B(KEYINPUT85), .ZN(new_n284_));
  XNOR2_X1  g083(.A(G127gat), .B(G134gat), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n284_), .B(new_n285_), .ZN(new_n286_));
  AND2_X1   g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287_));
  NOR2_X1   g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  NOR2_X1   g088(.A1(G141gat), .A2(G148gat), .ZN(new_n290_));
  XOR2_X1   g089(.A(new_n290_), .B(KEYINPUT3), .Z(new_n291_));
  NAND2_X1  g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292_));
  XOR2_X1   g091(.A(new_n292_), .B(KEYINPUT2), .Z(new_n293_));
  OAI21_X1  g092(.A(new_n289_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT1), .ZN(new_n295_));
  AOI21_X1  g094(.A(new_n288_), .B1(new_n287_), .B2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n296_), .B1(new_n295_), .B2(new_n287_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n290_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n297_), .A2(new_n298_), .A3(new_n292_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n294_), .A2(new_n299_), .ZN(new_n300_));
  NOR2_X1   g099(.A1(new_n300_), .A2(KEYINPUT86), .ZN(new_n301_));
  INV_X1    g100(.A(KEYINPUT86), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n302_), .B1(new_n294_), .B2(new_n299_), .ZN(new_n303_));
  OAI21_X1  g102(.A(new_n286_), .B1(new_n301_), .B2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(KEYINPUT4), .ZN(new_n305_));
  AND2_X1   g104(.A1(new_n304_), .A2(new_n305_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n286_), .A2(new_n300_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n305_), .B1(new_n304_), .B2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n282_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT93), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  OAI211_X1 g110(.A(KEYINPUT93), .B(new_n282_), .C1(new_n306_), .C2(new_n308_), .ZN(new_n312_));
  AND2_X1   g111(.A1(new_n304_), .A2(new_n307_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n313_), .A2(new_n281_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G1gat), .B(G29gat), .ZN(new_n316_));
  INV_X1    g115(.A(G85gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(KEYINPUT0), .B(G57gat), .ZN(new_n319_));
  XOR2_X1   g118(.A(new_n318_), .B(new_n319_), .Z(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n320_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n311_), .A2(new_n322_), .A3(new_n312_), .A4(new_n314_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n321_), .A2(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G22gat), .B(G50gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT28), .ZN(new_n327_));
  INV_X1    g126(.A(G233gat), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT88), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n329_), .A2(G228gat), .ZN(new_n330_));
  INV_X1    g129(.A(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n329_), .A2(G228gat), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n328_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n236_), .A2(new_n334_), .ZN(new_n335_));
  OR2_X1    g134(.A1(new_n301_), .A2(new_n303_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n335_), .B1(new_n336_), .B2(KEYINPUT29), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n300_), .A2(KEYINPUT29), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n334_), .B1(new_n236_), .B2(new_n338_), .ZN(new_n339_));
  OAI21_X1  g138(.A(G78gat), .B1(new_n337_), .B2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G78gat), .ZN(new_n341_));
  INV_X1    g140(.A(new_n339_), .ZN(new_n342_));
  NOR2_X1   g141(.A1(new_n301_), .A2(new_n303_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT29), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  OAI211_X1 g144(.A(new_n341_), .B(new_n342_), .C1(new_n345_), .C2(new_n335_), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n340_), .A2(G106gat), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT87), .ZN(new_n348_));
  AOI21_X1  g147(.A(G106gat), .B1(new_n340_), .B2(new_n346_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n327_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n340_), .A2(new_n346_), .ZN(new_n351_));
  INV_X1    g150(.A(G106gat), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n327_), .ZN(new_n354_));
  NAND4_X1  g153(.A1(new_n353_), .A2(KEYINPUT87), .A3(new_n354_), .A4(new_n347_), .ZN(new_n355_));
  NOR2_X1   g154(.A1(new_n336_), .A2(KEYINPUT29), .ZN(new_n356_));
  NAND3_X1  g155(.A1(new_n350_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n356_), .B1(new_n350_), .B2(new_n355_), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n280_), .B(new_n325_), .C1(new_n358_), .C2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT33), .ZN(new_n361_));
  AND2_X1   g160(.A1(new_n323_), .A2(new_n361_), .ZN(new_n362_));
  OAI21_X1  g161(.A(new_n281_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n363_));
  AOI21_X1  g162(.A(new_n322_), .B1(new_n313_), .B2(new_n282_), .ZN(new_n364_));
  AND2_X1   g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  NOR3_X1   g164(.A1(new_n362_), .A2(new_n279_), .A3(new_n365_), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n323_), .A2(new_n361_), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n272_), .A2(KEYINPUT32), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  OAI21_X1  g168(.A(KEYINPUT94), .B1(new_n277_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT94), .ZN(new_n371_));
  NAND4_X1  g170(.A1(new_n271_), .A2(new_n371_), .A3(new_n273_), .A4(new_n368_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n370_), .A2(new_n372_), .ZN(new_n373_));
  AOI21_X1  g172(.A(new_n368_), .B1(new_n253_), .B2(new_n263_), .ZN(new_n374_));
  NOR2_X1   g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  AOI22_X1  g174(.A1(new_n366_), .A2(new_n367_), .B1(new_n375_), .B2(new_n324_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n359_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n357_), .ZN(new_n378_));
  OAI21_X1  g177(.A(new_n360_), .B1(new_n376_), .B2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G227gat), .A2(G233gat), .ZN(new_n380_));
  INV_X1    g179(.A(new_n380_), .ZN(new_n381_));
  XNOR2_X1  g180(.A(new_n286_), .B(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G71gat), .B(G99gat), .ZN(new_n383_));
  XNOR2_X1  g182(.A(new_n382_), .B(new_n383_), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT84), .B(G15gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n383_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n382_), .B(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n385_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n388_), .A2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n386_), .A2(new_n390_), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n242_), .B(KEYINPUT30), .Z(new_n392_));
  XNOR2_X1  g191(.A(KEYINPUT83), .B(G43gat), .ZN(new_n393_));
  XNOR2_X1  g192(.A(new_n393_), .B(KEYINPUT31), .ZN(new_n394_));
  INV_X1    g193(.A(new_n394_), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n392_), .B(new_n395_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n391_), .A2(new_n396_), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n392_), .B(new_n394_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n398_), .A2(new_n390_), .A3(new_n386_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n397_), .A2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NOR2_X1   g200(.A1(new_n401_), .A2(new_n324_), .ZN(new_n402_));
  NAND4_X1  g201(.A1(new_n377_), .A2(new_n402_), .A3(new_n280_), .A4(new_n357_), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT96), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n403_), .A2(new_n404_), .ZN(new_n405_));
  NOR2_X1   g204(.A1(new_n358_), .A2(new_n359_), .ZN(new_n406_));
  NAND4_X1  g205(.A1(new_n406_), .A2(KEYINPUT96), .A3(new_n280_), .A4(new_n402_), .ZN(new_n407_));
  AOI22_X1  g206(.A1(new_n379_), .A2(new_n401_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(KEYINPUT10), .B(G99gat), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT65), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n409_), .A2(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT10), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n412_), .A2(G99gat), .ZN(new_n413_));
  INV_X1    g212(.A(G99gat), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n414_), .A2(KEYINPUT10), .ZN(new_n415_));
  OAI21_X1  g214(.A(KEYINPUT65), .B1(new_n413_), .B2(new_n415_), .ZN(new_n416_));
  AOI21_X1  g215(.A(G106gat), .B1(new_n411_), .B2(new_n416_), .ZN(new_n417_));
  NOR2_X1   g216(.A1(G85gat), .A2(G92gat), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(G85gat), .A2(G92gat), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n419_), .A2(KEYINPUT9), .A3(new_n420_), .ZN(new_n421_));
  AND3_X1   g220(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n422_));
  AOI21_X1  g221(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n423_));
  NOR2_X1   g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  OR2_X1    g223(.A1(new_n420_), .A2(KEYINPUT9), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n421_), .A2(new_n424_), .A3(new_n425_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n417_), .A2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NOR3_X1   g228(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n430_));
  NOR2_X1   g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G99gat), .A2(G106gat), .ZN(new_n432_));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n434_), .A2(KEYINPUT67), .A3(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT67), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n431_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(new_n420_), .ZN(new_n440_));
  NOR2_X1   g239(.A1(new_n440_), .A2(new_n418_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n439_), .A2(new_n441_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n442_), .A2(KEYINPUT8), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT7), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n444_), .A2(new_n414_), .A3(new_n352_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n445_), .A2(new_n434_), .A3(new_n435_), .A4(new_n428_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT66), .ZN(new_n447_));
  NOR3_X1   g246(.A1(new_n440_), .A2(new_n418_), .A3(KEYINPUT8), .ZN(new_n448_));
  AND3_X1   g247(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n447_), .B1(new_n446_), .B2(new_n448_), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n427_), .B1(new_n443_), .B2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G29gat), .B(G36gat), .Z(new_n453_));
  XNOR2_X1  g252(.A(G43gat), .B(G50gat), .ZN(new_n454_));
  OR2_X1    g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n453_), .A2(new_n454_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n455_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT35), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G232gat), .A2(G233gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n460_), .B(new_n461_), .ZN(new_n462_));
  AOI22_X1  g261(.A1(new_n452_), .A2(new_n458_), .B1(new_n459_), .B2(new_n462_), .ZN(new_n463_));
  NOR2_X1   g262(.A1(new_n409_), .A2(new_n410_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n413_), .A2(new_n415_), .A3(KEYINPUT65), .ZN(new_n465_));
  OAI21_X1  g264(.A(new_n352_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT71), .ZN(new_n467_));
  INV_X1    g266(.A(new_n426_), .ZN(new_n468_));
  NAND3_X1  g267(.A1(new_n466_), .A2(new_n467_), .A3(new_n468_), .ZN(new_n469_));
  OAI21_X1  g268(.A(KEYINPUT71), .B1(new_n417_), .B2(new_n426_), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT70), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n446_), .A2(new_n448_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(KEYINPUT66), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n446_), .A2(new_n447_), .A3(new_n448_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n474_), .A2(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n477_), .B1(new_n439_), .B2(new_n441_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n472_), .B1(new_n476_), .B2(new_n478_), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n443_), .A2(new_n451_), .A3(KEYINPUT70), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n471_), .B1(new_n479_), .B2(new_n480_), .ZN(new_n481_));
  XNOR2_X1  g280(.A(new_n457_), .B(KEYINPUT15), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n463_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(new_n462_), .A2(new_n459_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  OAI221_X1 g284(.A(new_n463_), .B1(new_n459_), .B2(new_n462_), .C1(new_n481_), .C2(new_n482_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n485_), .A2(new_n486_), .A3(KEYINPUT75), .ZN(new_n487_));
  XNOR2_X1  g286(.A(G190gat), .B(G218gat), .ZN(new_n488_));
  XNOR2_X1  g287(.A(G134gat), .B(G162gat), .ZN(new_n489_));
  XOR2_X1   g288(.A(new_n488_), .B(new_n489_), .Z(new_n490_));
  INV_X1    g289(.A(KEYINPUT36), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n490_), .A2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n487_), .A2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n485_), .A2(new_n486_), .ZN(new_n495_));
  INV_X1    g294(.A(new_n490_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(KEYINPUT36), .A3(new_n496_), .ZN(new_n497_));
  NAND4_X1  g296(.A1(new_n485_), .A2(new_n486_), .A3(KEYINPUT75), .A4(new_n492_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n494_), .A2(new_n497_), .A3(new_n498_), .ZN(new_n499_));
  INV_X1    g298(.A(KEYINPUT37), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n499_), .A2(new_n500_), .ZN(new_n501_));
  NAND4_X1  g300(.A1(new_n494_), .A2(new_n497_), .A3(KEYINPUT37), .A4(new_n498_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NOR2_X1   g303(.A1(G57gat), .A2(G64gat), .ZN(new_n505_));
  INV_X1    g304(.A(new_n505_), .ZN(new_n506_));
  NAND2_X1  g305(.A1(G57gat), .A2(G64gat), .ZN(new_n507_));
  AOI21_X1  g306(.A(KEYINPUT69), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n507_), .ZN(new_n509_));
  INV_X1    g308(.A(KEYINPUT69), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n509_), .A2(new_n505_), .A3(new_n510_), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT11), .B1(new_n508_), .B2(new_n511_), .ZN(new_n512_));
  OR2_X1    g311(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(KEYINPUT68), .A2(G71gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n515_), .A2(G78gat), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n513_), .A2(new_n341_), .A3(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(new_n506_), .A2(KEYINPUT69), .A3(new_n507_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n510_), .B1(new_n509_), .B2(new_n505_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT11), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n519_), .A2(new_n520_), .A3(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n512_), .A2(new_n518_), .A3(new_n522_), .ZN(new_n523_));
  AOI21_X1  g322(.A(new_n521_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n524_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n523_), .A2(new_n525_), .ZN(new_n526_));
  XNOR2_X1  g325(.A(G15gat), .B(G22gat), .ZN(new_n527_));
  INV_X1    g326(.A(G1gat), .ZN(new_n528_));
  INV_X1    g327(.A(G8gat), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT14), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G1gat), .B(G8gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n526_), .B(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(G231gat), .A2(G233gat), .ZN(new_n535_));
  OR2_X1    g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n534_), .A2(new_n535_), .ZN(new_n537_));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n538_));
  XOR2_X1   g337(.A(KEYINPUT76), .B(KEYINPUT16), .Z(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(G211gat), .ZN(new_n540_));
  XOR2_X1   g339(.A(G127gat), .B(G155gat), .Z(new_n541_));
  XNOR2_X1  g340(.A(new_n540_), .B(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT77), .B(G183gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  OAI211_X1 g343(.A(new_n536_), .B(new_n537_), .C1(new_n538_), .C2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(KEYINPUT17), .ZN(new_n546_));
  AND2_X1   g345(.A1(new_n536_), .A2(new_n537_), .ZN(new_n547_));
  OAI21_X1  g346(.A(new_n545_), .B1(new_n546_), .B2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(new_n548_), .B(KEYINPUT78), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n504_), .A2(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n551_), .B(KEYINPUT79), .ZN(new_n552_));
  NOR2_X1   g351(.A1(new_n408_), .A2(new_n552_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n533_), .A2(new_n457_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n482_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n554_), .B1(new_n555_), .B2(new_n533_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(G229gat), .A2(G233gat), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n556_), .A2(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n533_), .B(new_n457_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(G229gat), .A3(G233gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G113gat), .B(G141gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G169gat), .B(G197gat), .ZN(new_n562_));
  XNOR2_X1  g361(.A(new_n561_), .B(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n558_), .A2(new_n560_), .A3(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n565_), .A2(KEYINPUT80), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n558_), .A2(new_n560_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(new_n563_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n566_), .B(new_n568_), .ZN(new_n569_));
  INV_X1    g368(.A(new_n471_), .ZN(new_n570_));
  NOR3_X1   g369(.A1(new_n476_), .A2(new_n478_), .A3(new_n472_), .ZN(new_n571_));
  AOI21_X1  g370(.A(KEYINPUT70), .B1(new_n443_), .B2(new_n451_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n570_), .B1(new_n571_), .B2(new_n572_), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT12), .ZN(new_n574_));
  NOR2_X1   g373(.A1(new_n526_), .A2(new_n574_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n573_), .A2(new_n575_), .ZN(new_n576_));
  OAI22_X1  g375(.A1(new_n476_), .A2(new_n478_), .B1(new_n417_), .B2(new_n426_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n523_), .A2(new_n525_), .ZN(new_n578_));
  AOI21_X1  g377(.A(KEYINPUT12), .B1(new_n577_), .B2(new_n578_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n577_), .A2(new_n578_), .ZN(new_n580_));
  NOR2_X1   g379(.A1(new_n579_), .A2(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(G230gat), .A2(G233gat), .ZN(new_n582_));
  XOR2_X1   g381(.A(new_n582_), .B(KEYINPUT64), .Z(new_n583_));
  INV_X1    g382(.A(new_n583_), .ZN(new_n584_));
  NAND3_X1  g383(.A1(new_n576_), .A2(new_n581_), .A3(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n452_), .A2(new_n526_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n583_), .B1(new_n586_), .B2(new_n580_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  XOR2_X1   g387(.A(G120gat), .B(G148gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(G204gat), .ZN(new_n590_));
  XNOR2_X1  g389(.A(KEYINPUT5), .B(G176gat), .ZN(new_n591_));
  XOR2_X1   g390(.A(new_n590_), .B(new_n591_), .Z(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n588_), .A2(new_n593_), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n585_), .A2(new_n587_), .A3(new_n592_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(new_n596_), .B1(KEYINPUT72), .B2(KEYINPUT13), .ZN(new_n597_));
  XNOR2_X1  g396(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n594_), .A2(new_n595_), .A3(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  XOR2_X1   g399(.A(new_n600_), .B(KEYINPUT73), .Z(new_n601_));
  AND3_X1   g400(.A1(new_n553_), .A2(new_n569_), .A3(new_n601_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n602_), .A2(new_n528_), .A3(new_n324_), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n603_), .B(KEYINPUT38), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n600_), .A2(new_n569_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n605_), .A2(new_n550_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  XOR2_X1   g406(.A(new_n499_), .B(KEYINPUT97), .Z(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT98), .B1(new_n408_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n379_), .A2(new_n401_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n405_), .A2(new_n407_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n613_), .A2(new_n614_), .A3(new_n608_), .ZN(new_n615_));
  AOI21_X1  g414(.A(new_n607_), .B1(new_n610_), .B2(new_n615_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n616_), .A2(new_n324_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n604_), .B1(new_n528_), .B2(new_n617_), .ZN(G1324gat));
  INV_X1    g417(.A(new_n280_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n602_), .A2(new_n529_), .A3(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT39), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n616_), .A2(new_n619_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n621_), .B1(new_n622_), .B2(G8gat), .ZN(new_n623_));
  AOI211_X1 g422(.A(KEYINPUT39), .B(new_n529_), .C1(new_n616_), .C2(new_n619_), .ZN(new_n624_));
  OAI21_X1  g423(.A(new_n620_), .B1(new_n623_), .B2(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n625_), .B(new_n627_), .ZN(G1325gat));
  INV_X1    g427(.A(G15gat), .ZN(new_n629_));
  AOI21_X1  g428(.A(new_n629_), .B1(new_n616_), .B2(new_n400_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT41), .ZN(new_n631_));
  OR2_X1    g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n631_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n602_), .A2(new_n629_), .A3(new_n400_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n632_), .A2(new_n633_), .A3(new_n634_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  NAND4_X1  g436(.A1(new_n632_), .A2(KEYINPUT100), .A3(new_n633_), .A4(new_n634_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n637_), .A2(new_n638_), .ZN(G1326gat));
  INV_X1    g438(.A(G22gat), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n640_), .B1(new_n616_), .B2(new_n378_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT42), .Z(new_n642_));
  NAND3_X1  g441(.A1(new_n602_), .A2(new_n640_), .A3(new_n378_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(G1327gat));
  INV_X1    g443(.A(G29gat), .ZN(new_n645_));
  INV_X1    g444(.A(new_n605_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n499_), .ZN(new_n647_));
  NOR2_X1   g446(.A1(new_n549_), .A2(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n613_), .A2(new_n646_), .A3(new_n648_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n649_), .B2(new_n325_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n646_), .A2(new_n550_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(new_n651_), .B(KEYINPUT101), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  NOR3_X1   g452(.A1(new_n408_), .A2(KEYINPUT43), .A3(new_n503_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT43), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n655_), .B1(new_n613_), .B2(new_n504_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n653_), .B1(new_n654_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n659_), .A2(G29gat), .A3(new_n324_), .ZN(new_n660_));
  OAI21_X1  g459(.A(KEYINPUT43), .B1(new_n408_), .B2(new_n503_), .ZN(new_n661_));
  NAND3_X1  g460(.A1(new_n613_), .A2(new_n655_), .A3(new_n504_), .ZN(new_n662_));
  AOI21_X1  g461(.A(new_n652_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n663_), .A2(KEYINPUT44), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  OAI21_X1  g464(.A(new_n650_), .B1(new_n660_), .B2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT102), .ZN(new_n667_));
  XNOR2_X1  g466(.A(new_n666_), .B(new_n667_), .ZN(G1328gat));
  NAND2_X1  g467(.A1(KEYINPUT104), .A2(KEYINPUT46), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT46), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(G36gat), .ZN(new_n673_));
  AOI21_X1  g472(.A(new_n280_), .B1(new_n657_), .B2(new_n658_), .ZN(new_n674_));
  AOI21_X1  g473(.A(new_n673_), .B1(new_n674_), .B2(new_n664_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT45), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n280_), .A2(G36gat), .ZN(new_n677_));
  INV_X1    g476(.A(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT103), .B1(new_n649_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n679_), .ZN(new_n680_));
  NOR3_X1   g479(.A1(new_n649_), .A2(KEYINPUT103), .A3(new_n678_), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n676_), .B1(new_n680_), .B2(new_n681_), .ZN(new_n682_));
  OR3_X1    g481(.A1(new_n649_), .A2(KEYINPUT103), .A3(new_n678_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(KEYINPUT45), .A3(new_n679_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n682_), .A2(new_n684_), .ZN(new_n685_));
  OAI211_X1 g484(.A(new_n669_), .B(new_n672_), .C1(new_n675_), .C2(new_n685_), .ZN(new_n686_));
  NOR3_X1   g485(.A1(new_n680_), .A2(new_n681_), .A3(new_n676_), .ZN(new_n687_));
  AOI21_X1  g486(.A(KEYINPUT45), .B1(new_n683_), .B2(new_n679_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n619_), .B1(new_n663_), .B2(KEYINPUT44), .ZN(new_n690_));
  OAI21_X1  g489(.A(G36gat), .B1(new_n665_), .B2(new_n690_), .ZN(new_n691_));
  NAND4_X1  g490(.A1(new_n689_), .A2(new_n691_), .A3(new_n670_), .A4(new_n671_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n686_), .A2(new_n692_), .ZN(G1329gat));
  INV_X1    g492(.A(G43gat), .ZN(new_n694_));
  OAI21_X1  g493(.A(new_n694_), .B1(new_n649_), .B2(new_n401_), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n659_), .A2(G43gat), .A3(new_n400_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n695_), .B1(new_n696_), .B2(new_n665_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g497(.A(new_n649_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G50gat), .B1(new_n699_), .B2(new_n378_), .ZN(new_n700_));
  AND3_X1   g499(.A1(new_n659_), .A2(G50gat), .A3(new_n378_), .ZN(new_n701_));
  AOI21_X1  g500(.A(new_n700_), .B1(new_n701_), .B2(new_n664_), .ZN(G1331gat));
  INV_X1    g501(.A(G57gat), .ZN(new_n703_));
  NOR2_X1   g502(.A1(new_n600_), .A2(new_n569_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n553_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n703_), .B1(new_n705_), .B2(new_n325_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT105), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n601_), .A2(new_n569_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(new_n549_), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n610_), .B2(new_n615_), .ZN(new_n710_));
  INV_X1    g509(.A(new_n710_), .ZN(new_n711_));
  NOR3_X1   g510(.A1(new_n711_), .A2(new_n703_), .A3(new_n325_), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n707_), .A2(new_n712_), .ZN(G1332gat));
  INV_X1    g512(.A(new_n705_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(new_n280_), .A2(G64gat), .ZN(new_n715_));
  XNOR2_X1  g514(.A(new_n715_), .B(KEYINPUT106), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n710_), .A2(new_n619_), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT48), .ZN(new_n719_));
  AND3_X1   g518(.A1(new_n718_), .A2(new_n719_), .A3(G64gat), .ZN(new_n720_));
  AOI21_X1  g519(.A(new_n719_), .B1(new_n718_), .B2(G64gat), .ZN(new_n721_));
  OAI21_X1  g520(.A(new_n717_), .B1(new_n720_), .B2(new_n721_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(KEYINPUT107), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT107), .ZN(new_n724_));
  OAI211_X1 g523(.A(new_n724_), .B(new_n717_), .C1(new_n720_), .C2(new_n721_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n723_), .A2(new_n725_), .ZN(G1333gat));
  OR3_X1    g525(.A1(new_n705_), .A2(G71gat), .A3(new_n401_), .ZN(new_n727_));
  OAI21_X1  g526(.A(G71gat), .B1(new_n711_), .B2(new_n401_), .ZN(new_n728_));
  XOR2_X1   g527(.A(KEYINPUT108), .B(KEYINPUT49), .Z(new_n729_));
  AND2_X1   g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  NOR2_X1   g529(.A1(new_n728_), .A2(new_n729_), .ZN(new_n731_));
  OAI21_X1  g530(.A(new_n727_), .B1(new_n730_), .B2(new_n731_), .ZN(G1334gat));
  AOI21_X1  g531(.A(new_n341_), .B1(new_n710_), .B2(new_n378_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(KEYINPUT109), .B(KEYINPUT50), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n733_), .B(new_n734_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n714_), .A2(new_n341_), .A3(new_n378_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1335gat));
  NAND3_X1  g536(.A1(new_n613_), .A2(new_n648_), .A3(new_n708_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(G85gat), .B1(new_n739_), .B2(new_n324_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n704_), .A2(new_n550_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n741_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n742_));
  NOR2_X1   g541(.A1(new_n325_), .A2(new_n317_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n740_), .B1(new_n742_), .B2(new_n743_), .ZN(G1336gat));
  AOI21_X1  g543(.A(G92gat), .B1(new_n739_), .B2(new_n619_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n280_), .A2(new_n266_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n742_), .B2(new_n746_), .ZN(G1337gat));
  AOI211_X1 g546(.A(new_n401_), .B(new_n738_), .C1(new_n416_), .C2(new_n411_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n742_), .A2(new_n400_), .ZN(new_n749_));
  AOI21_X1  g548(.A(new_n748_), .B1(new_n749_), .B2(G99gat), .ZN(new_n750_));
  XNOR2_X1  g549(.A(KEYINPUT110), .B(KEYINPUT51), .ZN(new_n751_));
  XOR2_X1   g550(.A(new_n750_), .B(new_n751_), .Z(G1338gat));
  NAND3_X1  g551(.A1(new_n739_), .A2(new_n352_), .A3(new_n378_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n742_), .A2(new_n378_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n754_), .B1(new_n755_), .B2(G106gat), .ZN(new_n756_));
  AOI211_X1 g555(.A(KEYINPUT52), .B(new_n352_), .C1(new_n742_), .C2(new_n378_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n753_), .B1(new_n756_), .B2(new_n757_), .ZN(new_n758_));
  XNOR2_X1  g557(.A(new_n758_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g558(.A(KEYINPUT56), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n574_), .B1(new_n452_), .B2(new_n526_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n452_), .A2(new_n526_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n575_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n762_), .B(new_n763_), .C1(new_n481_), .C2(new_n764_), .ZN(new_n765_));
  AOI21_X1  g564(.A(new_n761_), .B1(new_n765_), .B2(new_n583_), .ZN(new_n766_));
  NOR2_X1   g565(.A1(new_n765_), .A2(new_n583_), .ZN(new_n767_));
  NOR2_X1   g566(.A1(new_n766_), .A2(new_n767_), .ZN(new_n768_));
  NOR3_X1   g567(.A1(new_n765_), .A2(new_n761_), .A3(new_n583_), .ZN(new_n769_));
  OAI211_X1 g568(.A(new_n760_), .B(new_n593_), .C1(new_n768_), .C2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n770_), .A2(new_n595_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n584_), .B1(new_n576_), .B2(new_n581_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n585_), .B1(new_n772_), .B2(new_n761_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n769_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n773_), .A2(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n760_), .B1(new_n775_), .B2(new_n593_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n564_), .B1(new_n559_), .B2(new_n557_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n556_), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n777_), .B1(new_n778_), .B2(new_n557_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n565_), .A2(new_n779_), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n771_), .A2(new_n776_), .A3(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n504_), .B1(new_n781_), .B2(KEYINPUT58), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT112), .ZN(new_n783_));
  OAI21_X1  g582(.A(new_n593_), .B1(new_n768_), .B2(new_n769_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n784_), .A2(KEYINPUT56), .ZN(new_n785_));
  INV_X1    g584(.A(new_n780_), .ZN(new_n786_));
  NAND4_X1  g585(.A1(new_n785_), .A2(new_n595_), .A3(new_n786_), .A4(new_n770_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT58), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n503_), .B1(new_n787_), .B2(new_n788_), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT112), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n789_), .A2(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n781_), .A2(KEYINPUT58), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n783_), .A2(new_n791_), .A3(new_n792_), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n785_), .A2(new_n569_), .A3(new_n595_), .A4(new_n770_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n596_), .A2(new_n786_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT57), .B1(new_n796_), .B2(new_n647_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  AOI211_X1 g597(.A(new_n798_), .B(new_n499_), .C1(new_n794_), .C2(new_n795_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(new_n797_), .A2(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n549_), .B1(new_n793_), .B2(new_n800_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n569_), .B1(new_n597_), .B2(new_n599_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n802_), .A2(new_n549_), .A3(new_n503_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n803_), .A2(KEYINPUT111), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT111), .ZN(new_n805_));
  NAND4_X1  g604(.A1(new_n802_), .A2(new_n805_), .A3(new_n503_), .A4(new_n549_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n804_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n804_), .A2(KEYINPUT54), .A3(new_n806_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n809_), .A2(new_n810_), .ZN(new_n811_));
  OAI21_X1  g610(.A(KEYINPUT113), .B1(new_n801_), .B2(new_n811_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n796_), .A2(new_n647_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n813_), .A2(new_n798_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n796_), .A2(KEYINPUT57), .A3(new_n647_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n792_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n816_));
  AOI211_X1 g615(.A(KEYINPUT112), .B(new_n503_), .C1(new_n787_), .C2(new_n788_), .ZN(new_n817_));
  OAI211_X1 g616(.A(new_n814_), .B(new_n815_), .C1(new_n816_), .C2(new_n817_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(new_n550_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n820_));
  AND3_X1   g619(.A1(new_n804_), .A2(KEYINPUT54), .A3(new_n806_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT54), .B1(new_n804_), .B2(new_n806_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n819_), .A2(new_n820_), .A3(new_n823_), .ZN(new_n824_));
  NOR4_X1   g623(.A1(new_n378_), .A2(new_n619_), .A3(new_n325_), .A4(new_n401_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n812_), .A2(new_n824_), .A3(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(G113gat), .B1(new_n827_), .B2(new_n569_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(KEYINPUT59), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n829_), .A2(KEYINPUT114), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n826_), .A2(new_n831_), .A3(KEYINPUT59), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(KEYINPUT59), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n834_), .B(new_n825_), .C1(new_n801_), .C2(new_n811_), .ZN(new_n835_));
  AND2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  AND2_X1   g635(.A1(new_n569_), .A2(G113gat), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n828_), .B1(new_n836_), .B2(new_n837_), .ZN(G1340gat));
  INV_X1    g637(.A(new_n601_), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n826_), .A2(new_n831_), .A3(KEYINPUT59), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n831_), .B1(new_n826_), .B2(KEYINPUT59), .ZN(new_n841_));
  OAI211_X1 g640(.A(new_n839_), .B(new_n835_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT115), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n833_), .A2(KEYINPUT115), .A3(new_n839_), .A4(new_n835_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n844_), .A2(new_n845_), .A3(G120gat), .ZN(new_n846_));
  INV_X1    g645(.A(G120gat), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n600_), .B2(KEYINPUT60), .ZN(new_n848_));
  OAI211_X1 g647(.A(new_n827_), .B(new_n848_), .C1(KEYINPUT60), .C2(new_n847_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n846_), .A2(new_n849_), .ZN(G1341gat));
  AOI21_X1  g649(.A(G127gat), .B1(new_n827_), .B2(new_n549_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n549_), .A2(G127gat), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT116), .ZN(new_n853_));
  AOI21_X1  g652(.A(new_n851_), .B1(new_n836_), .B2(new_n853_), .ZN(G1342gat));
  INV_X1    g653(.A(G134gat), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n503_), .A2(new_n855_), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n835_), .B(new_n856_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n855_), .B1(new_n826_), .B2(new_n608_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n857_), .A2(KEYINPUT117), .A3(new_n858_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n861_), .A2(new_n862_), .ZN(G1343gat));
  NOR4_X1   g662(.A1(new_n406_), .A2(new_n619_), .A3(new_n325_), .A4(new_n400_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n812_), .A2(new_n824_), .A3(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n865_), .A2(new_n866_), .ZN(new_n867_));
  NAND4_X1  g666(.A1(new_n812_), .A2(new_n824_), .A3(KEYINPUT118), .A4(new_n864_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n867_), .A2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n869_), .A2(new_n569_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(G141gat), .ZN(G1344gat));
  XNOR2_X1  g670(.A(KEYINPUT119), .B(G148gat), .ZN(new_n872_));
  INV_X1    g671(.A(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT120), .ZN(new_n874_));
  NAND3_X1  g673(.A1(new_n869_), .A2(new_n874_), .A3(new_n839_), .ZN(new_n875_));
  INV_X1    g674(.A(new_n875_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n874_), .B1(new_n869_), .B2(new_n839_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n873_), .B1(new_n876_), .B2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n877_), .ZN(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(new_n875_), .A3(new_n872_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n880_), .ZN(G1345gat));
  XNOR2_X1  g680(.A(KEYINPUT61), .B(G155gat), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n869_), .A2(new_n549_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(KEYINPUT121), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n869_), .A2(new_n885_), .A3(new_n549_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n882_), .B1(new_n884_), .B2(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n885_), .B1(new_n869_), .B2(new_n549_), .ZN(new_n888_));
  AOI211_X1 g687(.A(KEYINPUT121), .B(new_n550_), .C1(new_n867_), .C2(new_n868_), .ZN(new_n889_));
  INV_X1    g688(.A(new_n882_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n888_), .A2(new_n889_), .A3(new_n890_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n887_), .A2(new_n891_), .ZN(G1346gat));
  AOI21_X1  g691(.A(G162gat), .B1(new_n869_), .B2(new_n609_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n504_), .A2(G162gat), .ZN(new_n894_));
  AOI21_X1  g693(.A(new_n893_), .B1(new_n869_), .B2(new_n894_), .ZN(G1347gat));
  INV_X1    g694(.A(KEYINPUT62), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n896_), .A2(KEYINPUT123), .ZN(new_n897_));
  AOI21_X1  g696(.A(new_n378_), .B1(new_n819_), .B2(new_n823_), .ZN(new_n898_));
  NOR3_X1   g697(.A1(new_n280_), .A2(new_n324_), .A3(new_n401_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n569_), .ZN(new_n900_));
  XOR2_X1   g699(.A(new_n900_), .B(KEYINPUT122), .Z(new_n901_));
  NAND2_X1  g700(.A1(new_n898_), .A2(new_n901_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n897_), .B1(new_n902_), .B2(G169gat), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n896_), .A2(KEYINPUT123), .ZN(new_n904_));
  INV_X1    g703(.A(new_n904_), .ZN(new_n905_));
  OR2_X1    g704(.A1(new_n903_), .A2(new_n905_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n903_), .A2(new_n905_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n898_), .A2(new_n899_), .ZN(new_n908_));
  INV_X1    g707(.A(new_n908_), .ZN(new_n909_));
  NAND3_X1  g708(.A1(new_n909_), .A2(new_n202_), .A3(new_n569_), .ZN(new_n910_));
  NAND3_X1  g709(.A1(new_n906_), .A2(new_n907_), .A3(new_n910_), .ZN(new_n911_));
  XNOR2_X1  g710(.A(new_n911_), .B(KEYINPUT124), .ZN(G1348gat));
  OAI21_X1  g711(.A(new_n203_), .B1(new_n908_), .B2(new_n600_), .ZN(new_n913_));
  XOR2_X1   g712(.A(new_n913_), .B(KEYINPUT125), .Z(new_n914_));
  AND2_X1   g713(.A1(new_n812_), .A2(new_n824_), .ZN(new_n915_));
  AND2_X1   g714(.A1(new_n915_), .A2(new_n406_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n899_), .ZN(new_n917_));
  NOR3_X1   g716(.A1(new_n917_), .A2(new_n601_), .A3(new_n203_), .ZN(new_n918_));
  AOI21_X1  g717(.A(new_n914_), .B1(new_n916_), .B2(new_n918_), .ZN(G1349gat));
  NOR2_X1   g718(.A1(new_n917_), .A2(new_n550_), .ZN(new_n920_));
  AOI21_X1  g719(.A(G183gat), .B1(new_n916_), .B2(new_n920_), .ZN(new_n921_));
  NOR2_X1   g720(.A1(new_n550_), .A2(new_n215_), .ZN(new_n922_));
  INV_X1    g721(.A(new_n922_), .ZN(new_n923_));
  OR3_X1    g722(.A1(new_n908_), .A2(KEYINPUT126), .A3(new_n923_), .ZN(new_n924_));
  OAI21_X1  g723(.A(KEYINPUT126), .B1(new_n908_), .B2(new_n923_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT127), .ZN(new_n927_));
  OR3_X1    g726(.A1(new_n921_), .A2(new_n926_), .A3(new_n927_), .ZN(new_n928_));
  OAI21_X1  g727(.A(new_n927_), .B1(new_n921_), .B2(new_n926_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n928_), .A2(new_n929_), .ZN(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n908_), .B2(new_n503_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n609_), .A2(new_n216_), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n908_), .B2(new_n932_), .ZN(G1351gat));
  NOR4_X1   g732(.A1(new_n406_), .A2(new_n324_), .A3(new_n280_), .A4(new_n400_), .ZN(new_n934_));
  AND2_X1   g733(.A1(new_n915_), .A2(new_n934_), .ZN(new_n935_));
  NAND2_X1  g734(.A1(new_n935_), .A2(new_n569_), .ZN(new_n936_));
  XNOR2_X1  g735(.A(new_n936_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g736(.A1(new_n935_), .A2(new_n839_), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n938_), .B(G204gat), .ZN(G1353gat));
  AND2_X1   g738(.A1(new_n935_), .A2(new_n549_), .ZN(new_n940_));
  NOR3_X1   g739(.A1(new_n940_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941_));
  XOR2_X1   g740(.A(KEYINPUT63), .B(G211gat), .Z(new_n942_));
  AOI21_X1  g741(.A(new_n941_), .B1(new_n940_), .B2(new_n942_), .ZN(G1354gat));
  AOI21_X1  g742(.A(G218gat), .B1(new_n935_), .B2(new_n609_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n504_), .A2(G218gat), .ZN(new_n945_));
  AOI21_X1  g744(.A(new_n944_), .B1(new_n935_), .B2(new_n945_), .ZN(G1355gat));
endmodule


