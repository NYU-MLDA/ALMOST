//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 0 0 0 1 1 0 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n600_, new_n601_, new_n602_, new_n603_, new_n604_, new_n605_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n650_, new_n651_,
    new_n652_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n672_,
    new_n673_, new_n674_, new_n675_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n693_, new_n694_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n811_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n821_, new_n822_,
    new_n823_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n858_,
    new_n859_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n877_, new_n878_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT10), .B(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n204_));
  XNOR2_X1  g003(.A(new_n203_), .B(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(G106gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT66), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT6), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n209_), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NOR2_X1   g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  OAI21_X1  g011(.A(new_n208_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n209_), .A2(G99gat), .A3(G106gat), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT66), .ZN(new_n216_));
  AND2_X1   g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  NOR2_X1   g017(.A1(new_n218_), .A2(KEYINPUT9), .ZN(new_n219_));
  INV_X1    g018(.A(new_n218_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(G85gat), .A2(G92gat), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n219_), .B1(new_n222_), .B2(KEYINPUT9), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n207_), .A2(new_n217_), .A3(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT69), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n226_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT69), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT7), .ZN(new_n229_));
  INV_X1    g028(.A(G99gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(new_n206_), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n232_));
  AND2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n227_), .A2(new_n228_), .A3(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n235_));
  OAI21_X1  g034(.A(new_n235_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n236_));
  INV_X1    g035(.A(G85gat), .ZN(new_n237_));
  INV_X1    g036(.A(G92gat), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n239_), .A2(KEYINPUT67), .A3(new_n218_), .ZN(new_n240_));
  AND2_X1   g039(.A1(new_n236_), .A2(new_n240_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n234_), .A2(KEYINPUT70), .A3(new_n241_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n242_), .A2(KEYINPUT8), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT70), .B1(new_n234_), .B2(new_n241_), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NAND3_X1  g044(.A1(new_n213_), .A2(new_n216_), .A3(new_n233_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT8), .ZN(new_n247_));
  AND3_X1   g046(.A1(new_n236_), .A2(new_n240_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n246_), .A2(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT68), .ZN(new_n250_));
  INV_X1    g049(.A(KEYINPUT68), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n246_), .A2(new_n248_), .A3(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n225_), .B1(new_n245_), .B2(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(G64gat), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n255_), .A2(G57gat), .ZN(new_n256_));
  INV_X1    g055(.A(G57gat), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(G64gat), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n258_), .A3(KEYINPUT11), .ZN(new_n259_));
  INV_X1    g058(.A(G71gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n260_), .A2(KEYINPUT71), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT71), .ZN(new_n262_));
  NAND2_X1  g061(.A1(new_n262_), .A2(G71gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n261_), .A2(new_n263_), .ZN(new_n264_));
  NOR2_X1   g063(.A1(new_n264_), .A2(G78gat), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT71), .B(G71gat), .ZN(new_n266_));
  INV_X1    g065(.A(G78gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n259_), .B1(new_n265_), .B2(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n264_), .A2(G78gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n266_), .A2(new_n267_), .ZN(new_n271_));
  INV_X1    g070(.A(new_n259_), .ZN(new_n272_));
  AOI21_X1  g071(.A(KEYINPUT11), .B1(new_n256_), .B2(new_n258_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n270_), .B(new_n271_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n269_), .A2(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n254_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n277_));
  AND3_X1   g076(.A1(new_n214_), .A2(new_n215_), .A3(KEYINPUT69), .ZN(new_n278_));
  AOI21_X1  g077(.A(KEYINPUT69), .B1(new_n214_), .B2(new_n215_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n231_), .A2(new_n232_), .ZN(new_n280_));
  NOR3_X1   g079(.A1(new_n278_), .A2(new_n279_), .A3(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n236_), .A2(new_n240_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n277_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND3_X1  g082(.A1(new_n283_), .A2(KEYINPUT8), .A3(new_n242_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n246_), .A2(new_n248_), .A3(new_n251_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n251_), .B1(new_n246_), .B2(new_n248_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  AOI21_X1  g086(.A(new_n224_), .B1(new_n284_), .B2(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n275_), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n288_), .A2(new_n289_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n276_), .A2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(G230gat), .A2(G233gat), .ZN(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT64), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n291_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT12), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n295_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n296_));
  AOI21_X1  g095(.A(new_n293_), .B1(new_n288_), .B2(new_n289_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n298_));
  AND3_X1   g097(.A1(new_n269_), .A2(new_n274_), .A3(new_n298_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n298_), .B1(new_n269_), .B2(new_n274_), .ZN(new_n300_));
  OAI21_X1  g099(.A(KEYINPUT12), .B1(new_n299_), .B2(new_n300_), .ZN(new_n301_));
  INV_X1    g100(.A(new_n301_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n254_), .A2(new_n302_), .ZN(new_n303_));
  NAND3_X1  g102(.A1(new_n296_), .A2(new_n297_), .A3(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n294_), .A2(new_n304_), .ZN(new_n305_));
  XOR2_X1   g104(.A(G176gat), .B(G204gat), .Z(new_n306_));
  XNOR2_X1  g105(.A(new_n306_), .B(KEYINPUT74), .ZN(new_n307_));
  XOR2_X1   g106(.A(G120gat), .B(G148gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n309_), .B(new_n310_), .Z(new_n311_));
  NAND2_X1  g110(.A1(new_n305_), .A2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n311_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n294_), .A2(new_n304_), .A3(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n312_), .A2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT13), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n315_), .A2(new_n316_), .ZN(new_n317_));
  NAND3_X1  g116(.A1(new_n312_), .A2(KEYINPUT13), .A3(new_n314_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n317_), .A2(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G229gat), .A2(G233gat), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  XNOR2_X1  g121(.A(KEYINPUT79), .B(G8gat), .ZN(new_n323_));
  OAI21_X1  g122(.A(KEYINPUT14), .B1(new_n323_), .B2(new_n202_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G15gat), .B(G22gat), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  INV_X1    g125(.A(KEYINPUT80), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G1gat), .B(G8gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n326_), .B(KEYINPUT80), .ZN(new_n331_));
  INV_X1    g130(.A(new_n329_), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n331_), .A2(new_n332_), .ZN(new_n333_));
  XNOR2_X1  g132(.A(G29gat), .B(G36gat), .ZN(new_n334_));
  XNOR2_X1  g133(.A(G43gat), .B(G50gat), .ZN(new_n335_));
  XNOR2_X1  g134(.A(new_n334_), .B(new_n335_), .ZN(new_n336_));
  NAND3_X1  g135(.A1(new_n330_), .A2(new_n333_), .A3(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n336_), .B1(new_n330_), .B2(new_n333_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n322_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n330_), .A2(new_n333_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(KEYINPUT75), .B(KEYINPUT15), .ZN(new_n342_));
  XNOR2_X1  g141(.A(new_n336_), .B(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n341_), .A2(new_n343_), .ZN(new_n344_));
  NAND3_X1  g143(.A1(new_n344_), .A2(new_n337_), .A3(new_n321_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G113gat), .B(G141gat), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT82), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G169gat), .B(G197gat), .ZN(new_n348_));
  XOR2_X1   g147(.A(new_n347_), .B(new_n348_), .Z(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND3_X1  g149(.A1(new_n340_), .A2(new_n345_), .A3(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT84), .ZN(new_n352_));
  OR2_X1    g151(.A1(new_n351_), .A2(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n352_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n353_), .A2(new_n354_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n340_), .A2(new_n345_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n349_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT83), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT83), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n356_), .A2(new_n359_), .A3(new_n349_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n358_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n355_), .A2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n320_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT102), .ZN(new_n364_));
  AND2_X1   g163(.A1(G231gat), .A2(G233gat), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n341_), .B(new_n365_), .ZN(new_n366_));
  XOR2_X1   g165(.A(new_n366_), .B(KEYINPUT81), .Z(new_n367_));
  INV_X1    g166(.A(new_n299_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n300_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n367_), .A2(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT17), .ZN(new_n372_));
  XOR2_X1   g171(.A(G127gat), .B(G155gat), .Z(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(KEYINPUT16), .ZN(new_n374_));
  XNOR2_X1  g173(.A(G183gat), .B(G211gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  NOR3_X1   g175(.A1(new_n371_), .A2(new_n372_), .A3(new_n376_), .ZN(new_n377_));
  OAI21_X1  g176(.A(new_n377_), .B1(new_n370_), .B2(new_n367_), .ZN(new_n378_));
  OR2_X1    g177(.A1(new_n366_), .A2(new_n289_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n366_), .A2(new_n289_), .ZN(new_n380_));
  XNOR2_X1  g179(.A(new_n376_), .B(KEYINPUT17), .ZN(new_n381_));
  NAND3_X1  g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n378_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  AND3_X1   g183(.A1(new_n364_), .A2(KEYINPUT103), .A3(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT103), .B1(new_n364_), .B2(new_n384_), .ZN(new_n386_));
  XOR2_X1   g185(.A(KEYINPUT98), .B(KEYINPUT0), .Z(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(KEYINPUT99), .ZN(new_n388_));
  XOR2_X1   g187(.A(G1gat), .B(G29gat), .Z(new_n389_));
  XNOR2_X1  g188(.A(new_n388_), .B(new_n389_), .ZN(new_n390_));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391_));
  XOR2_X1   g190(.A(new_n390_), .B(new_n391_), .Z(new_n392_));
  INV_X1    g191(.A(KEYINPUT4), .ZN(new_n393_));
  XOR2_X1   g192(.A(G113gat), .B(G120gat), .Z(new_n394_));
  XNOR2_X1  g193(.A(new_n394_), .B(KEYINPUT89), .ZN(new_n395_));
  XOR2_X1   g194(.A(G127gat), .B(G134gat), .Z(new_n396_));
  XOR2_X1   g195(.A(new_n395_), .B(new_n396_), .Z(new_n397_));
  NAND2_X1  g196(.A1(new_n397_), .A2(KEYINPUT90), .ZN(new_n398_));
  OR3_X1    g197(.A1(new_n395_), .A2(KEYINPUT90), .A3(new_n396_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n398_), .A2(new_n399_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G155gat), .A2(G162gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NOR2_X1   g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403_));
  NOR2_X1   g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G141gat), .A2(G148gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n405_), .B(KEYINPUT92), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT2), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(new_n408_), .B(KEYINPUT93), .ZN(new_n409_));
  NOR2_X1   g208(.A1(G141gat), .A2(G148gat), .ZN(new_n410_));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  OAI21_X1  g211(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n412_), .B(new_n413_), .C1(new_n407_), .C2(new_n405_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n404_), .B1(new_n409_), .B2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT1), .ZN(new_n416_));
  OAI221_X1 g215(.A(new_n406_), .B1(new_n416_), .B2(new_n401_), .C1(G141gat), .C2(G148gat), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n417_), .B1(new_n416_), .B2(new_n404_), .ZN(new_n418_));
  INV_X1    g217(.A(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n415_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n400_), .A2(new_n420_), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n420_), .A2(new_n397_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n393_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT4), .B1(new_n400_), .B2(new_n420_), .ZN(new_n424_));
  NOR2_X1   g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426_));
  INV_X1    g225(.A(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n425_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  AOI21_X1  g228(.A(new_n427_), .B1(new_n421_), .B2(new_n422_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n392_), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT101), .ZN(new_n432_));
  INV_X1    g231(.A(new_n392_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n430_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n428_), .A2(new_n433_), .A3(new_n434_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n431_), .A2(new_n432_), .A3(new_n435_), .ZN(new_n436_));
  NAND4_X1  g235(.A1(new_n428_), .A2(KEYINPUT101), .A3(new_n433_), .A4(new_n434_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n436_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT27), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G211gat), .B(G218gat), .ZN(new_n440_));
  XOR2_X1   g239(.A(KEYINPUT95), .B(G204gat), .Z(new_n441_));
  NOR2_X1   g240(.A1(new_n441_), .A2(G197gat), .ZN(new_n442_));
  INV_X1    g241(.A(G197gat), .ZN(new_n443_));
  INV_X1    g242(.A(G204gat), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT21), .B1(new_n443_), .B2(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(G197gat), .A2(G204gat), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n446_), .B1(new_n441_), .B2(G197gat), .ZN(new_n447_));
  OAI221_X1 g246(.A(new_n440_), .B1(new_n442_), .B2(new_n445_), .C1(KEYINPUT21), .C2(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(new_n440_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(KEYINPUT21), .A3(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G183gat), .A2(G190gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(KEYINPUT23), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT24), .ZN(new_n455_));
  INV_X1    g254(.A(G169gat), .ZN(new_n456_));
  INV_X1    g255(.A(G176gat), .ZN(new_n457_));
  NAND3_X1  g256(.A1(new_n455_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n458_));
  AND2_X1   g257(.A1(new_n454_), .A2(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT25), .B(G183gat), .ZN(new_n460_));
  INV_X1    g259(.A(G190gat), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n461_), .A2(KEYINPUT26), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(KEYINPUT26), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n460_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n464_));
  OAI21_X1  g263(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G169gat), .A2(G176gat), .ZN(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  OAI211_X1 g266(.A(new_n459_), .B(new_n464_), .C1(new_n465_), .C2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n466_), .B(KEYINPUT87), .ZN(new_n469_));
  INV_X1    g268(.A(G183gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n470_), .A2(new_n461_), .ZN(new_n471_));
  AOI21_X1  g270(.A(new_n469_), .B1(new_n454_), .B2(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(KEYINPUT22), .B(G169gat), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n473_), .A2(new_n457_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  AND2_X1   g274(.A1(new_n468_), .A2(new_n475_), .ZN(new_n476_));
  OR3_X1    g275(.A1(new_n452_), .A2(new_n476_), .A3(KEYINPUT97), .ZN(new_n477_));
  OAI21_X1  g276(.A(KEYINPUT97), .B1(new_n452_), .B2(new_n476_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(new_n474_), .B(KEYINPUT88), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n472_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT86), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n463_), .A2(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n461_), .A2(KEYINPUT86), .A3(KEYINPUT26), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n460_), .A2(new_n482_), .A3(new_n462_), .A4(new_n483_), .ZN(new_n484_));
  OAI211_X1 g283(.A(new_n459_), .B(new_n484_), .C1(new_n465_), .C2(new_n469_), .ZN(new_n485_));
  AND2_X1   g284(.A1(new_n480_), .A2(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n452_), .A2(new_n486_), .ZN(new_n487_));
  NAND4_X1  g286(.A1(new_n477_), .A2(KEYINPUT20), .A3(new_n478_), .A4(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(G226gat), .A2(G233gat), .ZN(new_n489_));
  XNOR2_X1  g288(.A(new_n489_), .B(KEYINPUT19), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G8gat), .B(G36gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT18), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G64gat), .B(G92gat), .ZN(new_n494_));
  XOR2_X1   g293(.A(new_n493_), .B(new_n494_), .Z(new_n495_));
  NAND2_X1  g294(.A1(new_n452_), .A2(new_n476_), .ZN(new_n496_));
  OAI211_X1 g295(.A(new_n496_), .B(KEYINPUT20), .C1(new_n452_), .C2(new_n486_), .ZN(new_n497_));
  OR2_X1    g296(.A1(new_n497_), .A2(new_n490_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n491_), .A2(new_n495_), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n495_), .B1(new_n491_), .B2(new_n498_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n439_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  NOR2_X1   g300(.A1(new_n499_), .A2(new_n439_), .ZN(new_n502_));
  NOR2_X1   g301(.A1(new_n488_), .A2(new_n490_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n503_), .B1(new_n490_), .B2(new_n497_), .ZN(new_n504_));
  OAI21_X1  g303(.A(new_n502_), .B1(new_n495_), .B2(new_n504_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n438_), .A2(new_n501_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT29), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n415_), .A2(new_n508_), .A3(new_n419_), .ZN(new_n509_));
  XOR2_X1   g308(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n510_));
  XNOR2_X1  g309(.A(new_n509_), .B(new_n510_), .ZN(new_n511_));
  XOR2_X1   g310(.A(G22gat), .B(G50gat), .Z(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  OR2_X1    g312(.A1(new_n513_), .A2(KEYINPUT96), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(KEYINPUT96), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n452_), .B1(new_n420_), .B2(KEYINPUT29), .ZN(new_n516_));
  NAND2_X1  g315(.A1(G228gat), .A2(G233gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(new_n267_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(G106gat), .ZN(new_n519_));
  XOR2_X1   g318(.A(new_n516_), .B(new_n519_), .Z(new_n520_));
  NAND3_X1  g319(.A1(new_n514_), .A2(new_n515_), .A3(new_n520_), .ZN(new_n521_));
  OR2_X1    g320(.A1(new_n515_), .A2(new_n520_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  XOR2_X1   g322(.A(new_n400_), .B(KEYINPUT31), .Z(new_n524_));
  XNOR2_X1  g323(.A(G71gat), .B(G99gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(G43gat), .ZN(new_n526_));
  XNOR2_X1  g325(.A(new_n526_), .B(KEYINPUT30), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G227gat), .A2(G233gat), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n528_), .B(G15gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(new_n527_), .B(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(KEYINPUT91), .B1(new_n530_), .B2(new_n486_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n531_), .B1(new_n486_), .B2(new_n530_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n524_), .B(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  NOR2_X1   g333(.A1(new_n523_), .A2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n533_), .B1(new_n521_), .B2(new_n522_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n495_), .A2(KEYINPUT32), .ZN(new_n540_));
  OR2_X1    g339(.A1(new_n504_), .A2(new_n540_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n491_), .A2(new_n498_), .A3(new_n540_), .ZN(new_n542_));
  NAND4_X1  g341(.A1(new_n436_), .A2(new_n437_), .A3(new_n541_), .A4(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(KEYINPUT33), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n431_), .A2(KEYINPUT100), .A3(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n499_), .A2(new_n500_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(KEYINPUT100), .ZN(new_n547_));
  OAI211_X1 g346(.A(new_n392_), .B(new_n547_), .C1(new_n429_), .C2(new_n430_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n421_), .A2(new_n422_), .A3(new_n427_), .ZN(new_n549_));
  OAI211_X1 g348(.A(new_n549_), .B(new_n433_), .C1(new_n425_), .C2(new_n427_), .ZN(new_n550_));
  NAND4_X1  g349(.A1(new_n545_), .A2(new_n546_), .A3(new_n548_), .A4(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n543_), .A2(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n523_), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n553_), .A2(new_n534_), .ZN(new_n554_));
  AOI22_X1  g353(.A1(new_n507_), .A2(new_n539_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n254_), .A2(new_n343_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n288_), .A2(new_n336_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(G232gat), .A2(G233gat), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT34), .ZN(new_n559_));
  OAI211_X1 g358(.A(new_n556_), .B(new_n557_), .C1(KEYINPUT35), .C2(new_n559_), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n559_), .A2(KEYINPUT35), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT36), .ZN(new_n563_));
  XOR2_X1   g362(.A(G134gat), .B(G162gat), .Z(new_n564_));
  XNOR2_X1  g363(.A(new_n564_), .B(KEYINPUT78), .ZN(new_n565_));
  XOR2_X1   g364(.A(G190gat), .B(G218gat), .Z(new_n566_));
  XOR2_X1   g365(.A(new_n565_), .B(new_n566_), .Z(new_n567_));
  XNOR2_X1  g366(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n567_), .B(new_n568_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n562_), .A2(new_n563_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n569_), .B(new_n563_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n562_), .A2(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(new_n571_), .A2(new_n573_), .ZN(new_n574_));
  NOR4_X1   g373(.A1(new_n385_), .A2(new_n386_), .A3(new_n555_), .A4(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n438_), .ZN(new_n576_));
  AOI21_X1  g375(.A(new_n202_), .B1(new_n575_), .B2(new_n576_), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n577_), .B(KEYINPUT104), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n362_), .B(KEYINPUT85), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n555_), .A2(new_n579_), .ZN(new_n580_));
  OAI21_X1  g379(.A(KEYINPUT37), .B1(new_n571_), .B2(new_n573_), .ZN(new_n581_));
  INV_X1    g380(.A(KEYINPUT37), .ZN(new_n582_));
  OAI211_X1 g381(.A(new_n570_), .B(new_n582_), .C1(new_n562_), .C2(new_n572_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n581_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n584_), .ZN(new_n585_));
  NOR3_X1   g384(.A1(new_n383_), .A2(new_n585_), .A3(new_n319_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n580_), .A2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n588_), .A2(new_n202_), .A3(new_n576_), .ZN(new_n589_));
  XNOR2_X1  g388(.A(new_n589_), .B(KEYINPUT38), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n578_), .A2(new_n590_), .ZN(G1324gat));
  NAND2_X1  g390(.A1(new_n505_), .A2(new_n501_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n588_), .A2(new_n323_), .A3(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n575_), .A2(new_n592_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT39), .ZN(new_n595_));
  AND3_X1   g394(.A1(new_n594_), .A2(new_n595_), .A3(G8gat), .ZN(new_n596_));
  AOI21_X1  g395(.A(new_n595_), .B1(new_n594_), .B2(G8gat), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n593_), .B1(new_n596_), .B2(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT40), .Z(G1325gat));
  NAND2_X1  g398(.A1(new_n575_), .A2(new_n534_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n600_), .A2(G15gat), .ZN(new_n601_));
  OR2_X1    g400(.A1(new_n601_), .A2(KEYINPUT41), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(KEYINPUT41), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n587_), .A2(G15gat), .A3(new_n533_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT105), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n602_), .A2(new_n603_), .A3(new_n605_), .ZN(G1326gat));
  INV_X1    g405(.A(G22gat), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n588_), .A2(new_n607_), .A3(new_n553_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n607_), .B1(new_n575_), .B2(new_n553_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT42), .ZN(new_n610_));
  AND2_X1   g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n609_), .A2(new_n610_), .ZN(new_n612_));
  OAI21_X1  g411(.A(new_n608_), .B1(new_n611_), .B2(new_n612_), .ZN(new_n613_));
  XOR2_X1   g412(.A(new_n613_), .B(KEYINPUT106), .Z(G1327gat));
  INV_X1    g413(.A(new_n574_), .ZN(new_n615_));
  NOR3_X1   g414(.A1(new_n384_), .A2(new_n319_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n580_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n438_), .A2(G29gat), .ZN(new_n619_));
  XOR2_X1   g418(.A(new_n619_), .B(KEYINPUT108), .Z(new_n620_));
  NAND2_X1  g419(.A1(new_n618_), .A2(new_n620_), .ZN(new_n621_));
  AOI211_X1 g420(.A(new_n553_), .B(new_n534_), .C1(new_n543_), .C2(new_n551_), .ZN(new_n622_));
  AOI21_X1  g421(.A(new_n506_), .B1(new_n536_), .B2(new_n538_), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n585_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT43), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n384_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  OAI211_X1 g425(.A(KEYINPUT43), .B(new_n585_), .C1(new_n622_), .C2(new_n623_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n626_), .A2(KEYINPUT44), .A3(new_n364_), .A4(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(new_n625_), .B1(new_n555_), .B2(new_n584_), .ZN(new_n629_));
  NAND4_X1  g428(.A1(new_n629_), .A2(new_n627_), .A3(new_n364_), .A4(new_n383_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT44), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n630_), .A2(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n628_), .A2(new_n632_), .A3(new_n576_), .ZN(new_n633_));
  AND3_X1   g432(.A1(new_n633_), .A2(KEYINPUT107), .A3(G29gat), .ZN(new_n634_));
  AOI21_X1  g433(.A(KEYINPUT107), .B1(new_n633_), .B2(G29gat), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n621_), .B1(new_n634_), .B2(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT109), .ZN(new_n637_));
  INV_X1    g436(.A(KEYINPUT109), .ZN(new_n638_));
  OAI211_X1 g437(.A(new_n638_), .B(new_n621_), .C1(new_n634_), .C2(new_n635_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(G1328gat));
  XNOR2_X1  g439(.A(new_n592_), .B(KEYINPUT110), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NOR3_X1   g441(.A1(new_n617_), .A2(G36gat), .A3(new_n642_), .ZN(new_n643_));
  XOR2_X1   g442(.A(new_n643_), .B(KEYINPUT45), .Z(new_n644_));
  NAND3_X1  g443(.A1(new_n628_), .A2(new_n632_), .A3(new_n592_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(G36gat), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT46), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(G1329gat));
  NAND4_X1  g448(.A1(new_n628_), .A2(new_n632_), .A3(G43gat), .A4(new_n534_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n617_), .A2(new_n533_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n650_), .B1(G43gat), .B2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT47), .ZN(G1330gat));
  AND4_X1   g452(.A1(G50gat), .A2(new_n628_), .A3(new_n632_), .A4(new_n553_), .ZN(new_n654_));
  AOI21_X1  g453(.A(G50gat), .B1(new_n618_), .B2(new_n553_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1331gat));
  NAND3_X1  g455(.A1(new_n384_), .A2(new_n579_), .A3(new_n319_), .ZN(new_n657_));
  OR3_X1    g456(.A1(new_n555_), .A2(new_n574_), .A3(new_n657_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n658_), .A2(new_n257_), .A3(new_n438_), .ZN(new_n659_));
  XNOR2_X1  g458(.A(new_n659_), .B(KEYINPUT112), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n320_), .A2(new_n362_), .ZN(new_n661_));
  INV_X1    g460(.A(new_n661_), .ZN(new_n662_));
  NOR2_X1   g461(.A1(new_n555_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n383_), .A2(new_n585_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(G57gat), .B1(new_n666_), .B2(new_n576_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT111), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n667_), .A2(new_n668_), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n667_), .A2(new_n668_), .ZN(new_n670_));
  NOR3_X1   g469(.A1(new_n660_), .A2(new_n669_), .A3(new_n670_), .ZN(G1332gat));
  OAI21_X1  g470(.A(G64gat), .B1(new_n658_), .B2(new_n642_), .ZN(new_n672_));
  XOR2_X1   g471(.A(KEYINPUT113), .B(KEYINPUT48), .Z(new_n673_));
  XNOR2_X1  g472(.A(new_n672_), .B(new_n673_), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n666_), .A2(new_n255_), .A3(new_n641_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n674_), .A2(new_n675_), .ZN(G1333gat));
  OAI21_X1  g475(.A(G71gat), .B1(new_n658_), .B2(new_n533_), .ZN(new_n677_));
  XNOR2_X1  g476(.A(new_n677_), .B(KEYINPUT49), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n666_), .A2(new_n260_), .A3(new_n534_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  XOR2_X1   g479(.A(new_n680_), .B(KEYINPUT114), .Z(G1334gat));
  OAI21_X1  g480(.A(G78gat), .B1(new_n658_), .B2(new_n523_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT50), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n553_), .A2(new_n267_), .ZN(new_n684_));
  XNOR2_X1  g483(.A(new_n684_), .B(KEYINPUT115), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n683_), .B1(new_n665_), .B2(new_n685_), .ZN(G1335gat));
  NAND3_X1  g485(.A1(new_n626_), .A2(new_n627_), .A3(new_n661_), .ZN(new_n687_));
  OAI21_X1  g486(.A(G85gat), .B1(new_n687_), .B2(new_n438_), .ZN(new_n688_));
  NAND3_X1  g487(.A1(new_n663_), .A2(new_n383_), .A3(new_n574_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n690_), .A2(new_n237_), .A3(new_n576_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n688_), .A2(new_n691_), .ZN(G1336gat));
  OAI21_X1  g491(.A(G92gat), .B1(new_n687_), .B2(new_n642_), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n690_), .A2(new_n238_), .A3(new_n592_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n693_), .A2(new_n694_), .ZN(G1337gat));
  NAND3_X1  g494(.A1(new_n690_), .A2(new_n205_), .A3(new_n534_), .ZN(new_n696_));
  XNOR2_X1  g495(.A(new_n696_), .B(KEYINPUT116), .ZN(new_n697_));
  OAI21_X1  g496(.A(G99gat), .B1(new_n687_), .B2(new_n533_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n697_), .A2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g499(.A1(new_n690_), .A2(new_n206_), .A3(new_n553_), .ZN(new_n701_));
  NAND4_X1  g500(.A1(new_n626_), .A2(new_n553_), .A3(new_n627_), .A4(new_n661_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n703_));
  AND3_X1   g502(.A1(new_n702_), .A2(G106gat), .A3(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n703_), .B1(new_n702_), .B2(G106gat), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n701_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g506(.A(KEYINPUT122), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT57), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n574_), .A2(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n321_), .B1(new_n338_), .B2(new_n339_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n344_), .A2(new_n337_), .A3(new_n322_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n349_), .A3(new_n712_), .ZN(new_n713_));
  XOR2_X1   g512(.A(new_n713_), .B(KEYINPUT120), .Z(new_n714_));
  NAND3_X1  g513(.A1(new_n714_), .A2(new_n315_), .A3(new_n355_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n362_), .A2(new_n314_), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n296_), .A2(new_n303_), .A3(new_n290_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n304_), .A2(KEYINPUT55), .ZN(new_n718_));
  INV_X1    g517(.A(KEYINPUT55), .ZN(new_n719_));
  NAND4_X1  g518(.A1(new_n296_), .A2(new_n297_), .A3(new_n719_), .A4(new_n303_), .ZN(new_n720_));
  AOI221_X4 g519(.A(KEYINPUT118), .B1(new_n293_), .B2(new_n717_), .C1(new_n718_), .C2(new_n720_), .ZN(new_n721_));
  INV_X1    g520(.A(KEYINPUT118), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n718_), .A2(new_n720_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n717_), .A2(new_n293_), .ZN(new_n724_));
  AOI21_X1  g523(.A(new_n722_), .B1(new_n723_), .B2(new_n724_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n311_), .B1(new_n721_), .B2(new_n725_), .ZN(new_n726_));
  INV_X1    g525(.A(KEYINPUT56), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n726_), .A2(new_n727_), .ZN(new_n728_));
  OAI211_X1 g527(.A(KEYINPUT56), .B(new_n311_), .C1(new_n721_), .C2(new_n725_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n716_), .B1(new_n728_), .B2(new_n729_), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n715_), .B1(new_n730_), .B2(KEYINPUT119), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT119), .ZN(new_n732_));
  AOI211_X1 g531(.A(new_n732_), .B(new_n716_), .C1(new_n728_), .C2(new_n729_), .ZN(new_n733_));
  OAI21_X1  g532(.A(new_n710_), .B1(new_n731_), .B2(new_n733_), .ZN(new_n734_));
  AND3_X1   g533(.A1(new_n714_), .A2(new_n314_), .A3(new_n355_), .ZN(new_n735_));
  NAND2_X1  g534(.A1(new_n284_), .A2(new_n287_), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n301_), .B1(new_n736_), .B2(new_n225_), .ZN(new_n737_));
  AOI21_X1  g536(.A(new_n737_), .B1(new_n276_), .B2(new_n295_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n719_), .B1(new_n738_), .B2(new_n297_), .ZN(new_n739_));
  INV_X1    g538(.A(new_n720_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n724_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(KEYINPUT118), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n723_), .A2(new_n722_), .A3(new_n724_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n742_), .A2(new_n743_), .ZN(new_n744_));
  AOI21_X1  g543(.A(KEYINPUT56), .B1(new_n744_), .B2(new_n311_), .ZN(new_n745_));
  AOI211_X1 g544(.A(new_n727_), .B(new_n313_), .C1(new_n742_), .C2(new_n743_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n735_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT58), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n584_), .B1(new_n747_), .B2(new_n748_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n728_), .A2(new_n729_), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n750_), .A2(KEYINPUT121), .A3(KEYINPUT58), .A4(new_n735_), .ZN(new_n751_));
  OAI211_X1 g550(.A(KEYINPUT58), .B(new_n735_), .C1(new_n745_), .C2(new_n746_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT121), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n752_), .A2(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n749_), .A2(new_n751_), .A3(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n734_), .A2(new_n755_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n716_), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n757_), .B1(new_n745_), .B2(new_n746_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n758_), .A2(new_n732_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n730_), .A2(KEYINPUT119), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n759_), .A2(new_n760_), .A3(new_n715_), .ZN(new_n761_));
  AOI21_X1  g560(.A(KEYINPUT57), .B1(new_n761_), .B2(new_n615_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n708_), .B1(new_n756_), .B2(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n615_), .B1(new_n731_), .B2(new_n733_), .ZN(new_n764_));
  NAND2_X1  g563(.A1(new_n764_), .A2(new_n709_), .ZN(new_n765_));
  NAND4_X1  g564(.A1(new_n765_), .A2(KEYINPUT122), .A3(new_n734_), .A4(new_n755_), .ZN(new_n766_));
  NAND3_X1  g565(.A1(new_n763_), .A2(new_n383_), .A3(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n586_), .A2(new_n579_), .ZN(new_n768_));
  XNOR2_X1  g567(.A(new_n768_), .B(KEYINPUT54), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT123), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n770_), .A2(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n767_), .A2(KEYINPUT123), .A3(new_n769_), .ZN(new_n773_));
  NOR3_X1   g572(.A1(new_n538_), .A2(new_n438_), .A3(new_n592_), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n772_), .A2(new_n362_), .A3(new_n773_), .A4(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(G113gat), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n777_), .A2(KEYINPUT124), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT124), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n775_), .A2(new_n779_), .A3(new_n776_), .ZN(new_n780_));
  INV_X1    g579(.A(new_n769_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n383_), .B1(new_n756_), .B2(new_n762_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n781_), .A2(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n774_), .ZN(new_n785_));
  NOR3_X1   g584(.A1(new_n784_), .A2(KEYINPUT59), .A3(new_n785_), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n772_), .A2(new_n773_), .A3(new_n774_), .ZN(new_n787_));
  AOI21_X1  g586(.A(new_n786_), .B1(new_n787_), .B2(KEYINPUT59), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n579_), .A2(new_n776_), .ZN(new_n789_));
  AOI22_X1  g588(.A1(new_n778_), .A2(new_n780_), .B1(new_n788_), .B2(new_n789_), .ZN(G1340gat));
  AND3_X1   g589(.A1(new_n767_), .A2(KEYINPUT123), .A3(new_n769_), .ZN(new_n791_));
  AOI21_X1  g590(.A(KEYINPUT123), .B1(new_n767_), .B2(new_n769_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(new_n792_), .ZN(new_n793_));
  NOR2_X1   g592(.A1(new_n320_), .A2(KEYINPUT60), .ZN(new_n794_));
  INV_X1    g593(.A(G120gat), .ZN(new_n795_));
  MUX2_X1   g594(.A(KEYINPUT60), .B(new_n794_), .S(new_n795_), .Z(new_n796_));
  NAND4_X1  g595(.A1(new_n793_), .A2(KEYINPUT125), .A3(new_n774_), .A4(new_n796_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n772_), .A2(new_n773_), .A3(new_n774_), .A4(new_n796_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT125), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(new_n799_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n797_), .A2(new_n800_), .ZN(new_n801_));
  AOI211_X1 g600(.A(new_n320_), .B(new_n786_), .C1(new_n787_), .C2(KEYINPUT59), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n801_), .B1(new_n802_), .B2(new_n795_), .ZN(G1341gat));
  INV_X1    g602(.A(new_n787_), .ZN(new_n804_));
  INV_X1    g603(.A(G127gat), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n804_), .A2(new_n805_), .A3(new_n384_), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n383_), .B(new_n786_), .C1(new_n787_), .C2(KEYINPUT59), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n805_), .ZN(G1342gat));
  INV_X1    g607(.A(G134gat), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n804_), .A2(new_n809_), .A3(new_n574_), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n584_), .B(new_n786_), .C1(new_n787_), .C2(KEYINPUT59), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n810_), .B1(new_n811_), .B2(new_n809_), .ZN(G1343gat));
  NOR3_X1   g611(.A1(new_n791_), .A2(new_n792_), .A3(new_n536_), .ZN(new_n813_));
  NOR2_X1   g612(.A1(new_n641_), .A2(new_n438_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n813_), .A2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n362_), .ZN(new_n816_));
  OAI21_X1  g615(.A(G141gat), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(G141gat), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n813_), .A2(new_n818_), .A3(new_n362_), .A4(new_n814_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n817_), .A2(new_n819_), .ZN(G1344gat));
  OAI21_X1  g619(.A(G148gat), .B1(new_n815_), .B2(new_n320_), .ZN(new_n821_));
  INV_X1    g620(.A(G148gat), .ZN(new_n822_));
  NAND4_X1  g621(.A1(new_n813_), .A2(new_n822_), .A3(new_n319_), .A4(new_n814_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n821_), .A2(new_n823_), .ZN(G1345gat));
  XNOR2_X1  g623(.A(KEYINPUT61), .B(G155gat), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n825_), .B1(new_n815_), .B2(new_n383_), .ZN(new_n826_));
  INV_X1    g625(.A(new_n825_), .ZN(new_n827_));
  NAND4_X1  g626(.A1(new_n813_), .A2(new_n384_), .A3(new_n814_), .A4(new_n827_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n826_), .A2(new_n828_), .ZN(G1346gat));
  OAI21_X1  g628(.A(G162gat), .B1(new_n815_), .B2(new_n584_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n615_), .A2(G162gat), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n813_), .A2(new_n814_), .A3(new_n831_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n830_), .A2(new_n832_), .ZN(G1347gat));
  NAND2_X1  g632(.A1(new_n641_), .A2(new_n438_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(new_n537_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n836_), .ZN(new_n837_));
  OAI211_X1 g636(.A(new_n362_), .B(new_n837_), .C1(new_n781_), .C2(new_n783_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n838_), .A2(G169gat), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT126), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT126), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n838_), .A2(new_n841_), .A3(G169gat), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  INV_X1    g642(.A(KEYINPUT62), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n843_), .A2(new_n844_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n840_), .A2(new_n842_), .A3(KEYINPUT62), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n784_), .A2(new_n836_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n847_), .A2(new_n362_), .A3(new_n473_), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n845_), .A2(new_n846_), .A3(new_n848_), .ZN(G1348gat));
  AOI21_X1  g648(.A(G176gat), .B1(new_n847_), .B2(new_n319_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n791_), .A2(new_n792_), .A3(new_n553_), .ZN(new_n851_));
  NOR4_X1   g650(.A1(new_n834_), .A2(new_n457_), .A3(new_n320_), .A4(new_n533_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n850_), .B1(new_n851_), .B2(new_n852_), .ZN(G1349gat));
  INV_X1    g652(.A(new_n847_), .ZN(new_n854_));
  NOR3_X1   g653(.A1(new_n854_), .A2(new_n383_), .A3(new_n460_), .ZN(new_n855_));
  NAND4_X1  g654(.A1(new_n851_), .A2(new_n384_), .A3(new_n534_), .A4(new_n835_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n855_), .B1(new_n856_), .B2(new_n470_), .ZN(G1350gat));
  OAI21_X1  g656(.A(G190gat), .B1(new_n854_), .B2(new_n584_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n574_), .A2(new_n462_), .A3(new_n463_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n854_), .B2(new_n859_), .ZN(G1351gat));
  NAND4_X1  g659(.A1(new_n813_), .A2(G197gat), .A3(new_n362_), .A4(new_n835_), .ZN(new_n861_));
  NAND4_X1  g660(.A1(new_n772_), .A2(new_n535_), .A3(new_n773_), .A4(new_n835_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n443_), .B1(new_n862_), .B2(new_n816_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n861_), .A2(new_n863_), .ZN(G1352gat));
  NAND4_X1  g663(.A1(new_n813_), .A2(new_n319_), .A3(new_n441_), .A4(new_n835_), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n444_), .B1(new_n862_), .B2(new_n320_), .ZN(new_n866_));
  AND2_X1   g665(.A1(new_n865_), .A2(new_n866_), .ZN(G1353gat));
  INV_X1    g666(.A(KEYINPUT63), .ZN(new_n868_));
  INV_X1    g667(.A(G211gat), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n384_), .B1(new_n868_), .B2(new_n869_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(new_n870_), .B(KEYINPUT127), .ZN(new_n871_));
  INV_X1    g670(.A(new_n871_), .ZN(new_n872_));
  OAI211_X1 g671(.A(new_n868_), .B(new_n869_), .C1(new_n862_), .C2(new_n872_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n868_), .A2(new_n869_), .ZN(new_n874_));
  NAND4_X1  g673(.A1(new_n813_), .A2(new_n835_), .A3(new_n874_), .A4(new_n871_), .ZN(new_n875_));
  AND2_X1   g674(.A1(new_n873_), .A2(new_n875_), .ZN(G1354gat));
  OAI21_X1  g675(.A(G218gat), .B1(new_n862_), .B2(new_n584_), .ZN(new_n877_));
  OR2_X1    g676(.A1(new_n615_), .A2(G218gat), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n877_), .B1(new_n862_), .B2(new_n878_), .ZN(G1355gat));
endmodule


