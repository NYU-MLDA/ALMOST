//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n658_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n760_,
    new_n761_, new_n762_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n849_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_;
  XOR2_X1   g000(.A(G127gat), .B(G134gat), .Z(new_n202_));
  INV_X1    g001(.A(G120gat), .ZN(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G113gat), .ZN(new_n204_));
  INV_X1    g003(.A(G113gat), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(G120gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n204_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n202_), .A2(new_n207_), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G127gat), .B(G134gat), .ZN(new_n209_));
  NAND3_X1  g008(.A1(new_n209_), .A2(new_n204_), .A3(new_n206_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n208_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n211_), .B(KEYINPUT31), .ZN(new_n212_));
  XNOR2_X1  g011(.A(KEYINPUT26), .B(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT80), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT25), .ZN(new_n215_));
  NAND3_X1  g014(.A1(new_n214_), .A2(new_n215_), .A3(G183gat), .ZN(new_n216_));
  INV_X1    g015(.A(G183gat), .ZN(new_n217_));
  OAI21_X1  g016(.A(KEYINPUT25), .B1(new_n217_), .B2(KEYINPUT80), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n213_), .A2(new_n216_), .A3(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(G169gat), .ZN(new_n220_));
  INV_X1    g019(.A(G176gat), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n220_), .A2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n222_), .A2(KEYINPUT24), .A3(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(KEYINPUT81), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n219_), .A2(KEYINPUT81), .A3(new_n224_), .ZN(new_n228_));
  AND3_X1   g027(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n229_));
  AOI21_X1  g028(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT24), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n232_), .A2(new_n220_), .A3(new_n221_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT82), .ZN(new_n235_));
  NAND2_X1  g034(.A1(G183gat), .A2(G190gat), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT23), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n239_));
  AND3_X1   g038(.A1(new_n233_), .A2(new_n238_), .A3(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(KEYINPUT82), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  NAND4_X1  g041(.A1(new_n227_), .A2(new_n228_), .A3(new_n235_), .A4(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n220_), .A2(KEYINPUT22), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT22), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n245_), .A2(G169gat), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n244_), .A2(new_n246_), .A3(new_n221_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT83), .ZN(new_n248_));
  INV_X1    g047(.A(G190gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n217_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n238_), .A2(new_n250_), .A3(new_n239_), .ZN(new_n251_));
  NAND3_X1  g050(.A1(new_n248_), .A2(new_n251_), .A3(new_n223_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n243_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(G71gat), .B(G99gat), .ZN(new_n254_));
  XNOR2_X1  g053(.A(new_n254_), .B(G43gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(new_n253_), .B(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(G227gat), .A2(G233gat), .ZN(new_n257_));
  INV_X1    g056(.A(G15gat), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n259_), .B(KEYINPUT30), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n256_), .B(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n212_), .B1(new_n261_), .B2(KEYINPUT84), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n262_), .B1(KEYINPUT84), .B2(new_n261_), .ZN(new_n263_));
  NOR2_X1   g062(.A1(new_n261_), .A2(KEYINPUT84), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n264_), .A2(new_n212_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n215_), .A2(G183gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n249_), .A2(KEYINPUT26), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT26), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(G190gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n217_), .A2(KEYINPUT25), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n267_), .A2(new_n268_), .A3(new_n270_), .A4(new_n271_), .ZN(new_n272_));
  NAND4_X1  g071(.A1(new_n272_), .A2(new_n231_), .A3(new_n224_), .A4(new_n233_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT91), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND4_X1  g074(.A1(new_n240_), .A2(KEYINPUT91), .A3(new_n224_), .A4(new_n272_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n223_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT22), .B(G169gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n277_), .B1(new_n278_), .B2(new_n221_), .ZN(new_n279_));
  AOI21_X1  g078(.A(KEYINPUT92), .B1(new_n279_), .B2(new_n251_), .ZN(new_n280_));
  AND4_X1   g079(.A1(KEYINPUT92), .A2(new_n251_), .A3(new_n223_), .A4(new_n247_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n275_), .B(new_n276_), .C1(new_n280_), .C2(new_n281_), .ZN(new_n282_));
  OR2_X1    g081(.A1(G197gat), .A2(G204gat), .ZN(new_n283_));
  NAND2_X1  g082(.A1(G197gat), .A2(G204gat), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n283_), .A2(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(G211gat), .B(G218gat), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n285_), .B(KEYINPUT21), .C1(new_n286_), .C2(KEYINPUT88), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT21), .ZN(new_n288_));
  XOR2_X1   g087(.A(G211gat), .B(G218gat), .Z(new_n289_));
  INV_X1    g088(.A(KEYINPUT88), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n283_), .B(new_n284_), .C1(new_n286_), .C2(KEYINPUT21), .ZN(new_n292_));
  OAI21_X1  g091(.A(new_n287_), .B1(new_n291_), .B2(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n282_), .A2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n293_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n227_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n228_), .A2(new_n235_), .A3(new_n242_), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n295_), .B(new_n252_), .C1(new_n296_), .C2(new_n297_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n294_), .A2(new_n298_), .A3(KEYINPUT20), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G226gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT19), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(KEYINPUT20), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n301_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n304_), .B1(new_n282_), .B2(new_n293_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n295_), .B1(new_n243_), .B2(new_n252_), .ZN(new_n306_));
  OR2_X1    g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(G8gat), .B(G36gat), .Z(new_n308_));
  XNOR2_X1  g107(.A(KEYINPUT93), .B(KEYINPUT18), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n308_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G64gat), .B(G92gat), .ZN(new_n311_));
  XNOR2_X1  g110(.A(new_n310_), .B(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n302_), .A2(new_n307_), .A3(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n312_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n301_), .ZN(new_n315_));
  AOI21_X1  g114(.A(new_n303_), .B1(new_n282_), .B2(new_n293_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n315_), .B1(new_n316_), .B2(new_n298_), .ZN(new_n317_));
  NOR2_X1   g116(.A1(new_n305_), .A2(new_n306_), .ZN(new_n318_));
  OAI21_X1  g117(.A(new_n314_), .B1(new_n317_), .B2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n313_), .A2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT27), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  XOR2_X1   g121(.A(new_n312_), .B(KEYINPUT98), .Z(new_n323_));
  NOR2_X1   g122(.A1(new_n299_), .A2(new_n301_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n253_), .A2(new_n293_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n279_), .A2(new_n251_), .ZN(new_n326_));
  AOI21_X1  g125(.A(KEYINPUT96), .B1(new_n326_), .B2(new_n273_), .ZN(new_n327_));
  NOR2_X1   g126(.A1(new_n327_), .A2(new_n293_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n273_), .A3(KEYINPUT96), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n303_), .B1(new_n328_), .B2(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n315_), .B1(new_n325_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n323_), .B1(new_n324_), .B2(new_n331_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n332_), .A2(KEYINPUT27), .A3(new_n313_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n322_), .A2(new_n333_), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G78gat), .B(G106gat), .ZN(new_n336_));
  XNOR2_X1  g135(.A(new_n336_), .B(KEYINPUT89), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(G155gat), .A2(G162gat), .ZN(new_n339_));
  INV_X1    g138(.A(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(G155gat), .A2(G162gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  INV_X1    g141(.A(new_n342_), .ZN(new_n343_));
  OAI21_X1  g142(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(KEYINPUT85), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT85), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n346_), .B(KEYINPUT3), .C1(G141gat), .C2(G148gat), .ZN(new_n347_));
  AND2_X1   g146(.A1(new_n345_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(G141gat), .A2(G148gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT2), .ZN(new_n350_));
  INV_X1    g149(.A(KEYINPUT2), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(G141gat), .A3(G148gat), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT3), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G141gat), .A2(G148gat), .ZN(new_n354_));
  AOI22_X1  g153(.A1(new_n350_), .A2(new_n352_), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  AOI21_X1  g154(.A(new_n343_), .B1(new_n348_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n339_), .A2(KEYINPUT1), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT1), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(G155gat), .A3(G162gat), .ZN(new_n359_));
  OAI211_X1 g158(.A(new_n357_), .B(new_n359_), .C1(G155gat), .C2(G162gat), .ZN(new_n360_));
  INV_X1    g159(.A(new_n349_), .ZN(new_n361_));
  NOR2_X1   g160(.A1(new_n361_), .A2(new_n354_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n360_), .A2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(new_n363_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n356_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366_));
  OAI21_X1  g165(.A(new_n293_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n367_));
  AND2_X1   g166(.A1(G228gat), .A2(G233gat), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n368_), .B1(new_n293_), .B2(KEYINPUT87), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(new_n369_), .ZN(new_n370_));
  OAI221_X1 g169(.A(new_n293_), .B1(KEYINPUT87), .B2(new_n368_), .C1(new_n365_), .C2(new_n366_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n338_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n372_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n370_), .A2(new_n371_), .A3(new_n338_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n373_), .A2(new_n374_), .ZN(new_n375_));
  NOR2_X1   g174(.A1(new_n372_), .A2(KEYINPUT90), .ZN(new_n376_));
  XOR2_X1   g175(.A(G22gat), .B(G50gat), .Z(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  XNOR2_X1  g177(.A(KEYINPUT86), .B(KEYINPUT28), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  NAND3_X1  g179(.A1(new_n365_), .A2(new_n366_), .A3(new_n380_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n380_), .B1(new_n365_), .B2(new_n366_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n378_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(new_n383_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n385_), .A2(new_n377_), .A3(new_n381_), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(new_n386_), .ZN(new_n387_));
  OAI21_X1  g186(.A(new_n375_), .B1(new_n376_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n387_), .ZN(new_n389_));
  NAND4_X1  g188(.A1(new_n389_), .A2(KEYINPUT90), .A3(new_n373_), .A4(new_n374_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n335_), .A2(new_n391_), .ZN(new_n392_));
  AND2_X1   g191(.A1(new_n208_), .A2(new_n210_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n393_), .B1(new_n356_), .B2(new_n364_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n354_), .A2(new_n353_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n351_), .B1(G141gat), .B2(G148gat), .ZN(new_n396_));
  NOR2_X1   g195(.A1(new_n349_), .A2(KEYINPUT2), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n395_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n345_), .A2(new_n347_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n342_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  NAND3_X1  g199(.A1(new_n400_), .A2(new_n363_), .A3(new_n211_), .ZN(new_n401_));
  NAND3_X1  g200(.A1(new_n394_), .A2(KEYINPUT4), .A3(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403_));
  AOI21_X1  g202(.A(new_n211_), .B1(new_n400_), .B2(new_n363_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n403_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n406_));
  AND3_X1   g205(.A1(new_n400_), .A2(new_n211_), .A3(new_n363_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n407_), .A2(new_n404_), .ZN(new_n408_));
  AOI22_X1  g207(.A1(new_n402_), .A2(new_n406_), .B1(new_n408_), .B2(new_n403_), .ZN(new_n409_));
  XNOR2_X1  g208(.A(G1gat), .B(G29gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(G85gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(KEYINPUT0), .B(G57gat), .Z(new_n412_));
  XNOR2_X1  g211(.A(new_n411_), .B(new_n412_), .ZN(new_n413_));
  OR2_X1    g212(.A1(new_n409_), .A2(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n413_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NOR3_X1   g215(.A1(new_n266_), .A2(new_n392_), .A3(new_n416_), .ZN(new_n417_));
  NOR3_X1   g216(.A1(new_n334_), .A2(new_n391_), .A3(new_n416_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n313_), .A2(KEYINPUT94), .A3(new_n319_), .ZN(new_n419_));
  AOI21_X1  g218(.A(KEYINPUT94), .B1(new_n313_), .B2(new_n319_), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT33), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n421_), .B1(new_n409_), .B2(new_n413_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n406_), .A2(new_n402_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n394_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n424_));
  AND4_X1   g223(.A1(new_n421_), .A2(new_n423_), .A3(new_n424_), .A4(new_n413_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n403_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n404_), .B2(new_n405_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n427_), .A2(new_n402_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT95), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n394_), .A2(new_n401_), .A3(new_n426_), .ZN(new_n430_));
  XOR2_X1   g229(.A(new_n411_), .B(new_n412_), .Z(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n428_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n433_));
  AOI21_X1  g232(.A(new_n413_), .B1(new_n408_), .B2(new_n426_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n402_), .ZN(new_n435_));
  AOI21_X1  g234(.A(KEYINPUT95), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  OAI22_X1  g235(.A1(new_n422_), .A2(new_n425_), .B1(new_n433_), .B2(new_n436_), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n419_), .A2(new_n420_), .A3(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n312_), .A2(KEYINPUT32), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n302_), .A2(new_n307_), .A3(new_n439_), .ZN(new_n440_));
  OAI211_X1 g239(.A(KEYINPUT32), .B(new_n312_), .C1(new_n324_), .C2(new_n331_), .ZN(new_n441_));
  NAND3_X1  g240(.A1(new_n416_), .A2(new_n440_), .A3(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  OAI21_X1  g242(.A(new_n391_), .B1(new_n438_), .B2(new_n443_), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n418_), .B1(new_n444_), .B2(KEYINPUT97), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n388_), .A2(new_n390_), .ZN(new_n446_));
  INV_X1    g245(.A(new_n420_), .ZN(new_n447_));
  INV_X1    g246(.A(new_n437_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n313_), .A2(new_n319_), .A3(KEYINPUT94), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n447_), .A2(new_n448_), .A3(new_n449_), .ZN(new_n450_));
  AOI21_X1  g249(.A(new_n446_), .B1(new_n450_), .B2(new_n442_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT97), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n445_), .A2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n417_), .B1(new_n454_), .B2(new_n266_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(G230gat), .A2(G233gat), .ZN(new_n456_));
  XOR2_X1   g255(.A(new_n456_), .B(KEYINPUT64), .Z(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  OR2_X1    g257(.A1(G85gat), .A2(G92gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  AND2_X1   g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(G99gat), .ZN(new_n462_));
  INV_X1    g261(.A(G106gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n464_), .B(KEYINPUT7), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G99gat), .A2(G106gat), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  OAI21_X1  g267(.A(new_n461_), .B1(new_n465_), .B2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(KEYINPUT67), .A2(KEYINPUT8), .ZN(new_n470_));
  INV_X1    g269(.A(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n469_), .B(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT9), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n459_), .B1(new_n473_), .B2(new_n460_), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n460_), .A2(new_n473_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT65), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n475_), .A2(new_n476_), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n460_), .A2(KEYINPUT65), .A3(new_n473_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n474_), .B1(new_n477_), .B2(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n468_), .ZN(new_n481_));
  XOR2_X1   g280(.A(KEYINPUT10), .B(G99gat), .Z(new_n482_));
  NAND2_X1  g281(.A1(new_n482_), .A2(new_n463_), .ZN(new_n483_));
  NAND4_X1  g282(.A1(new_n480_), .A2(KEYINPUT66), .A3(new_n481_), .A4(new_n483_), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT66), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n481_), .A2(new_n483_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n485_), .B1(new_n486_), .B2(new_n479_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n472_), .A2(new_n484_), .A3(new_n487_), .ZN(new_n488_));
  XOR2_X1   g287(.A(G71gat), .B(G78gat), .Z(new_n489_));
  XNOR2_X1  g288(.A(G57gat), .B(G64gat), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n489_), .B1(KEYINPUT11), .B2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT68), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n492_), .A3(KEYINPUT11), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n492_), .B1(new_n490_), .B2(KEYINPUT11), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n491_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n490_), .A2(KEYINPUT11), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(KEYINPUT68), .ZN(new_n498_));
  OR2_X1    g297(.A1(new_n490_), .A2(KEYINPUT11), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n498_), .A2(new_n499_), .A3(new_n489_), .A4(new_n493_), .ZN(new_n500_));
  AND2_X1   g299(.A1(new_n496_), .A2(new_n500_), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT12), .B1(new_n488_), .B2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n488_), .A2(new_n501_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n502_), .A2(new_n503_), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n469_), .B(new_n470_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n484_), .A2(new_n487_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT69), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  NAND3_X1  g307(.A1(new_n484_), .A2(KEYINPUT69), .A3(new_n487_), .ZN(new_n509_));
  AOI21_X1  g308(.A(new_n505_), .B1(new_n508_), .B2(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(KEYINPUT70), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n501_), .A2(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n511_), .B1(new_n496_), .B2(new_n500_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n512_), .A2(KEYINPUT12), .A3(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT71), .ZN(new_n516_));
  NOR3_X1   g315(.A1(new_n510_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n484_), .A2(KEYINPUT69), .A3(new_n487_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT69), .B1(new_n484_), .B2(new_n487_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n472_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n496_), .A2(new_n500_), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT12), .B1(new_n521_), .B2(KEYINPUT70), .ZN(new_n522_));
  NOR2_X1   g321(.A1(new_n522_), .A2(new_n513_), .ZN(new_n523_));
  AOI21_X1  g322(.A(KEYINPUT71), .B1(new_n520_), .B2(new_n523_), .ZN(new_n524_));
  OAI211_X1 g323(.A(new_n458_), .B(new_n504_), .C1(new_n517_), .C2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(new_n503_), .ZN(new_n526_));
  NOR2_X1   g325(.A1(new_n488_), .A2(new_n501_), .ZN(new_n527_));
  OAI21_X1  g326(.A(new_n457_), .B1(new_n526_), .B2(new_n527_), .ZN(new_n528_));
  XOR2_X1   g327(.A(G120gat), .B(G148gat), .Z(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT72), .B(KEYINPUT5), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n529_), .B(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n531_), .B(new_n532_), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n525_), .A2(new_n528_), .A3(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  AOI21_X1  g334(.A(new_n533_), .B1(new_n525_), .B2(new_n528_), .ZN(new_n536_));
  OAI21_X1  g335(.A(KEYINPUT13), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n536_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT13), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(new_n534_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n537_), .A2(new_n540_), .ZN(new_n541_));
  INV_X1    g340(.A(KEYINPUT14), .ZN(new_n542_));
  XNOR2_X1  g341(.A(KEYINPUT76), .B(G8gat), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n542_), .B1(new_n543_), .B2(G1gat), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT77), .ZN(new_n545_));
  XNOR2_X1  g344(.A(new_n544_), .B(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n546_), .A2(new_n547_), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G1gat), .B(G8gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G29gat), .B(G36gat), .ZN(new_n551_));
  XNOR2_X1  g350(.A(G43gat), .B(G50gat), .ZN(new_n552_));
  XNOR2_X1  g351(.A(new_n551_), .B(new_n552_), .ZN(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(KEYINPUT79), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n550_), .B(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(G229gat), .A2(G233gat), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n550_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n554_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n553_), .B(KEYINPUT15), .ZN(new_n560_));
  NAND2_X1  g359(.A1(new_n550_), .A2(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n559_), .A2(new_n561_), .A3(new_n556_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G113gat), .B(G141gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(G169gat), .B(G197gat), .ZN(new_n564_));
  XOR2_X1   g363(.A(new_n563_), .B(new_n564_), .Z(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  OR3_X1    g365(.A1(new_n557_), .A2(new_n562_), .A3(new_n566_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n566_), .B1(new_n557_), .B2(new_n562_), .ZN(new_n568_));
  NAND2_X1  g367(.A1(new_n567_), .A2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n541_), .A2(new_n569_), .ZN(new_n570_));
  NOR2_X1   g369(.A1(new_n455_), .A2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(G190gat), .B(G218gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(G134gat), .B(G162gat), .ZN(new_n573_));
  XNOR2_X1  g372(.A(new_n572_), .B(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(KEYINPUT75), .B(KEYINPUT36), .ZN(new_n575_));
  XOR2_X1   g374(.A(new_n574_), .B(new_n575_), .Z(new_n576_));
  INV_X1    g375(.A(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n578_), .B(KEYINPUT34), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT35), .ZN(new_n581_));
  NOR2_X1   g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n520_), .A2(new_n560_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n505_), .A2(new_n506_), .ZN(new_n585_));
  AOI22_X1  g384(.A1(new_n585_), .A2(new_n553_), .B1(new_n581_), .B2(new_n580_), .ZN(new_n586_));
  AOI21_X1  g385(.A(new_n583_), .B1(new_n584_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  NAND3_X1  g387(.A1(new_n584_), .A2(new_n586_), .A3(new_n583_), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n577_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  INV_X1    g389(.A(KEYINPUT74), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT37), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n589_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n576_), .B1(new_n593_), .B2(new_n587_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(KEYINPUT73), .B(KEYINPUT36), .ZN(new_n595_));
  NOR2_X1   g394(.A1(new_n574_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n588_), .A2(new_n589_), .A3(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n594_), .A2(new_n597_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(new_n592_), .B(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n521_), .B(new_n600_), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n550_), .B(new_n601_), .ZN(new_n602_));
  XOR2_X1   g401(.A(G127gat), .B(G155gat), .Z(new_n603_));
  XNOR2_X1  g402(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G183gat), .B(G211gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n605_), .B(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(KEYINPUT70), .A2(KEYINPUT17), .ZN(new_n609_));
  AOI21_X1  g408(.A(new_n602_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n609_), .ZN(new_n611_));
  OAI21_X1  g410(.A(new_n611_), .B1(KEYINPUT17), .B2(new_n608_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n602_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n610_), .A2(new_n613_), .ZN(new_n614_));
  NOR2_X1   g413(.A1(new_n599_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n571_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT99), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT99), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n571_), .A2(new_n618_), .A3(new_n615_), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(G1gat), .ZN(new_n621_));
  NAND3_X1  g420(.A1(new_n620_), .A2(new_n621_), .A3(new_n416_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT38), .ZN(new_n623_));
  AND2_X1   g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n598_), .ZN(new_n625_));
  NOR2_X1   g424(.A1(new_n455_), .A2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n570_), .A2(new_n614_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT100), .Z(new_n629_));
  AOI21_X1  g428(.A(new_n621_), .B1(new_n629_), .B2(new_n416_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n624_), .A2(new_n630_), .ZN(new_n631_));
  OAI21_X1  g430(.A(new_n631_), .B1(new_n623_), .B2(new_n622_), .ZN(G1324gat));
  NAND3_X1  g431(.A1(new_n626_), .A2(new_n334_), .A3(new_n627_), .ZN(new_n633_));
  AOI21_X1  g432(.A(KEYINPUT101), .B1(new_n633_), .B2(G8gat), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT39), .ZN(new_n635_));
  NOR2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n633_), .A2(G8gat), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n636_), .B1(new_n637_), .B2(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n634_), .A2(new_n635_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n335_), .A2(new_n543_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n617_), .A2(new_n619_), .A3(new_n642_), .ZN(new_n643_));
  NAND4_X1  g442(.A1(new_n639_), .A2(new_n640_), .A3(new_n641_), .A4(new_n643_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n638_), .A2(new_n637_), .ZN(new_n645_));
  NOR3_X1   g444(.A1(new_n645_), .A2(new_n635_), .A3(new_n634_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n641_), .A2(new_n643_), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT40), .B1(new_n646_), .B2(new_n647_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n644_), .A2(new_n648_), .ZN(new_n649_));
  XNOR2_X1  g448(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n650_));
  INV_X1    g449(.A(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n644_), .A2(new_n648_), .A3(new_n650_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(G1325gat));
  INV_X1    g453(.A(new_n266_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n258_), .B1(new_n629_), .B2(new_n655_), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n656_), .B(KEYINPUT41), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n620_), .A2(new_n258_), .A3(new_n655_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(G1326gat));
  INV_X1    g458(.A(G22gat), .ZN(new_n660_));
  XNOR2_X1  g459(.A(new_n446_), .B(KEYINPUT104), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n629_), .B2(new_n661_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT42), .Z(new_n663_));
  NAND3_X1  g462(.A1(new_n620_), .A2(new_n660_), .A3(new_n661_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1327gat));
  INV_X1    g464(.A(new_n614_), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n666_), .A2(new_n598_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n571_), .A2(new_n667_), .ZN(new_n668_));
  AOI21_X1  g467(.A(G29gat), .B1(new_n668_), .B2(new_n416_), .ZN(new_n669_));
  INV_X1    g468(.A(KEYINPUT43), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n655_), .B1(new_n445_), .B2(new_n453_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n670_), .B(new_n599_), .C1(new_n671_), .C2(new_n417_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n391_), .A2(new_n416_), .ZN(new_n675_));
  NAND2_X1  g474(.A1(new_n675_), .A2(new_n335_), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(new_n451_), .B2(new_n452_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n444_), .A2(KEYINPUT97), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n266_), .B1(new_n677_), .B2(new_n678_), .ZN(new_n679_));
  INV_X1    g478(.A(new_n417_), .ZN(new_n680_));
  NAND2_X1  g479(.A1(new_n679_), .A2(new_n680_), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n681_), .A2(KEYINPUT105), .A3(new_n670_), .A4(new_n599_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n599_), .ZN(new_n683_));
  OAI21_X1  g482(.A(KEYINPUT43), .B1(new_n455_), .B2(new_n683_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n674_), .A2(new_n682_), .A3(new_n684_), .ZN(new_n685_));
  NOR2_X1   g484(.A1(new_n570_), .A2(new_n666_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n688_));
  AOI21_X1  g487(.A(KEYINPUT106), .B1(new_n687_), .B2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n690_));
  AOI211_X1 g489(.A(new_n690_), .B(KEYINPUT44), .C1(new_n685_), .C2(new_n686_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n689_), .A2(new_n691_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n685_), .A2(KEYINPUT44), .A3(new_n686_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n692_), .A2(new_n693_), .ZN(new_n694_));
  AND2_X1   g493(.A1(new_n416_), .A2(G29gat), .ZN(new_n695_));
  AOI21_X1  g494(.A(new_n669_), .B1(new_n694_), .B2(new_n695_), .ZN(G1328gat));
  XNOR2_X1  g495(.A(KEYINPUT107), .B(KEYINPUT46), .ZN(new_n697_));
  OAI211_X1 g496(.A(new_n334_), .B(new_n693_), .C1(new_n689_), .C2(new_n691_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(G36gat), .ZN(new_n699_));
  INV_X1    g498(.A(G36gat), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n668_), .A2(new_n700_), .A3(new_n334_), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT45), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n701_), .B(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n703_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n697_), .B1(new_n699_), .B2(new_n704_), .ZN(new_n705_));
  INV_X1    g504(.A(new_n697_), .ZN(new_n706_));
  AOI211_X1 g505(.A(new_n703_), .B(new_n706_), .C1(new_n698_), .C2(G36gat), .ZN(new_n707_));
  NOR2_X1   g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1329gat));
  INV_X1    g507(.A(G43gat), .ZN(new_n709_));
  NOR2_X1   g508(.A1(new_n266_), .A2(new_n709_), .ZN(new_n710_));
  OAI211_X1 g509(.A(new_n693_), .B(new_n710_), .C1(new_n689_), .C2(new_n691_), .ZN(new_n711_));
  INV_X1    g510(.A(new_n668_), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n709_), .B1(new_n712_), .B2(new_n266_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n711_), .A2(new_n713_), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g514(.A(G50gat), .ZN(new_n716_));
  NAND3_X1  g515(.A1(new_n668_), .A2(new_n716_), .A3(new_n661_), .ZN(new_n717_));
  OAI211_X1 g516(.A(new_n446_), .B(new_n693_), .C1(new_n689_), .C2(new_n691_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n718_), .A2(KEYINPUT108), .A3(G50gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT108), .B1(new_n718_), .B2(G50gat), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n717_), .B1(new_n719_), .B2(new_n720_), .ZN(G1331gat));
  NAND3_X1  g520(.A1(new_n666_), .A2(new_n567_), .A3(new_n568_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n541_), .A2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n626_), .A2(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(G57gat), .ZN(new_n725_));
  INV_X1    g524(.A(new_n416_), .ZN(new_n726_));
  NOR3_X1   g525(.A1(new_n724_), .A2(new_n725_), .A3(new_n726_), .ZN(new_n727_));
  NOR3_X1   g526(.A1(new_n455_), .A2(new_n569_), .A3(new_n541_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(new_n615_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n726_), .B1(new_n729_), .B2(KEYINPUT109), .ZN(new_n730_));
  OAI21_X1  g529(.A(new_n730_), .B1(KEYINPUT109), .B2(new_n729_), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n727_), .B1(new_n731_), .B2(new_n725_), .ZN(G1332gat));
  OAI21_X1  g531(.A(G64gat), .B1(new_n724_), .B2(new_n335_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT48), .ZN(new_n734_));
  OR2_X1    g533(.A1(new_n335_), .A2(G64gat), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n734_), .B1(new_n729_), .B2(new_n735_), .ZN(G1333gat));
  OAI21_X1  g535(.A(G71gat), .B1(new_n724_), .B2(new_n266_), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n737_), .B(KEYINPUT49), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n266_), .A2(G71gat), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT110), .Z(new_n740_));
  OAI21_X1  g539(.A(new_n738_), .B1(new_n729_), .B2(new_n740_), .ZN(G1334gat));
  NAND3_X1  g540(.A1(new_n626_), .A2(new_n661_), .A3(new_n723_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(G78gat), .ZN(new_n743_));
  XNOR2_X1  g542(.A(new_n743_), .B(KEYINPUT50), .ZN(new_n744_));
  INV_X1    g543(.A(G78gat), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n661_), .A2(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(new_n744_), .B1(new_n729_), .B2(new_n746_), .ZN(G1335gat));
  NAND2_X1  g546(.A1(new_n728_), .A2(new_n667_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT111), .ZN(new_n749_));
  AOI21_X1  g548(.A(G85gat), .B1(new_n749_), .B2(new_n416_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n541_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n569_), .ZN(new_n752_));
  NAND3_X1  g551(.A1(new_n751_), .A2(new_n614_), .A3(new_n752_), .ZN(new_n753_));
  OR2_X1    g552(.A1(new_n685_), .A2(KEYINPUT112), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n685_), .A2(KEYINPUT112), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n753_), .B1(new_n754_), .B2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n416_), .A2(G85gat), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT113), .Z(new_n758_));
  AOI21_X1  g557(.A(new_n750_), .B1(new_n756_), .B2(new_n758_), .ZN(G1336gat));
  INV_X1    g558(.A(G92gat), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n749_), .A2(new_n760_), .A3(new_n334_), .ZN(new_n761_));
  AND2_X1   g560(.A1(new_n756_), .A2(new_n334_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n761_), .B1(new_n762_), .B2(new_n760_), .ZN(G1337gat));
  AOI21_X1  g562(.A(new_n462_), .B1(new_n756_), .B2(new_n655_), .ZN(new_n764_));
  AND3_X1   g563(.A1(new_n749_), .A2(new_n482_), .A3(new_n655_), .ZN(new_n765_));
  OR3_X1    g564(.A1(new_n764_), .A2(KEYINPUT51), .A3(new_n765_), .ZN(new_n766_));
  OAI21_X1  g565(.A(KEYINPUT51), .B1(new_n764_), .B2(new_n765_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n766_), .A2(new_n767_), .ZN(G1338gat));
  NOR2_X1   g567(.A1(new_n753_), .A2(new_n391_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n463_), .B1(new_n685_), .B2(new_n769_), .ZN(new_n770_));
  XOR2_X1   g569(.A(new_n770_), .B(KEYINPUT52), .Z(new_n771_));
  NAND3_X1  g570(.A1(new_n749_), .A2(new_n463_), .A3(new_n446_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(KEYINPUT114), .B(KEYINPUT53), .ZN(new_n773_));
  AND3_X1   g572(.A1(new_n771_), .A2(new_n772_), .A3(new_n773_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(new_n775_), .ZN(G1339gat));
  AOI21_X1  g575(.A(new_n722_), .B1(new_n537_), .B2(new_n540_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n599_), .B1(new_n777_), .B2(KEYINPUT115), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n541_), .A2(new_n666_), .A3(new_n752_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AND3_X1   g581(.A1(new_n778_), .A2(new_n779_), .A3(new_n782_), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n779_), .B1(new_n778_), .B2(new_n782_), .ZN(new_n784_));
  NOR2_X1   g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n569_), .A2(new_n534_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT116), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n525_), .A2(new_n787_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n788_), .A2(KEYINPUT55), .ZN(new_n789_));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n525_), .A2(new_n787_), .A3(new_n790_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n504_), .B1(new_n517_), .B2(new_n524_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n792_), .A2(new_n457_), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n789_), .A2(new_n791_), .A3(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n533_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n794_), .A2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT56), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND3_X1  g597(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n795_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n786_), .B1(new_n798_), .B2(new_n799_), .ZN(new_n800_));
  INV_X1    g599(.A(new_n556_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n559_), .A2(new_n561_), .A3(new_n801_), .ZN(new_n802_));
  OAI211_X1 g601(.A(new_n802_), .B(new_n566_), .C1(new_n555_), .C2(new_n801_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n567_), .A2(new_n803_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n804_), .B1(new_n538_), .B2(new_n534_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n598_), .B1(new_n800_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT57), .ZN(new_n807_));
  NAND2_X1  g606(.A1(new_n806_), .A2(new_n807_), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n804_), .A2(new_n535_), .ZN(new_n809_));
  AND3_X1   g608(.A1(new_n794_), .A2(KEYINPUT56), .A3(new_n795_), .ZN(new_n810_));
  AOI21_X1  g609(.A(KEYINPUT56), .B1(new_n794_), .B2(new_n795_), .ZN(new_n811_));
  OAI21_X1  g610(.A(new_n809_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT58), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n683_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT58), .B(new_n809_), .C1(new_n810_), .C2(new_n811_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  OAI211_X1 g615(.A(KEYINPUT57), .B(new_n598_), .C1(new_n800_), .C2(new_n805_), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n808_), .A2(new_n816_), .A3(new_n817_), .ZN(new_n818_));
  AOI21_X1  g617(.A(new_n785_), .B1(new_n818_), .B2(new_n614_), .ZN(new_n819_));
  NOR2_X1   g618(.A1(new_n819_), .A2(new_n726_), .ZN(new_n820_));
  NOR2_X1   g619(.A1(new_n266_), .A2(new_n392_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n823_), .A2(new_n205_), .A3(new_n569_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT59), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(new_n826_));
  NAND3_X1  g625(.A1(new_n820_), .A2(KEYINPUT59), .A3(new_n821_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n752_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n824_), .B1(new_n828_), .B2(new_n205_), .ZN(G1340gat));
  OAI21_X1  g628(.A(new_n203_), .B1(new_n541_), .B2(KEYINPUT60), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n823_), .B(new_n830_), .C1(KEYINPUT60), .C2(new_n203_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n541_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n831_), .B1(new_n832_), .B2(new_n203_), .ZN(G1341gat));
  INV_X1    g632(.A(G127gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n823_), .A2(new_n834_), .A3(new_n666_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n614_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n834_), .ZN(G1342gat));
  INV_X1    g636(.A(G134gat), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(new_n822_), .B2(new_n598_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT117), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n839_), .A2(new_n840_), .ZN(new_n841_));
  OAI211_X1 g640(.A(KEYINPUT117), .B(new_n838_), .C1(new_n822_), .C2(new_n598_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n826_), .A2(new_n827_), .ZN(new_n843_));
  NOR2_X1   g642(.A1(new_n683_), .A2(new_n838_), .ZN(new_n844_));
  AOI22_X1  g643(.A1(new_n841_), .A2(new_n842_), .B1(new_n843_), .B2(new_n844_), .ZN(G1343gat));
  NOR3_X1   g644(.A1(new_n655_), .A2(new_n334_), .A3(new_n391_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n820_), .A2(new_n569_), .A3(new_n846_), .ZN(new_n847_));
  XNOR2_X1  g646(.A(new_n847_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g647(.A1(new_n820_), .A2(new_n751_), .A3(new_n846_), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n849_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g649(.A1(new_n820_), .A2(new_n846_), .ZN(new_n851_));
  NOR2_X1   g650(.A1(new_n851_), .A2(new_n614_), .ZN(new_n852_));
  XOR2_X1   g651(.A(KEYINPUT61), .B(G155gat), .Z(new_n853_));
  XNOR2_X1  g652(.A(new_n852_), .B(new_n853_), .ZN(G1346gat));
  OAI21_X1  g653(.A(G162gat), .B1(new_n851_), .B2(new_n683_), .ZN(new_n855_));
  OR2_X1    g654(.A1(new_n598_), .A2(G162gat), .ZN(new_n856_));
  OAI21_X1  g655(.A(new_n855_), .B1(new_n851_), .B2(new_n856_), .ZN(G1347gat));
  NAND3_X1  g656(.A1(new_n655_), .A2(new_n726_), .A3(new_n334_), .ZN(new_n858_));
  NOR3_X1   g657(.A1(new_n819_), .A2(new_n661_), .A3(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n220_), .B1(new_n859_), .B2(new_n569_), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n860_), .A2(KEYINPUT118), .A3(KEYINPUT62), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n569_), .A2(new_n278_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(KEYINPUT119), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n859_), .A2(new_n863_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT118), .B(KEYINPUT62), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n861_), .B(new_n864_), .C1(new_n860_), .C2(new_n865_), .ZN(G1348gat));
  INV_X1    g665(.A(new_n819_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(new_n391_), .ZN(new_n868_));
  NOR4_X1   g667(.A1(new_n868_), .A2(new_n221_), .A3(new_n541_), .A4(new_n858_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n859_), .A2(new_n751_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n221_), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n871_), .A2(KEYINPUT120), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n873_), .A3(new_n221_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n869_), .B1(new_n872_), .B2(new_n874_), .ZN(G1349gat));
  OR3_X1    g674(.A1(new_n868_), .A2(new_n614_), .A3(new_n858_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n614_), .B1(new_n267_), .B2(new_n271_), .ZN(new_n877_));
  AOI22_X1  g676(.A1(new_n876_), .A2(new_n217_), .B1(new_n859_), .B2(new_n877_), .ZN(G1350gat));
  NAND3_X1  g677(.A1(new_n859_), .A2(new_n625_), .A3(new_n213_), .ZN(new_n879_));
  AND2_X1   g678(.A1(new_n859_), .A2(new_n599_), .ZN(new_n880_));
  OAI21_X1  g679(.A(new_n879_), .B1(new_n880_), .B2(new_n249_), .ZN(G1351gat));
  NAND2_X1  g680(.A1(new_n266_), .A2(new_n675_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n883_), .A2(KEYINPUT121), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(KEYINPUT121), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n884_), .A2(new_n334_), .A3(new_n885_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n818_), .A2(new_n614_), .ZN(new_n887_));
  INV_X1    g686(.A(new_n785_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n887_), .B2(new_n888_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n889_), .A2(new_n569_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(new_n890_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n751_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g692(.A(new_n889_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n666_), .A2(new_n895_), .ZN(new_n896_));
  XOR2_X1   g695(.A(new_n896_), .B(KEYINPUT122), .Z(new_n897_));
  NOR2_X1   g696(.A1(new_n894_), .A2(new_n897_), .ZN(new_n898_));
  NOR2_X1   g697(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT124), .B1(new_n898_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902_));
  OAI211_X1 g701(.A(new_n902_), .B(new_n899_), .C1(new_n894_), .C2(new_n897_), .ZN(new_n903_));
  INV_X1    g702(.A(new_n897_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n889_), .A2(new_n900_), .A3(new_n904_), .ZN(new_n905_));
  INV_X1    g704(.A(KEYINPUT123), .ZN(new_n906_));
  OR2_X1    g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n905_), .A2(new_n906_), .ZN(new_n908_));
  AOI22_X1  g707(.A1(new_n901_), .A2(new_n903_), .B1(new_n907_), .B2(new_n908_), .ZN(G1354gat));
  INV_X1    g708(.A(KEYINPUT127), .ZN(new_n910_));
  XNOR2_X1  g709(.A(KEYINPUT126), .B(G218gat), .ZN(new_n911_));
  INV_X1    g710(.A(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(new_n886_), .ZN(new_n913_));
  AOI22_X1  g712(.A1(new_n807_), .A2(new_n806_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n914_));
  AOI21_X1  g713(.A(new_n666_), .B1(new_n914_), .B2(new_n817_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n625_), .B(new_n913_), .C1(new_n915_), .C2(new_n785_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(KEYINPUT125), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n918_));
  NAND3_X1  g717(.A1(new_n889_), .A2(new_n918_), .A3(new_n625_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n912_), .B1(new_n917_), .B2(new_n919_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n889_), .A2(new_n599_), .A3(new_n912_), .ZN(new_n921_));
  INV_X1    g720(.A(new_n921_), .ZN(new_n922_));
  OAI21_X1  g721(.A(new_n910_), .B1(new_n920_), .B2(new_n922_), .ZN(new_n923_));
  AOI21_X1  g722(.A(new_n918_), .B1(new_n889_), .B2(new_n625_), .ZN(new_n924_));
  NOR4_X1   g723(.A1(new_n819_), .A2(KEYINPUT125), .A3(new_n598_), .A4(new_n886_), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n911_), .B1(new_n924_), .B2(new_n925_), .ZN(new_n926_));
  NAND3_X1  g725(.A1(new_n926_), .A2(KEYINPUT127), .A3(new_n921_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n923_), .A2(new_n927_), .ZN(G1355gat));
endmodule


