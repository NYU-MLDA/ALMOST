//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 1 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n643_, new_n644_, new_n645_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n690_, new_n691_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n704_, new_n705_, new_n706_, new_n707_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n727_, new_n728_, new_n729_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n839_, new_n840_, new_n841_, new_n843_, new_n844_, new_n845_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n850_, new_n851_,
    new_n852_, new_n853_, new_n855_, new_n856_, new_n857_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n883_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n897_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_;
  INV_X1    g000(.A(KEYINPUT22), .ZN(new_n202_));
  OAI21_X1  g001(.A(G169gat), .B1(new_n202_), .B2(KEYINPUT78), .ZN(new_n203_));
  INV_X1    g002(.A(KEYINPUT78), .ZN(new_n204_));
  INV_X1    g003(.A(G169gat), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(new_n205_), .A3(KEYINPUT22), .ZN(new_n206_));
  INV_X1    g005(.A(G176gat), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n203_), .A2(new_n206_), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n208_), .A2(KEYINPUT79), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT79), .ZN(new_n211_));
  NAND4_X1  g010(.A1(new_n203_), .A2(new_n206_), .A3(new_n211_), .A4(new_n207_), .ZN(new_n212_));
  AOI21_X1  g011(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  NAND3_X1  g013(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n215_));
  INV_X1    g014(.A(G183gat), .ZN(new_n216_));
  INV_X1    g015(.A(G190gat), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n216_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n214_), .A2(new_n215_), .A3(new_n218_), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n209_), .A2(new_n210_), .A3(new_n212_), .A4(new_n219_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n221_));
  OAI21_X1  g020(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n222_));
  INV_X1    g021(.A(new_n222_), .ZN(new_n223_));
  AOI21_X1  g022(.A(new_n221_), .B1(new_n223_), .B2(new_n210_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n215_), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n225_), .A2(new_n213_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT25), .B(G183gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n217_), .A2(KEYINPUT26), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n227_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n232_), .A2(G190gat), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n229_), .B1(new_n228_), .B2(new_n233_), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n224_), .B(new_n226_), .C1(new_n231_), .C2(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n220_), .A2(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT80), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT80), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n220_), .A2(new_n238_), .A3(new_n235_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n237_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G227gat), .A2(G233gat), .ZN(new_n241_));
  INV_X1    g040(.A(G15gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(new_n241_), .B(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n243_), .B(KEYINPUT30), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n240_), .B(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G127gat), .B(G134gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G113gat), .B(G120gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT81), .ZN(new_n249_));
  XNOR2_X1  g048(.A(new_n248_), .B(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n245_), .B(new_n250_), .ZN(new_n251_));
  XOR2_X1   g050(.A(G71gat), .B(G99gat), .Z(new_n252_));
  XNOR2_X1  g051(.A(new_n252_), .B(G43gat), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n253_), .B(KEYINPUT31), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  OR2_X1    g054(.A1(new_n251_), .A2(new_n255_), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n251_), .A2(new_n255_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(G197gat), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n260_), .A2(G204gat), .ZN(new_n261_));
  INV_X1    g060(.A(G204gat), .ZN(new_n262_));
  OAI21_X1  g061(.A(KEYINPUT86), .B1(new_n262_), .B2(G197gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT86), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(new_n260_), .A3(G204gat), .ZN(new_n265_));
  AOI21_X1  g064(.A(new_n261_), .B1(new_n263_), .B2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT21), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G211gat), .B(G218gat), .ZN(new_n268_));
  NOR3_X1   g067(.A1(new_n266_), .A2(new_n267_), .A3(new_n268_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n262_), .A2(G197gat), .ZN(new_n270_));
  AOI21_X1  g069(.A(new_n264_), .B1(new_n260_), .B2(G204gat), .ZN(new_n271_));
  NOR3_X1   g070(.A1(new_n262_), .A2(KEYINPUT86), .A3(G197gat), .ZN(new_n272_));
  OAI211_X1 g071(.A(new_n267_), .B(new_n270_), .C1(new_n271_), .C2(new_n272_), .ZN(new_n273_));
  INV_X1    g072(.A(KEYINPUT87), .ZN(new_n274_));
  NAND2_X1  g073(.A1(new_n273_), .A2(new_n274_), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n266_), .A2(KEYINPUT87), .A3(new_n267_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n275_), .A2(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n268_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n270_), .A2(KEYINPUT85), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT85), .ZN(new_n280_));
  NAND3_X1  g079(.A1(new_n280_), .A2(new_n262_), .A3(G197gat), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n260_), .A2(G204gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n279_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n278_), .B1(new_n283_), .B2(KEYINPUT21), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n269_), .B1(new_n277_), .B2(new_n284_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT29), .ZN(new_n286_));
  OR3_X1    g085(.A1(KEYINPUT82), .A2(G155gat), .A3(G162gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT1), .ZN(new_n289_));
  INV_X1    g088(.A(KEYINPUT1), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n290_), .A2(G155gat), .A3(G162gat), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n287_), .A2(new_n289_), .A3(new_n291_), .A4(new_n292_), .ZN(new_n293_));
  INV_X1    g092(.A(G141gat), .ZN(new_n294_));
  INV_X1    g093(.A(G148gat), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(G141gat), .A2(G148gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n296_), .A3(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT3), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n299_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT2), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n297_), .A2(new_n301_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n303_));
  OAI21_X1  g102(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n304_));
  NAND4_X1  g103(.A1(new_n300_), .A2(new_n302_), .A3(new_n303_), .A4(new_n304_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n305_), .A2(new_n287_), .A3(new_n292_), .A4(new_n288_), .ZN(new_n306_));
  AOI21_X1  g105(.A(new_n286_), .B1(new_n298_), .B2(new_n306_), .ZN(new_n307_));
  OAI21_X1  g106(.A(KEYINPUT84), .B1(new_n285_), .B2(new_n307_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n263_), .A2(new_n265_), .ZN(new_n309_));
  AND4_X1   g108(.A1(KEYINPUT87), .A2(new_n309_), .A3(new_n267_), .A4(new_n270_), .ZN(new_n310_));
  AOI21_X1  g109(.A(KEYINPUT87), .B1(new_n266_), .B2(new_n267_), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n284_), .B1(new_n310_), .B2(new_n311_), .ZN(new_n312_));
  INV_X1    g111(.A(new_n269_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT84), .ZN(new_n315_));
  INV_X1    g114(.A(new_n307_), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n314_), .A2(new_n315_), .A3(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n308_), .A2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(G228gat), .ZN(new_n319_));
  INV_X1    g118(.A(G233gat), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n318_), .A2(new_n322_), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n308_), .A2(new_n317_), .A3(G228gat), .A4(G233gat), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  AND2_X1   g124(.A1(new_n298_), .A2(new_n306_), .ZN(new_n326_));
  XOR2_X1   g125(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n326_), .A2(new_n286_), .A3(new_n328_), .ZN(new_n329_));
  XOR2_X1   g128(.A(G22gat), .B(G50gat), .Z(new_n330_));
  NAND2_X1  g129(.A1(new_n298_), .A2(new_n306_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n327_), .B1(new_n331_), .B2(KEYINPUT29), .ZN(new_n332_));
  AND3_X1   g131(.A1(new_n329_), .A2(new_n330_), .A3(new_n332_), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n330_), .B1(new_n329_), .B2(new_n332_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(G78gat), .B(G106gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n335_), .A2(new_n336_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n325_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n338_), .ZN(new_n339_));
  XNOR2_X1  g138(.A(new_n336_), .B(KEYINPUT88), .ZN(new_n340_));
  INV_X1    g139(.A(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n341_), .B1(new_n323_), .B2(new_n324_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(new_n323_), .A2(new_n324_), .A3(new_n341_), .ZN(new_n343_));
  INV_X1    g142(.A(KEYINPUT89), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n335_), .A2(new_n344_), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n342_), .B1(new_n343_), .B2(new_n345_), .ZN(new_n346_));
  AND3_X1   g145(.A1(new_n345_), .A2(new_n325_), .A3(new_n340_), .ZN(new_n347_));
  OAI21_X1  g146(.A(new_n339_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n250_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT93), .B(KEYINPUT4), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n350_), .A2(new_n331_), .A3(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n326_), .A2(new_n248_), .ZN(new_n353_));
  OAI211_X1 g152(.A(KEYINPUT4), .B(new_n353_), .C1(new_n250_), .C2(new_n326_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G225gat), .A2(G233gat), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n352_), .A2(new_n354_), .A3(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(G1gat), .B(G29gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n357_), .B(G85gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT0), .B(G57gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n358_), .B(new_n359_), .Z(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n350_), .A2(new_n331_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n355_), .ZN(new_n363_));
  NAND3_X1  g162(.A1(new_n362_), .A2(new_n353_), .A3(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n356_), .A2(new_n361_), .A3(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n352_), .A2(new_n354_), .A3(new_n363_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n366_), .A2(KEYINPUT94), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT94), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n352_), .A2(new_n354_), .A3(new_n368_), .A4(new_n363_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n362_), .A2(new_n353_), .A3(new_n355_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n367_), .A2(new_n360_), .A3(new_n369_), .A4(new_n370_), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT95), .ZN(new_n372_));
  NOR2_X1   g171(.A1(new_n372_), .A2(KEYINPUT33), .ZN(new_n373_));
  OAI21_X1  g172(.A(new_n365_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n374_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n375_));
  XNOR2_X1  g174(.A(G8gat), .B(G36gat), .ZN(new_n376_));
  XNOR2_X1  g175(.A(new_n376_), .B(KEYINPUT18), .ZN(new_n377_));
  XNOR2_X1  g176(.A(G64gat), .B(G92gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n377_), .B(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT92), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n216_), .A2(KEYINPUT25), .ZN(new_n382_));
  INV_X1    g181(.A(KEYINPUT25), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(G183gat), .ZN(new_n384_));
  NAND4_X1  g183(.A1(new_n228_), .A2(new_n233_), .A3(new_n382_), .A4(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n224_), .A2(new_n226_), .A3(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(KEYINPUT22), .B(G169gat), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(new_n207_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n388_), .A2(new_n219_), .A3(new_n210_), .ZN(new_n389_));
  AND2_X1   g188(.A1(new_n386_), .A2(new_n389_), .ZN(new_n390_));
  AOI21_X1  g189(.A(KEYINPUT91), .B1(new_n285_), .B2(new_n390_), .ZN(new_n391_));
  AND4_X1   g190(.A1(KEYINPUT91), .A2(new_n312_), .A3(new_n313_), .A4(new_n390_), .ZN(new_n392_));
  NOR2_X1   g191(.A1(new_n391_), .A2(new_n392_), .ZN(new_n393_));
  AND3_X1   g192(.A1(new_n220_), .A2(new_n238_), .A3(new_n235_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n238_), .B1(new_n220_), .B2(new_n235_), .ZN(new_n395_));
  OAI21_X1  g194(.A(new_n314_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n397_), .B(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT20), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n396_), .A2(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n381_), .B1(new_n393_), .B2(new_n402_), .ZN(new_n403_));
  INV_X1    g202(.A(new_n401_), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n404_), .B1(new_n240_), .B2(new_n314_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n312_), .A2(new_n313_), .A3(new_n390_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT91), .ZN(new_n407_));
  NAND2_X1  g206(.A1(new_n406_), .A2(new_n407_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n285_), .A2(KEYINPUT91), .A3(new_n390_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n405_), .A2(KEYINPUT92), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n403_), .A2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(new_n399_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n390_), .ZN(new_n414_));
  AOI21_X1  g213(.A(new_n400_), .B1(new_n314_), .B2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n237_), .A2(new_n285_), .A3(new_n239_), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n413_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n380_), .B1(new_n412_), .B2(new_n418_), .ZN(new_n419_));
  AOI211_X1 g218(.A(new_n379_), .B(new_n417_), .C1(new_n403_), .C2(new_n411_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n375_), .A2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n367_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n423_), .A2(new_n361_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n424_), .A2(new_n371_), .ZN(new_n425_));
  XOR2_X1   g224(.A(KEYINPUT96), .B(KEYINPUT20), .Z(new_n426_));
  XNOR2_X1  g225(.A(new_n390_), .B(KEYINPUT97), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n426_), .B1(new_n427_), .B2(new_n314_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n396_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n399_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n415_), .A2(new_n416_), .A3(new_n413_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AND2_X1   g231(.A1(new_n380_), .A2(KEYINPUT32), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n412_), .A2(new_n418_), .ZN(new_n435_));
  OAI211_X1 g234(.A(new_n425_), .B(new_n434_), .C1(new_n433_), .C2(new_n435_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n349_), .B1(new_n422_), .B2(new_n436_), .ZN(new_n437_));
  NOR3_X1   g236(.A1(new_n393_), .A2(new_n402_), .A3(new_n381_), .ZN(new_n438_));
  AOI21_X1  g237(.A(KEYINPUT92), .B1(new_n405_), .B2(new_n410_), .ZN(new_n439_));
  OAI211_X1 g238(.A(new_n380_), .B(new_n418_), .C1(new_n438_), .C2(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT98), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n440_), .A2(new_n441_), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n412_), .A2(KEYINPUT98), .A3(new_n380_), .A4(new_n418_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT27), .ZN(new_n444_));
  AOI21_X1  g243(.A(new_n444_), .B1(new_n432_), .B2(new_n379_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n442_), .A2(new_n443_), .A3(new_n445_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n444_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NOR3_X1   g247(.A1(new_n448_), .A2(new_n348_), .A3(new_n425_), .ZN(new_n449_));
  OAI21_X1  g248(.A(new_n259_), .B1(new_n437_), .B2(new_n449_), .ZN(new_n450_));
  NAND3_X1  g249(.A1(new_n446_), .A2(new_n447_), .A3(new_n348_), .ZN(new_n451_));
  INV_X1    g250(.A(KEYINPUT99), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n446_), .A2(new_n447_), .A3(new_n348_), .A4(KEYINPUT99), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(new_n425_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n258_), .A2(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(new_n457_), .ZN(new_n458_));
  AOI21_X1  g257(.A(KEYINPUT100), .B1(new_n455_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT100), .ZN(new_n460_));
  AOI211_X1 g259(.A(new_n460_), .B(new_n457_), .C1(new_n453_), .C2(new_n454_), .ZN(new_n461_));
  OAI21_X1  g260(.A(new_n450_), .B1(new_n459_), .B2(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G29gat), .B(G36gat), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G43gat), .B(G50gat), .ZN(new_n464_));
  OR2_X1    g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n463_), .A2(new_n464_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n465_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n467_), .B(KEYINPUT74), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G15gat), .B(G22gat), .ZN(new_n469_));
  INV_X1    g268(.A(G1gat), .ZN(new_n470_));
  INV_X1    g269(.A(G8gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT14), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n469_), .A2(new_n472_), .ZN(new_n473_));
  XNOR2_X1  g272(.A(G1gat), .B(G8gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(new_n473_), .B(new_n474_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n468_), .A2(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n467_), .B(KEYINPUT15), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(new_n475_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G229gat), .A2(G233gat), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n477_), .A2(new_n479_), .A3(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(KEYINPUT74), .ZN(new_n482_));
  XNOR2_X1  g281(.A(new_n467_), .B(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(new_n475_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n477_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n480_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  AND2_X1   g286(.A1(new_n487_), .A2(KEYINPUT75), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n487_), .A2(KEYINPUT75), .ZN(new_n489_));
  OAI21_X1  g288(.A(new_n481_), .B1(new_n488_), .B2(new_n489_), .ZN(new_n490_));
  XNOR2_X1  g289(.A(G113gat), .B(G141gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(G169gat), .B(G197gat), .ZN(new_n492_));
  XOR2_X1   g291(.A(new_n491_), .B(new_n492_), .Z(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n490_), .A2(new_n494_), .ZN(new_n495_));
  OAI211_X1 g294(.A(new_n481_), .B(new_n493_), .C1(new_n488_), .C2(new_n489_), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n495_), .A2(KEYINPUT76), .A3(new_n496_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT76), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n490_), .A2(new_n498_), .A3(new_n494_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n497_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(new_n500_), .ZN(new_n501_));
  AND2_X1   g300(.A1(new_n462_), .A2(new_n501_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G230gat), .A2(G233gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(G99gat), .A2(G106gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n504_), .B(KEYINPUT6), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT64), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(G85gat), .ZN(new_n508_));
  INV_X1    g307(.A(G92gat), .ZN(new_n509_));
  NOR3_X1   g308(.A1(new_n508_), .A2(new_n509_), .A3(KEYINPUT9), .ZN(new_n510_));
  XOR2_X1   g309(.A(G85gat), .B(G92gat), .Z(new_n511_));
  AOI21_X1  g310(.A(new_n510_), .B1(new_n511_), .B2(KEYINPUT9), .ZN(new_n512_));
  XNOR2_X1  g311(.A(KEYINPUT10), .B(G99gat), .ZN(new_n513_));
  OAI211_X1 g312(.A(new_n507_), .B(new_n512_), .C1(G106gat), .C2(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT8), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  NOR3_X1   g315(.A1(KEYINPUT65), .A2(G99gat), .A3(G106gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n517_), .B(KEYINPUT7), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n516_), .B1(new_n507_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n505_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n515_), .B1(new_n520_), .B2(new_n511_), .ZN(new_n521_));
  OAI21_X1  g320(.A(new_n514_), .B1(new_n519_), .B2(new_n521_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(G57gat), .B(G64gat), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G71gat), .B(G78gat), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n523_), .A2(new_n524_), .A3(KEYINPUT11), .ZN(new_n525_));
  AND2_X1   g324(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n526_));
  OR2_X1    g325(.A1(new_n526_), .A2(new_n524_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n523_), .A2(KEYINPUT11), .ZN(new_n528_));
  OAI21_X1  g327(.A(new_n525_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n522_), .A2(new_n530_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n514_), .B(new_n529_), .C1(new_n519_), .C2(new_n521_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n503_), .B1(new_n531_), .B2(new_n532_), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT66), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n503_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT67), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT67), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n532_), .A2(new_n537_), .A3(new_n503_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n536_), .A2(new_n538_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT12), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n540_), .B1(new_n522_), .B2(new_n530_), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n522_), .A2(new_n540_), .A3(new_n530_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n542_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n539_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n544_));
  AND2_X1   g343(.A1(new_n534_), .A2(new_n544_), .ZN(new_n545_));
  XNOR2_X1  g344(.A(G120gat), .B(G148gat), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n546_), .B(KEYINPUT5), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G176gat), .B(G204gat), .ZN(new_n548_));
  XOR2_X1   g347(.A(new_n547_), .B(new_n548_), .Z(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n545_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT13), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n545_), .A2(new_n550_), .ZN(new_n554_));
  OR3_X1    g353(.A1(new_n552_), .A2(new_n553_), .A3(new_n554_), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n553_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n555_), .A2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(G183gat), .B(G211gat), .ZN(new_n559_));
  XNOR2_X1  g358(.A(new_n559_), .B(KEYINPUT72), .ZN(new_n560_));
  XOR2_X1   g359(.A(KEYINPUT71), .B(KEYINPUT16), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  XNOR2_X1  g361(.A(G127gat), .B(G155gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n562_), .B(new_n563_), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n564_), .A2(KEYINPUT17), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n564_), .A2(KEYINPUT17), .ZN(new_n566_));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567_));
  XNOR2_X1  g366(.A(new_n475_), .B(new_n567_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(new_n529_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n565_), .A2(new_n566_), .A3(new_n569_), .ZN(new_n570_));
  OR2_X1    g369(.A1(new_n569_), .A2(new_n566_), .ZN(new_n571_));
  AND2_X1   g370(.A1(new_n570_), .A2(new_n571_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT73), .ZN(new_n573_));
  XNOR2_X1  g372(.A(KEYINPUT70), .B(KEYINPUT37), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(new_n467_), .ZN(new_n576_));
  XNOR2_X1  g375(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n577_));
  NAND2_X1  g376(.A1(G232gat), .A2(G233gat), .ZN(new_n578_));
  XNOR2_X1  g377(.A(new_n577_), .B(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  OAI22_X1  g379(.A1(new_n522_), .A2(new_n576_), .B1(KEYINPUT35), .B2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n581_), .B1(new_n478_), .B2(new_n522_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(KEYINPUT35), .ZN(new_n583_));
  OR2_X1    g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n582_), .A2(new_n583_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  XNOR2_X1  g385(.A(G190gat), .B(G218gat), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n587_), .B(KEYINPUT69), .ZN(new_n588_));
  XOR2_X1   g387(.A(G134gat), .B(G162gat), .Z(new_n589_));
  XNOR2_X1  g388(.A(new_n588_), .B(new_n589_), .ZN(new_n590_));
  XNOR2_X1  g389(.A(new_n590_), .B(KEYINPUT36), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n586_), .A2(new_n591_), .ZN(new_n592_));
  INV_X1    g391(.A(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n590_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n594_), .A2(KEYINPUT36), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n584_), .A2(new_n595_), .A3(new_n585_), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  OAI21_X1  g396(.A(new_n575_), .B1(new_n593_), .B2(new_n597_), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n592_), .A2(new_n596_), .A3(new_n574_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n598_), .A2(new_n599_), .ZN(new_n600_));
  AND4_X1   g399(.A1(new_n502_), .A2(new_n558_), .A3(new_n573_), .A4(new_n600_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n601_), .A2(new_n470_), .A3(new_n425_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT38), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n602_), .A2(new_n603_), .ZN(new_n604_));
  OR3_X1    g403(.A1(new_n593_), .A2(KEYINPUT101), .A3(new_n597_), .ZN(new_n605_));
  OAI21_X1  g404(.A(KEYINPUT101), .B1(new_n593_), .B2(new_n597_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n607_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n462_), .A2(new_n608_), .ZN(new_n609_));
  INV_X1    g408(.A(new_n572_), .ZN(new_n610_));
  NOR3_X1   g409(.A1(new_n557_), .A2(new_n500_), .A3(new_n610_), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  OAI21_X1  g411(.A(G1gat), .B1(new_n612_), .B2(new_n456_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n602_), .A2(new_n603_), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n604_), .A2(new_n613_), .A3(new_n614_), .ZN(G1324gat));
  NAND3_X1  g414(.A1(new_n601_), .A2(new_n471_), .A3(new_n448_), .ZN(new_n616_));
  AND2_X1   g415(.A1(new_n609_), .A2(new_n611_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n617_), .A2(new_n448_), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n618_), .A2(G8gat), .ZN(new_n619_));
  AND2_X1   g418(.A1(new_n619_), .A2(KEYINPUT39), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n619_), .A2(KEYINPUT39), .ZN(new_n621_));
  OAI21_X1  g420(.A(new_n616_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(G1325gat));
  INV_X1    g423(.A(KEYINPUT41), .ZN(new_n625_));
  OAI21_X1  g424(.A(G15gat), .B1(new_n612_), .B2(new_n259_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n626_), .A2(KEYINPUT102), .ZN(new_n627_));
  INV_X1    g426(.A(new_n627_), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n626_), .A2(KEYINPUT102), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n625_), .B1(new_n628_), .B2(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n629_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n631_), .A2(KEYINPUT41), .A3(new_n627_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n601_), .A2(new_n242_), .A3(new_n258_), .ZN(new_n633_));
  NAND3_X1  g432(.A1(new_n630_), .A2(new_n632_), .A3(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n634_), .A2(KEYINPUT103), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n636_));
  NAND4_X1  g435(.A1(new_n630_), .A2(new_n632_), .A3(new_n636_), .A4(new_n633_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n635_), .A2(new_n637_), .ZN(G1326gat));
  INV_X1    g437(.A(G22gat), .ZN(new_n639_));
  XNOR2_X1  g438(.A(new_n348_), .B(KEYINPUT104), .ZN(new_n640_));
  AOI21_X1  g439(.A(new_n639_), .B1(new_n617_), .B2(new_n640_), .ZN(new_n641_));
  XOR2_X1   g440(.A(new_n641_), .B(KEYINPUT42), .Z(new_n642_));
  NAND2_X1  g441(.A1(new_n640_), .A2(new_n639_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT105), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n601_), .A2(new_n644_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n642_), .A2(new_n645_), .ZN(G1327gat));
  INV_X1    g445(.A(new_n573_), .ZN(new_n647_));
  AND4_X1   g446(.A1(new_n502_), .A2(new_n558_), .A3(new_n647_), .A4(new_n607_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n456_), .A2(G29gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT107), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n648_), .A2(new_n650_), .ZN(new_n651_));
  NOR3_X1   g450(.A1(new_n557_), .A2(new_n500_), .A3(new_n573_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT43), .ZN(new_n653_));
  INV_X1    g452(.A(new_n600_), .ZN(new_n654_));
  AND3_X1   g453(.A1(new_n462_), .A2(new_n653_), .A3(new_n654_), .ZN(new_n655_));
  AOI21_X1  g454(.A(new_n653_), .B1(new_n462_), .B2(new_n654_), .ZN(new_n656_));
  OAI21_X1  g455(.A(new_n652_), .B1(new_n655_), .B2(new_n656_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n657_), .A2(new_n658_), .ZN(new_n659_));
  OAI211_X1 g458(.A(KEYINPUT44), .B(new_n652_), .C1(new_n655_), .C2(new_n656_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n659_), .A2(new_n425_), .A3(new_n660_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT106), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n661_), .A2(new_n662_), .A3(G29gat), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n662_), .B1(new_n661_), .B2(G29gat), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n651_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT108), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT108), .ZN(new_n667_));
  OAI211_X1 g466(.A(new_n667_), .B(new_n651_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n666_), .A2(new_n668_), .ZN(G1328gat));
  NAND3_X1  g468(.A1(new_n659_), .A2(new_n448_), .A3(new_n660_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT109), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT109), .ZN(new_n672_));
  NAND4_X1  g471(.A1(new_n659_), .A2(new_n672_), .A3(new_n448_), .A4(new_n660_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n671_), .A2(G36gat), .A3(new_n673_), .ZN(new_n674_));
  INV_X1    g473(.A(G36gat), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n648_), .A2(new_n675_), .A3(new_n448_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT45), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n674_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT46), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n678_), .A2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n674_), .A2(KEYINPUT46), .A3(new_n677_), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n680_), .A2(new_n681_), .ZN(G1329gat));
  AND2_X1   g481(.A1(new_n659_), .A2(new_n660_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n683_), .A2(G43gat), .A3(new_n258_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n648_), .A2(new_n258_), .ZN(new_n685_));
  XNOR2_X1  g484(.A(KEYINPUT110), .B(G43gat), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n685_), .A2(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n684_), .A2(new_n687_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g488(.A(G50gat), .B1(new_n648_), .B2(new_n640_), .ZN(new_n690_));
  AND2_X1   g489(.A1(new_n349_), .A2(G50gat), .ZN(new_n691_));
  AOI21_X1  g490(.A(new_n690_), .B1(new_n683_), .B2(new_n691_), .ZN(G1331gat));
  NOR2_X1   g491(.A1(new_n501_), .A2(new_n647_), .ZN(new_n693_));
  INV_X1    g492(.A(new_n693_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n558_), .A2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n609_), .A2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(new_n696_), .ZN(new_n697_));
  OAI21_X1  g496(.A(G57gat), .B1(new_n697_), .B2(new_n456_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n462_), .A2(new_n500_), .ZN(new_n699_));
  NOR4_X1   g498(.A1(new_n699_), .A2(new_n558_), .A3(new_n647_), .A4(new_n654_), .ZN(new_n700_));
  INV_X1    g499(.A(G57gat), .ZN(new_n701_));
  NAND3_X1  g500(.A1(new_n700_), .A2(new_n701_), .A3(new_n425_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n698_), .A2(new_n702_), .ZN(G1332gat));
  INV_X1    g502(.A(G64gat), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n704_), .B1(new_n696_), .B2(new_n448_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT48), .Z(new_n706_));
  NAND3_X1  g505(.A1(new_n700_), .A2(new_n704_), .A3(new_n448_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(G1333gat));
  INV_X1    g507(.A(G71gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(new_n709_), .B1(new_n696_), .B2(new_n258_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(KEYINPUT111), .B(KEYINPUT49), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n710_), .B(new_n711_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n700_), .A2(new_n709_), .A3(new_n258_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1334gat));
  INV_X1    g513(.A(G78gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n715_), .B1(new_n696_), .B2(new_n640_), .ZN(new_n716_));
  XOR2_X1   g515(.A(new_n716_), .B(KEYINPUT50), .Z(new_n717_));
  NAND3_X1  g516(.A1(new_n700_), .A2(new_n715_), .A3(new_n640_), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n717_), .A2(new_n718_), .ZN(G1335gat));
  NAND3_X1  g518(.A1(new_n557_), .A2(new_n647_), .A3(new_n607_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n699_), .A2(new_n720_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n721_), .A2(new_n508_), .A3(new_n425_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n655_), .A2(new_n656_), .ZN(new_n723_));
  NOR4_X1   g522(.A1(new_n723_), .A2(new_n501_), .A3(new_n558_), .A4(new_n573_), .ZN(new_n724_));
  AND2_X1   g523(.A1(new_n724_), .A2(new_n425_), .ZN(new_n725_));
  OAI21_X1  g524(.A(new_n722_), .B1(new_n725_), .B2(new_n508_), .ZN(G1336gat));
  AND3_X1   g525(.A1(new_n721_), .A2(new_n509_), .A3(new_n448_), .ZN(new_n727_));
  NAND2_X1  g526(.A1(new_n724_), .A2(new_n448_), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n727_), .B1(new_n728_), .B2(G92gat), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT112), .ZN(G1337gat));
  NAND2_X1  g529(.A1(new_n724_), .A2(new_n258_), .ZN(new_n731_));
  INV_X1    g530(.A(new_n513_), .ZN(new_n732_));
  NAND3_X1  g531(.A1(new_n721_), .A2(new_n258_), .A3(new_n732_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n733_), .A2(KEYINPUT113), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n733_), .A2(KEYINPUT113), .ZN(new_n735_));
  AOI22_X1  g534(.A1(new_n731_), .A2(G99gat), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT51), .ZN(new_n737_));
  XNOR2_X1  g536(.A(new_n736_), .B(new_n737_), .ZN(G1338gat));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n724_), .A2(new_n349_), .ZN(new_n740_));
  INV_X1    g539(.A(G106gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n739_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n741_), .B1(new_n724_), .B2(new_n349_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(KEYINPUT52), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n721_), .A2(new_n741_), .A3(new_n349_), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n746_), .B(KEYINPUT114), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n742_), .A2(new_n743_), .A3(new_n745_), .A4(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n744_), .B2(KEYINPUT52), .ZN(new_n749_));
  AOI211_X1 g548(.A(new_n739_), .B(new_n741_), .C1(new_n724_), .C2(new_n349_), .ZN(new_n750_));
  OAI21_X1  g549(.A(KEYINPUT53), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n748_), .A2(new_n751_), .ZN(G1339gat));
  NAND3_X1  g551(.A1(new_n455_), .A2(new_n258_), .A3(new_n425_), .ZN(new_n753_));
  INV_X1    g552(.A(new_n753_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n551_), .A2(new_n497_), .A3(new_n499_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT117), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND4_X1  g556(.A1(new_n551_), .A2(new_n497_), .A3(KEYINPUT117), .A4(new_n499_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT55), .ZN(new_n759_));
  NAND3_X1  g558(.A1(new_n544_), .A2(KEYINPUT118), .A3(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n541_), .ZN(new_n761_));
  AOI22_X1  g560(.A1(new_n536_), .A2(new_n538_), .B1(new_n761_), .B2(new_n542_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT118), .ZN(new_n763_));
  OAI21_X1  g562(.A(KEYINPUT55), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n532_), .B1(new_n543_), .B2(new_n541_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n503_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT119), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT119), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n765_), .A2(new_n769_), .A3(new_n766_), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n760_), .A2(new_n764_), .A3(new_n768_), .A4(new_n770_), .ZN(new_n771_));
  NAND3_X1  g570(.A1(new_n771_), .A2(KEYINPUT56), .A3(new_n549_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(KEYINPUT56), .B1(new_n771_), .B2(new_n549_), .ZN(new_n774_));
  OAI211_X1 g573(.A(new_n757_), .B(new_n758_), .C1(new_n773_), .C2(new_n774_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n496_), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n477_), .A2(new_n479_), .A3(new_n486_), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AOI211_X1 g577(.A(new_n493_), .B(new_n778_), .C1(new_n485_), .C2(new_n480_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n776_), .A2(new_n779_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n780_), .B1(new_n552_), .B2(new_n554_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n775_), .A2(new_n781_), .ZN(new_n782_));
  AOI21_X1  g581(.A(KEYINPUT57), .B1(new_n782_), .B2(new_n608_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n784_));
  AOI211_X1 g583(.A(new_n784_), .B(new_n607_), .C1(new_n775_), .C2(new_n781_), .ZN(new_n785_));
  NOR2_X1   g584(.A1(new_n783_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n551_), .A2(new_n780_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n771_), .A2(new_n549_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT56), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n787_), .B1(new_n790_), .B2(new_n772_), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n654_), .B1(new_n791_), .B2(KEYINPUT58), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT120), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  OAI211_X1 g593(.A(KEYINPUT120), .B(new_n654_), .C1(new_n791_), .C2(KEYINPUT58), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n791_), .A2(KEYINPUT58), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n794_), .A2(new_n795_), .A3(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n572_), .B1(new_n786_), .B2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT115), .B1(new_n557_), .B2(new_n694_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n555_), .A2(new_n693_), .A3(new_n800_), .A4(new_n556_), .ZN(new_n801_));
  NAND3_X1  g600(.A1(new_n799_), .A2(new_n600_), .A3(new_n801_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(KEYINPUT116), .B(KEYINPUT54), .ZN(new_n803_));
  INV_X1    g602(.A(new_n803_), .ZN(new_n804_));
  XNOR2_X1  g603(.A(new_n802_), .B(new_n804_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n754_), .B1(new_n798_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(G113gat), .ZN(new_n808_));
  NAND3_X1  g607(.A1(new_n807_), .A2(new_n808_), .A3(new_n501_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n782_), .A2(new_n608_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n810_), .A2(new_n784_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n782_), .A2(KEYINPUT57), .A3(new_n608_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n797_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n647_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n802_), .B(new_n803_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n815_), .A2(new_n816_), .ZN(new_n817_));
  NOR2_X1   g616(.A1(new_n753_), .A2(KEYINPUT59), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n806_), .A2(KEYINPUT59), .B1(new_n817_), .B2(new_n818_), .ZN(new_n819_));
  AND2_X1   g618(.A1(new_n819_), .A2(new_n501_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n809_), .B1(new_n820_), .B2(new_n808_), .ZN(G1340gat));
  XOR2_X1   g620(.A(KEYINPUT121), .B(G120gat), .Z(new_n822_));
  OAI21_X1  g621(.A(new_n822_), .B1(new_n558_), .B2(KEYINPUT60), .ZN(new_n823_));
  OAI211_X1 g622(.A(new_n807_), .B(new_n823_), .C1(KEYINPUT60), .C2(new_n822_), .ZN(new_n824_));
  AND2_X1   g623(.A1(new_n819_), .A2(new_n557_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n824_), .B1(new_n825_), .B2(new_n822_), .ZN(G1341gat));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n827_));
  INV_X1    g626(.A(G127gat), .ZN(new_n828_));
  AOI21_X1  g627(.A(new_n828_), .B1(new_n819_), .B2(new_n572_), .ZN(new_n829_));
  NOR3_X1   g628(.A1(new_n806_), .A2(G127gat), .A3(new_n647_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n827_), .B1(new_n829_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n806_), .A2(KEYINPUT59), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n817_), .A2(new_n818_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n572_), .A3(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n834_), .A2(G127gat), .ZN(new_n835_));
  INV_X1    g634(.A(new_n830_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n835_), .A2(KEYINPUT122), .A3(new_n836_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n831_), .A2(new_n837_), .ZN(G1342gat));
  AOI21_X1  g637(.A(G134gat), .B1(new_n807_), .B2(new_n607_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n654_), .A2(G134gat), .ZN(new_n840_));
  XNOR2_X1  g639(.A(new_n840_), .B(KEYINPUT123), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n839_), .B1(new_n819_), .B2(new_n841_), .ZN(G1343gat));
  NOR2_X1   g641(.A1(new_n258_), .A2(new_n348_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n610_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n844_), .B1(new_n845_), .B2(new_n816_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n448_), .A2(new_n456_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(KEYINPUT124), .A3(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  AOI21_X1  g648(.A(KEYINPUT124), .B1(new_n846_), .B2(new_n847_), .ZN(new_n850_));
  OAI21_X1  g649(.A(new_n501_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(G141gat), .ZN(new_n852_));
  OAI211_X1 g651(.A(new_n294_), .B(new_n501_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1344gat));
  OAI21_X1  g653(.A(new_n557_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n855_), .A2(G148gat), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n295_), .B(new_n557_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n856_), .A2(new_n857_), .ZN(G1345gat));
  OAI21_X1  g657(.A(new_n573_), .B1(new_n849_), .B2(new_n850_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT61), .B(G155gat), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(new_n861_));
  INV_X1    g660(.A(new_n860_), .ZN(new_n862_));
  OAI211_X1 g661(.A(new_n573_), .B(new_n862_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n861_), .A2(new_n863_), .ZN(G1346gat));
  INV_X1    g663(.A(G162gat), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n865_), .B(new_n607_), .C1(new_n849_), .C2(new_n850_), .ZN(new_n866_));
  INV_X1    g665(.A(new_n850_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n600_), .B1(new_n867_), .B2(new_n848_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n866_), .B1(new_n868_), .B2(new_n865_), .ZN(G1347gat));
  AOI21_X1  g668(.A(new_n425_), .B1(new_n446_), .B2(new_n447_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(new_n258_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n640_), .ZN(new_n872_));
  AND2_X1   g671(.A1(new_n817_), .A2(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n205_), .B1(new_n873_), .B2(new_n501_), .ZN(new_n874_));
  OR2_X1    g673(.A1(new_n874_), .A2(KEYINPUT62), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(KEYINPUT62), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n873_), .A2(new_n387_), .A3(new_n501_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n875_), .A2(new_n876_), .A3(new_n877_), .ZN(G1348gat));
  AOI21_X1  g677(.A(G176gat), .B1(new_n873_), .B2(new_n557_), .ZN(new_n879_));
  AOI21_X1  g678(.A(new_n349_), .B1(new_n845_), .B2(new_n816_), .ZN(new_n880_));
  NOR3_X1   g679(.A1(new_n558_), .A2(new_n207_), .A3(new_n871_), .ZN(new_n881_));
  AOI21_X1  g680(.A(new_n879_), .B1(new_n880_), .B2(new_n881_), .ZN(G1349gat));
  INV_X1    g681(.A(new_n873_), .ZN(new_n883_));
  NOR3_X1   g682(.A1(new_n883_), .A2(new_n227_), .A3(new_n610_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n880_), .A2(new_n258_), .A3(new_n573_), .A4(new_n870_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n216_), .B2(new_n885_), .ZN(G1350gat));
  OAI21_X1  g685(.A(G190gat), .B1(new_n883_), .B2(new_n600_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n607_), .A2(new_n228_), .A3(new_n233_), .ZN(new_n888_));
  OAI21_X1  g687(.A(new_n887_), .B1(new_n883_), .B2(new_n888_), .ZN(G1351gat));
  NAND2_X1  g688(.A1(new_n846_), .A2(new_n870_), .ZN(new_n890_));
  OAI21_X1  g689(.A(new_n260_), .B1(new_n890_), .B2(new_n500_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT125), .ZN(new_n892_));
  INV_X1    g691(.A(KEYINPUT125), .ZN(new_n893_));
  OAI211_X1 g692(.A(new_n893_), .B(new_n260_), .C1(new_n890_), .C2(new_n500_), .ZN(new_n894_));
  NAND4_X1  g693(.A1(new_n846_), .A2(G197gat), .A3(new_n501_), .A4(new_n870_), .ZN(new_n895_));
  AND3_X1   g694(.A1(new_n892_), .A2(new_n894_), .A3(new_n895_), .ZN(G1352gat));
  NOR2_X1   g695(.A1(new_n890_), .A2(new_n558_), .ZN(new_n897_));
  XNOR2_X1  g696(.A(new_n897_), .B(new_n262_), .ZN(G1353gat));
  AOI21_X1  g697(.A(new_n610_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n899_));
  INV_X1    g698(.A(new_n899_), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT126), .B1(new_n890_), .B2(new_n900_), .ZN(new_n901_));
  INV_X1    g700(.A(KEYINPUT126), .ZN(new_n902_));
  NAND4_X1  g701(.A1(new_n846_), .A2(new_n902_), .A3(new_n870_), .A4(new_n899_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n901_), .A2(new_n903_), .ZN(new_n904_));
  INV_X1    g703(.A(KEYINPUT63), .ZN(new_n905_));
  INV_X1    g704(.A(G211gat), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n904_), .A2(new_n907_), .ZN(new_n908_));
  NAND4_X1  g707(.A1(new_n901_), .A2(new_n905_), .A3(new_n906_), .A4(new_n903_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n908_), .A2(new_n909_), .ZN(G1354gat));
  OAI21_X1  g709(.A(G218gat), .B1(new_n890_), .B2(new_n600_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n608_), .A2(G218gat), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n846_), .A2(new_n870_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n911_), .A2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n911_), .A2(KEYINPUT127), .A3(new_n913_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1355gat));
endmodule


