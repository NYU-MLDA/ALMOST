//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n654_, new_n655_, new_n656_, new_n658_, new_n659_, new_n660_,
    new_n661_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n718_,
    new_n719_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n764_, new_n765_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n878_, new_n879_, new_n881_, new_n882_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n906_, new_n907_, new_n908_, new_n910_, new_n911_,
    new_n913_, new_n914_, new_n916_, new_n917_, new_n918_, new_n920_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n927_, new_n928_,
    new_n929_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  XNOR2_X1  g002(.A(G211gat), .B(G218gat), .ZN(new_n204_));
  INV_X1    g003(.A(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(new_n205_), .A2(KEYINPUT21), .ZN(new_n206_));
  INV_X1    g005(.A(G204gat), .ZN(new_n207_));
  NOR2_X1   g006(.A1(new_n207_), .A2(G197gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(G197gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n209_), .A2(KEYINPUT91), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT91), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n211_), .A2(new_n207_), .A3(G197gat), .ZN(new_n212_));
  AOI21_X1  g011(.A(new_n208_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n206_), .A2(new_n213_), .ZN(new_n214_));
  OR2_X1    g013(.A1(new_n208_), .A2(KEYINPUT90), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n208_), .A2(KEYINPUT90), .ZN(new_n216_));
  NAND3_X1  g015(.A1(new_n215_), .A2(new_n216_), .A3(new_n209_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n217_), .A2(KEYINPUT21), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT21), .ZN(new_n219_));
  AOI21_X1  g018(.A(new_n205_), .B1(new_n213_), .B2(new_n219_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n214_), .B1(new_n218_), .B2(new_n220_), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  XNOR2_X1  g021(.A(KEYINPUT83), .B(KEYINPUT23), .ZN(new_n223_));
  NAND2_X1  g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n223_), .A2(new_n224_), .ZN(new_n225_));
  OR3_X1    g024(.A1(new_n224_), .A2(KEYINPUT84), .A3(KEYINPUT23), .ZN(new_n226_));
  OAI21_X1  g025(.A(KEYINPUT84), .B1(new_n224_), .B2(KEYINPUT23), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  OR2_X1    g027(.A1(G183gat), .A2(G190gat), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G169gat), .A2(G176gat), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G169gat), .ZN(new_n232_));
  INV_X1    g031(.A(new_n232_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n231_), .B1(new_n233_), .B2(G176gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT96), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  AOI21_X1  g035(.A(new_n222_), .B1(new_n230_), .B2(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n224_), .A2(KEYINPUT23), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT87), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n224_), .A2(KEYINPUT87), .A3(KEYINPUT23), .ZN(new_n241_));
  OAI211_X1 g040(.A(new_n240_), .B(new_n241_), .C1(new_n223_), .C2(new_n224_), .ZN(new_n242_));
  INV_X1    g041(.A(G169gat), .ZN(new_n243_));
  INV_X1    g042(.A(G176gat), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n243_), .A2(new_n244_), .ZN(new_n245_));
  NOR2_X1   g044(.A1(new_n245_), .A2(KEYINPUT24), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n242_), .A2(new_n247_), .ZN(new_n248_));
  AND2_X1   g047(.A1(new_n248_), .A2(KEYINPUT95), .ZN(new_n249_));
  NOR2_X1   g048(.A1(new_n248_), .A2(KEYINPUT95), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n231_), .A2(KEYINPUT24), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT93), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n251_), .A2(new_n252_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n252_), .B2(new_n251_), .ZN(new_n254_));
  XNOR2_X1  g053(.A(KEYINPUT26), .B(G190gat), .ZN(new_n255_));
  XNOR2_X1  g054(.A(KEYINPUT25), .B(G183gat), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  AND3_X1   g056(.A1(new_n254_), .A2(KEYINPUT94), .A3(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(KEYINPUT94), .B1(new_n254_), .B2(new_n257_), .ZN(new_n259_));
  OAI22_X1  g058(.A1(new_n249_), .A2(new_n250_), .B1(new_n258_), .B2(new_n259_), .ZN(new_n260_));
  AND2_X1   g059(.A1(new_n237_), .A2(new_n260_), .ZN(new_n261_));
  INV_X1    g060(.A(KEYINPUT20), .ZN(new_n262_));
  XNOR2_X1  g061(.A(KEYINPUT81), .B(G183gat), .ZN(new_n263_));
  INV_X1    g062(.A(G190gat), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  AOI21_X1  g064(.A(G176gat), .B1(new_n243_), .B2(KEYINPUT22), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT22), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(KEYINPUT85), .A3(G169gat), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n266_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(KEYINPUT85), .B1(new_n267_), .B2(G169gat), .ZN(new_n270_));
  OAI21_X1  g069(.A(new_n231_), .B1(new_n269_), .B2(new_n270_), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT86), .ZN(new_n272_));
  AOI22_X1  g071(.A1(new_n242_), .A2(new_n265_), .B1(new_n271_), .B2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(new_n273_), .B1(new_n272_), .B2(new_n271_), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT25), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n263_), .A2(new_n275_), .ZN(new_n276_));
  NOR2_X1   g075(.A1(KEYINPUT25), .A2(G183gat), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n255_), .B1(new_n276_), .B2(new_n277_), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n245_), .A2(KEYINPUT24), .A3(new_n231_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n279_), .A2(KEYINPUT82), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n246_), .B1(new_n279_), .B2(KEYINPUT82), .ZN(new_n281_));
  NAND4_X1  g080(.A1(new_n278_), .A2(new_n228_), .A3(new_n280_), .A4(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n274_), .A2(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(new_n262_), .B1(new_n283_), .B2(new_n222_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n284_), .ZN(new_n285_));
  OAI21_X1  g084(.A(new_n203_), .B1(new_n261_), .B2(new_n285_), .ZN(new_n286_));
  OAI21_X1  g085(.A(KEYINPUT20), .B1(new_n283_), .B2(new_n222_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT97), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n234_), .B(KEYINPUT96), .ZN(new_n289_));
  INV_X1    g088(.A(new_n230_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n288_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND3_X1  g090(.A1(new_n236_), .A2(KEYINPUT97), .A3(new_n230_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n291_), .A2(new_n260_), .A3(new_n292_), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n287_), .B1(new_n222_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(new_n203_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(new_n286_), .ZN(new_n297_));
  MUX2_X1   g096(.A(new_n286_), .B(new_n297_), .S(KEYINPUT106), .Z(new_n298_));
  XNOR2_X1  g097(.A(G8gat), .B(G36gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT18), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G64gat), .B(G92gat), .ZN(new_n301_));
  XOR2_X1   g100(.A(new_n300_), .B(new_n301_), .Z(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n298_), .A2(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(KEYINPUT98), .B1(new_n294_), .B2(new_n295_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n293_), .A2(new_n222_), .ZN(new_n306_));
  AND2_X1   g105(.A1(new_n274_), .A2(new_n282_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n262_), .B1(new_n307_), .B2(new_n221_), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n306_), .A2(new_n308_), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT98), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n309_), .A2(new_n310_), .A3(new_n203_), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n305_), .A2(new_n311_), .ZN(new_n312_));
  NAND4_X1  g111(.A1(new_n291_), .A2(new_n260_), .A3(new_n292_), .A4(new_n221_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(new_n284_), .A3(new_n295_), .ZN(new_n314_));
  INV_X1    g113(.A(KEYINPUT99), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n314_), .A2(new_n315_), .ZN(new_n316_));
  NAND4_X1  g115(.A1(new_n313_), .A2(new_n284_), .A3(KEYINPUT99), .A4(new_n295_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n316_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n312_), .A2(new_n302_), .A3(new_n318_), .ZN(new_n319_));
  NAND3_X1  g118(.A1(new_n304_), .A2(KEYINPUT27), .A3(new_n319_), .ZN(new_n320_));
  NOR3_X1   g119(.A1(new_n294_), .A2(KEYINPUT98), .A3(new_n295_), .ZN(new_n321_));
  AOI21_X1  g120(.A(new_n310_), .B1(new_n309_), .B2(new_n203_), .ZN(new_n322_));
  OAI21_X1  g121(.A(new_n318_), .B1(new_n321_), .B2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(new_n303_), .ZN(new_n324_));
  AOI21_X1  g123(.A(KEYINPUT27), .B1(new_n324_), .B2(new_n319_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n320_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328_));
  NOR2_X1   g127(.A1(G155gat), .A2(G162gat), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331_));
  XOR2_X1   g130(.A(new_n331_), .B(KEYINPUT3), .Z(new_n332_));
  NAND2_X1  g131(.A1(G141gat), .A2(G148gat), .ZN(new_n333_));
  XOR2_X1   g132(.A(new_n333_), .B(KEYINPUT2), .Z(new_n334_));
  OAI211_X1 g133(.A(new_n328_), .B(new_n330_), .C1(new_n332_), .C2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n329_), .B1(KEYINPUT1), .B2(new_n328_), .ZN(new_n336_));
  OAI21_X1  g135(.A(new_n336_), .B1(KEYINPUT1), .B2(new_n328_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n331_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n337_), .A2(new_n338_), .A3(new_n333_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n339_), .ZN(new_n340_));
  NOR2_X1   g139(.A1(new_n340_), .A2(KEYINPUT29), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT28), .ZN(new_n342_));
  XOR2_X1   g141(.A(G22gat), .B(G50gat), .Z(new_n343_));
  XNOR2_X1  g142(.A(new_n342_), .B(new_n343_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(new_n344_), .B(KEYINPUT89), .ZN(new_n345_));
  AOI21_X1  g144(.A(new_n221_), .B1(KEYINPUT29), .B2(new_n340_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G228gat), .A2(G233gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n346_), .B(new_n347_), .Z(new_n348_));
  XNOR2_X1  g147(.A(G78gat), .B(G106gat), .ZN(new_n349_));
  XOR2_X1   g148(.A(new_n348_), .B(new_n349_), .Z(new_n350_));
  NAND2_X1  g149(.A1(new_n345_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT92), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n349_), .A2(new_n352_), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n348_), .A2(new_n353_), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n348_), .A2(new_n353_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n354_), .A2(new_n344_), .A3(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n351_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(G227gat), .A2(G233gat), .ZN(new_n358_));
  XNOR2_X1  g157(.A(new_n358_), .B(G15gat), .ZN(new_n359_));
  XOR2_X1   g158(.A(new_n359_), .B(KEYINPUT30), .Z(new_n360_));
  XNOR2_X1  g159(.A(new_n283_), .B(new_n360_), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G127gat), .B(G134gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(G113gat), .B(G120gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n362_), .B(new_n363_), .ZN(new_n364_));
  XNOR2_X1  g163(.A(new_n364_), .B(KEYINPUT88), .ZN(new_n365_));
  XNOR2_X1  g164(.A(new_n361_), .B(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G71gat), .B(G99gat), .ZN(new_n367_));
  INV_X1    g166(.A(G43gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  XNOR2_X1  g168(.A(new_n369_), .B(KEYINPUT31), .ZN(new_n370_));
  OR2_X1    g169(.A1(new_n366_), .A2(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n370_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n365_), .A2(new_n340_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n335_), .A2(new_n364_), .A3(new_n339_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(KEYINPUT4), .ZN(new_n377_));
  AOI21_X1  g176(.A(KEYINPUT4), .B1(new_n365_), .B2(new_n340_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND4_X1  g178(.A1(new_n377_), .A2(G225gat), .A3(G233gat), .A4(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(G225gat), .A2(G233gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n376_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n380_), .A2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(G1gat), .B(G29gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G85gat), .ZN(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT0), .B(G57gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  INV_X1    g186(.A(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n380_), .A2(new_n387_), .A3(new_n382_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n373_), .A2(new_n392_), .ZN(new_n393_));
  NOR3_X1   g192(.A1(new_n327_), .A2(new_n357_), .A3(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n357_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n302_), .A2(KEYINPUT32), .ZN(new_n396_));
  INV_X1    g195(.A(new_n396_), .ZN(new_n397_));
  AOI21_X1  g196(.A(new_n392_), .B1(new_n298_), .B2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n398_), .B1(new_n323_), .B2(new_n397_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n387_), .B1(new_n376_), .B2(new_n381_), .ZN(new_n400_));
  INV_X1    g199(.A(KEYINPUT102), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  OAI211_X1 g201(.A(KEYINPUT102), .B(new_n387_), .C1(new_n376_), .C2(new_n381_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT4), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n406_));
  OAI211_X1 g205(.A(KEYINPUT103), .B(new_n381_), .C1(new_n406_), .C2(new_n378_), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n381_), .B1(new_n406_), .B2(new_n378_), .ZN(new_n408_));
  INV_X1    g207(.A(KEYINPUT103), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n404_), .A2(new_n407_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(KEYINPUT104), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT104), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n404_), .A2(new_n410_), .A3(new_n413_), .A4(new_n407_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n389_), .A2(KEYINPUT101), .A3(KEYINPUT33), .ZN(new_n416_));
  OR2_X1    g215(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n417_));
  NAND2_X1  g216(.A1(KEYINPUT101), .A2(KEYINPUT33), .ZN(new_n418_));
  NAND4_X1  g217(.A1(new_n383_), .A2(new_n388_), .A3(new_n417_), .A4(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n416_), .A2(new_n419_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n415_), .A2(new_n420_), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT100), .ZN(new_n422_));
  NOR2_X1   g221(.A1(new_n323_), .A2(new_n303_), .ZN(new_n423_));
  AOI21_X1  g222(.A(new_n302_), .B1(new_n312_), .B2(new_n318_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n324_), .A2(KEYINPUT100), .A3(new_n319_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n421_), .B1(new_n425_), .B2(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n399_), .B1(new_n427_), .B2(KEYINPUT105), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT105), .ZN(new_n429_));
  AOI211_X1 g228(.A(new_n429_), .B(new_n421_), .C1(new_n425_), .C2(new_n426_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n395_), .B1(new_n428_), .B2(new_n430_), .ZN(new_n431_));
  NOR3_X1   g230(.A1(new_n327_), .A2(new_n391_), .A3(new_n395_), .ZN(new_n432_));
  INV_X1    g231(.A(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n431_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n373_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n394_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G29gat), .B(G36gat), .ZN(new_n437_));
  AND2_X1   g236(.A1(new_n437_), .A2(KEYINPUT71), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n437_), .A2(KEYINPUT71), .ZN(new_n439_));
  XOR2_X1   g238(.A(G43gat), .B(G50gat), .Z(new_n440_));
  OR3_X1    g239(.A1(new_n438_), .A2(new_n439_), .A3(new_n440_), .ZN(new_n441_));
  OAI21_X1  g240(.A(new_n440_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n441_), .A2(new_n442_), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(KEYINPUT15), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  XNOR2_X1  g244(.A(KEYINPUT76), .B(G15gat), .ZN(new_n446_));
  INV_X1    g245(.A(G22gat), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n446_), .B(new_n447_), .ZN(new_n448_));
  INV_X1    g247(.A(G1gat), .ZN(new_n449_));
  INV_X1    g248(.A(G8gat), .ZN(new_n450_));
  OAI21_X1  g249(.A(KEYINPUT14), .B1(new_n449_), .B2(new_n450_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n448_), .A2(new_n451_), .ZN(new_n452_));
  XOR2_X1   g251(.A(G1gat), .B(G8gat), .Z(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n454_), .ZN(new_n455_));
  NAND2_X1  g254(.A1(new_n445_), .A2(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n443_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT79), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT79), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n443_), .A2(new_n459_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n458_), .A2(new_n454_), .A3(new_n460_), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G229gat), .A2(G233gat), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n456_), .A2(new_n461_), .A3(new_n462_), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G113gat), .B(G141gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G169gat), .B(G197gat), .ZN(new_n465_));
  XOR2_X1   g264(.A(new_n464_), .B(new_n465_), .Z(new_n466_));
  NOR2_X1   g265(.A1(new_n466_), .A2(KEYINPUT80), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n462_), .ZN(new_n469_));
  AND3_X1   g268(.A1(new_n458_), .A2(new_n454_), .A3(new_n460_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n454_), .B1(new_n458_), .B2(new_n460_), .ZN(new_n471_));
  OAI21_X1  g270(.A(new_n469_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  AND3_X1   g271(.A1(new_n463_), .A2(new_n468_), .A3(new_n472_), .ZN(new_n473_));
  AOI21_X1  g272(.A(new_n468_), .B1(new_n463_), .B2(new_n472_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n473_), .A2(new_n474_), .ZN(new_n475_));
  NOR2_X1   g274(.A1(new_n436_), .A2(new_n475_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(G232gat), .A2(G233gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT34), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n478_), .A2(KEYINPUT35), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT73), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n479_), .A2(new_n480_), .ZN(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n478_), .A2(KEYINPUT73), .A3(KEYINPUT35), .ZN(new_n483_));
  OR2_X1    g282(.A1(new_n478_), .A2(KEYINPUT35), .ZN(new_n484_));
  XNOR2_X1  g283(.A(G85gat), .B(G92gat), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(G99gat), .A2(G106gat), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n487_), .A2(KEYINPUT6), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n489_), .A2(G99gat), .A3(G106gat), .ZN(new_n490_));
  AND2_X1   g289(.A1(new_n488_), .A2(new_n490_), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n492_));
  INV_X1    g291(.A(G99gat), .ZN(new_n493_));
  INV_X1    g292(.A(G106gat), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n492_), .A2(new_n493_), .A3(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n495_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n486_), .B1(new_n491_), .B2(new_n497_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(KEYINPUT8), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n488_), .A2(new_n490_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n500_), .A2(new_n496_), .A3(new_n495_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT8), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n501_), .A2(new_n502_), .A3(new_n486_), .ZN(new_n503_));
  OR2_X1    g302(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n504_));
  NAND2_X1  g303(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n494_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT64), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  AND2_X1   g307(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n511_), .A2(KEYINPUT64), .A3(new_n494_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n491_), .B1(new_n508_), .B2(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(G85gat), .A2(G92gat), .ZN(new_n514_));
  AND2_X1   g313(.A1(G85gat), .A2(G92gat), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n514_), .B1(new_n515_), .B2(KEYINPUT9), .ZN(new_n516_));
  OAI21_X1  g315(.A(KEYINPUT65), .B1(new_n515_), .B2(KEYINPUT9), .ZN(new_n517_));
  NAND2_X1  g316(.A1(G85gat), .A2(G92gat), .ZN(new_n518_));
  INV_X1    g317(.A(KEYINPUT65), .ZN(new_n519_));
  INV_X1    g318(.A(KEYINPUT9), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n518_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n516_), .A2(new_n517_), .A3(new_n521_), .ZN(new_n522_));
  AOI22_X1  g321(.A1(new_n499_), .A2(new_n503_), .B1(new_n513_), .B2(new_n522_), .ZN(new_n523_));
  OAI211_X1 g322(.A(new_n483_), .B(new_n484_), .C1(new_n444_), .C2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(KEYINPUT66), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n499_), .A2(new_n503_), .ZN(new_n526_));
  AOI21_X1  g325(.A(KEYINPUT64), .B1(new_n511_), .B2(new_n494_), .ZN(new_n527_));
  NOR4_X1   g326(.A1(new_n509_), .A2(new_n510_), .A3(new_n507_), .A4(G106gat), .ZN(new_n528_));
  OAI211_X1 g327(.A(new_n522_), .B(new_n500_), .C1(new_n527_), .C2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n525_), .B1(new_n526_), .B2(new_n529_), .ZN(new_n530_));
  AND2_X1   g329(.A1(new_n495_), .A2(new_n496_), .ZN(new_n531_));
  AOI211_X1 g330(.A(KEYINPUT8), .B(new_n485_), .C1(new_n531_), .C2(new_n500_), .ZN(new_n532_));
  AOI21_X1  g331(.A(new_n502_), .B1(new_n501_), .B2(new_n486_), .ZN(new_n533_));
  OAI211_X1 g332(.A(new_n529_), .B(new_n525_), .C1(new_n532_), .C2(new_n533_), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n530_), .A2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n536_), .A2(new_n457_), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n537_), .A2(KEYINPUT72), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT72), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n536_), .A2(new_n539_), .A3(new_n457_), .ZN(new_n540_));
  AOI211_X1 g339(.A(new_n482_), .B(new_n524_), .C1(new_n538_), .C2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n538_), .A2(new_n540_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n524_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n481_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n541_), .A2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT75), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(G190gat), .B(G218gat), .ZN(new_n548_));
  XNOR2_X1  g347(.A(G134gat), .B(G162gat), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n548_), .B(new_n549_), .ZN(new_n550_));
  XOR2_X1   g349(.A(new_n550_), .B(KEYINPUT36), .Z(new_n551_));
  OAI21_X1  g350(.A(KEYINPUT75), .B1(new_n541_), .B2(new_n544_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n547_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT37), .ZN(new_n554_));
  NOR2_X1   g353(.A1(new_n550_), .A2(KEYINPUT36), .ZN(new_n555_));
  OAI21_X1  g354(.A(new_n555_), .B1(new_n541_), .B2(new_n544_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n553_), .A2(new_n554_), .A3(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT74), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n542_), .A2(new_n543_), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n559_), .A2(new_n482_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n542_), .A2(new_n481_), .A3(new_n543_), .ZN(new_n561_));
  NAND3_X1  g360(.A1(new_n560_), .A2(new_n561_), .A3(new_n551_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n558_), .B1(new_n556_), .B2(new_n562_), .ZN(new_n563_));
  AOI21_X1  g362(.A(KEYINPUT74), .B1(new_n545_), .B2(new_n551_), .ZN(new_n564_));
  OAI21_X1  g363(.A(KEYINPUT37), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n557_), .A2(new_n565_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(G57gat), .B(G64gat), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n567_), .A2(KEYINPUT11), .ZN(new_n568_));
  XNOR2_X1  g367(.A(G71gat), .B(G78gat), .ZN(new_n569_));
  INV_X1    g368(.A(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n568_), .A2(new_n570_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n567_), .A2(KEYINPUT11), .ZN(new_n572_));
  OR2_X1    g371(.A1(new_n571_), .A2(new_n572_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n567_), .A2(new_n569_), .A3(KEYINPUT11), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n573_), .A2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(new_n454_), .B(new_n575_), .ZN(new_n576_));
  AND2_X1   g375(.A1(G231gat), .A2(G233gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(KEYINPUT17), .ZN(new_n579_));
  XOR2_X1   g378(.A(G127gat), .B(G155gat), .Z(new_n580_));
  XNOR2_X1  g379(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n580_), .B(new_n581_), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G183gat), .B(G211gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  OR3_X1    g383(.A1(new_n578_), .A2(new_n579_), .A3(new_n584_), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n584_), .B(KEYINPUT17), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n578_), .A2(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n585_), .A2(new_n587_), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n588_), .B(KEYINPUT78), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n566_), .A2(new_n589_), .ZN(new_n590_));
  OAI211_X1 g389(.A(KEYINPUT12), .B(new_n574_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n591_));
  OAI21_X1  g390(.A(KEYINPUT67), .B1(new_n523_), .B2(new_n591_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n529_), .B1(new_n532_), .B2(new_n533_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT67), .ZN(new_n594_));
  INV_X1    g393(.A(new_n591_), .ZN(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n594_), .A3(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n592_), .A2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n593_), .A2(KEYINPUT66), .ZN(new_n598_));
  AOI21_X1  g397(.A(new_n575_), .B1(new_n598_), .B2(new_n534_), .ZN(new_n599_));
  OAI21_X1  g398(.A(new_n597_), .B1(new_n599_), .B2(KEYINPUT12), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n598_), .A2(new_n575_), .A3(new_n534_), .ZN(new_n601_));
  NAND2_X1  g400(.A1(G230gat), .A2(G233gat), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT68), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NAND3_X1  g404(.A1(new_n601_), .A2(KEYINPUT68), .A3(new_n602_), .ZN(new_n606_));
  AOI21_X1  g405(.A(new_n600_), .B1(new_n605_), .B2(new_n606_), .ZN(new_n607_));
  INV_X1    g406(.A(new_n599_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n602_), .B1(new_n608_), .B2(new_n601_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n607_), .A2(new_n609_), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G120gat), .B(G148gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT5), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G176gat), .B(G204gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(KEYINPUT69), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  XOR2_X1   g417(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT13), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n615_), .B(new_n617_), .C1(KEYINPUT70), .C2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n620_), .A2(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n590_), .A2(new_n624_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n476_), .A2(new_n625_), .ZN(new_n626_));
  NOR3_X1   g425(.A1(new_n626_), .A2(G1gat), .A3(new_n392_), .ZN(new_n627_));
  OR2_X1    g426(.A1(new_n627_), .A2(KEYINPUT38), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n627_), .A2(KEYINPUT38), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n553_), .A2(new_n556_), .ZN(new_n630_));
  INV_X1    g429(.A(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n436_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n475_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n623_), .A2(new_n633_), .ZN(new_n634_));
  NOR2_X1   g433(.A1(new_n634_), .A2(new_n588_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n632_), .A2(new_n635_), .ZN(new_n636_));
  OAI21_X1  g435(.A(G1gat), .B1(new_n636_), .B2(new_n392_), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n628_), .A2(new_n629_), .A3(new_n637_), .ZN(G1324gat));
  INV_X1    g437(.A(new_n626_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n639_), .A2(new_n450_), .A3(new_n327_), .ZN(new_n640_));
  INV_X1    g439(.A(new_n327_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n636_), .A2(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(new_n450_), .B1(new_n642_), .B2(KEYINPUT107), .ZN(new_n643_));
  INV_X1    g442(.A(KEYINPUT39), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT107), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n645_), .B1(new_n636_), .B2(new_n641_), .ZN(new_n646_));
  AND3_X1   g445(.A1(new_n643_), .A2(new_n644_), .A3(new_n646_), .ZN(new_n647_));
  AOI21_X1  g446(.A(new_n644_), .B1(new_n643_), .B2(new_n646_), .ZN(new_n648_));
  OAI21_X1  g447(.A(new_n640_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT40), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  OAI211_X1 g450(.A(KEYINPUT40), .B(new_n640_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n652_));
  NAND2_X1  g451(.A1(new_n651_), .A2(new_n652_), .ZN(G1325gat));
  OAI21_X1  g452(.A(G15gat), .B1(new_n636_), .B2(new_n435_), .ZN(new_n654_));
  XNOR2_X1  g453(.A(new_n654_), .B(KEYINPUT41), .ZN(new_n655_));
  NOR3_X1   g454(.A1(new_n626_), .A2(G15gat), .A3(new_n435_), .ZN(new_n656_));
  OR2_X1    g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1326gat));
  OAI21_X1  g456(.A(G22gat), .B1(new_n636_), .B2(new_n395_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n658_), .B(KEYINPUT42), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n639_), .A2(new_n447_), .A3(new_n357_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n659_), .A2(new_n660_), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n661_), .B(KEYINPUT108), .ZN(G1327gat));
  INV_X1    g461(.A(new_n394_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n415_), .A2(new_n420_), .ZN(new_n664_));
  NOR3_X1   g463(.A1(new_n423_), .A2(new_n424_), .A3(new_n422_), .ZN(new_n665_));
  AOI21_X1  g464(.A(KEYINPUT100), .B1(new_n324_), .B2(new_n319_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n664_), .B1(new_n665_), .B2(new_n666_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(new_n429_), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n427_), .A2(KEYINPUT105), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n668_), .A2(new_n669_), .A3(new_n399_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n432_), .B1(new_n670_), .B2(new_n395_), .ZN(new_n671_));
  OAI21_X1  g470(.A(new_n663_), .B1(new_n671_), .B2(new_n373_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n589_), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n673_), .A2(new_n631_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n674_), .A2(new_n624_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n672_), .A2(new_n633_), .A3(new_n675_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  AOI21_X1  g476(.A(G29gat), .B1(new_n677_), .B2(new_n391_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT43), .ZN(new_n679_));
  INV_X1    g478(.A(new_n566_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n373_), .B1(new_n431_), .B2(new_n433_), .ZN(new_n681_));
  OAI211_X1 g480(.A(new_n679_), .B(new_n680_), .C1(new_n681_), .C2(new_n394_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n436_), .B2(new_n566_), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n672_), .A2(KEYINPUT109), .A3(new_n679_), .A4(new_n680_), .ZN(new_n686_));
  NAND3_X1  g485(.A1(new_n684_), .A2(new_n685_), .A3(new_n686_), .ZN(new_n687_));
  NOR2_X1   g486(.A1(new_n589_), .A2(new_n634_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n689_), .A2(new_n690_), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n687_), .A2(KEYINPUT44), .A3(new_n688_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n691_), .A2(new_n692_), .ZN(new_n693_));
  AND2_X1   g492(.A1(new_n391_), .A2(G29gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n678_), .B1(new_n693_), .B2(new_n694_), .ZN(G1328gat));
  OR2_X1    g494(.A1(new_n641_), .A2(G36gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n676_), .A2(new_n696_), .ZN(new_n697_));
  INV_X1    g496(.A(KEYINPUT45), .ZN(new_n698_));
  XNOR2_X1  g497(.A(new_n697_), .B(new_n698_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT46), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT110), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  NAND3_X1  g501(.A1(new_n691_), .A2(new_n327_), .A3(new_n692_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n703_), .B2(G36gat), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n700_), .A2(KEYINPUT110), .ZN(new_n705_));
  XNOR2_X1  g504(.A(new_n704_), .B(new_n705_), .ZN(G1329gat));
  NOR2_X1   g505(.A1(new_n435_), .A2(new_n368_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n691_), .A2(new_n692_), .A3(new_n707_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT111), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND4_X1  g509(.A1(new_n691_), .A2(KEYINPUT111), .A3(new_n692_), .A4(new_n707_), .ZN(new_n711_));
  OAI21_X1  g510(.A(new_n368_), .B1(new_n676_), .B2(new_n435_), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n710_), .A2(new_n711_), .A3(new_n712_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n713_), .A2(KEYINPUT47), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT47), .ZN(new_n715_));
  NAND4_X1  g514(.A1(new_n710_), .A2(new_n715_), .A3(new_n711_), .A4(new_n712_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(new_n716_), .ZN(G1330gat));
  AOI21_X1  g516(.A(G50gat), .B1(new_n677_), .B2(new_n357_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n357_), .A2(G50gat), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n718_), .B1(new_n693_), .B2(new_n719_), .ZN(G1331gat));
  INV_X1    g519(.A(G57gat), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n623_), .A2(new_n633_), .ZN(new_n722_));
  NAND3_X1  g521(.A1(new_n632_), .A2(new_n589_), .A3(new_n722_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT113), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  NAND4_X1  g524(.A1(new_n632_), .A2(KEYINPUT113), .A3(new_n589_), .A4(new_n722_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n721_), .B1(new_n727_), .B2(new_n391_), .ZN(new_n728_));
  NOR2_X1   g527(.A1(new_n436_), .A2(new_n633_), .ZN(new_n729_));
  NOR2_X1   g528(.A1(new_n590_), .A2(new_n623_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT112), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n732_), .A2(G57gat), .A3(new_n392_), .ZN(new_n733_));
  OR2_X1    g532(.A1(new_n728_), .A2(new_n733_), .ZN(G1332gat));
  OR3_X1    g533(.A1(new_n732_), .A2(G64gat), .A3(new_n641_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n725_), .A2(new_n327_), .A3(new_n726_), .ZN(new_n736_));
  INV_X1    g535(.A(KEYINPUT48), .ZN(new_n737_));
  AND3_X1   g536(.A1(new_n736_), .A2(new_n737_), .A3(G64gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n737_), .B1(new_n736_), .B2(G64gat), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n735_), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n740_), .A2(KEYINPUT114), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT114), .ZN(new_n742_));
  OAI211_X1 g541(.A(new_n742_), .B(new_n735_), .C1(new_n738_), .C2(new_n739_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n741_), .A2(new_n743_), .ZN(G1333gat));
  OR3_X1    g543(.A1(new_n732_), .A2(G71gat), .A3(new_n435_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n727_), .A2(new_n373_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n746_), .A2(G71gat), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n747_), .A2(KEYINPUT49), .ZN(new_n748_));
  NOR2_X1   g547(.A1(new_n747_), .A2(KEYINPUT49), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n745_), .B1(new_n748_), .B2(new_n749_), .ZN(G1334gat));
  OR3_X1    g549(.A1(new_n732_), .A2(G78gat), .A3(new_n395_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n727_), .A2(new_n357_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n752_), .A2(G78gat), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n753_), .A2(KEYINPUT50), .ZN(new_n754_));
  NOR2_X1   g553(.A1(new_n753_), .A2(KEYINPUT50), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(G1335gat));
  NOR3_X1   g555(.A1(new_n589_), .A2(new_n633_), .A3(new_n623_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n687_), .A2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G85gat), .B1(new_n758_), .B2(new_n392_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n674_), .A2(new_n623_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n729_), .A2(new_n760_), .ZN(new_n761_));
  OR2_X1    g560(.A1(new_n392_), .A2(G85gat), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n759_), .B1(new_n761_), .B2(new_n762_), .ZN(G1336gat));
  OAI21_X1  g562(.A(G92gat), .B1(new_n758_), .B2(new_n641_), .ZN(new_n764_));
  OR2_X1    g563(.A1(new_n641_), .A2(G92gat), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n764_), .B1(new_n761_), .B2(new_n765_), .ZN(G1337gat));
  OAI21_X1  g565(.A(G99gat), .B1(new_n758_), .B2(new_n435_), .ZN(new_n767_));
  INV_X1    g566(.A(new_n761_), .ZN(new_n768_));
  NAND3_X1  g567(.A1(new_n768_), .A2(new_n373_), .A3(new_n511_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n767_), .A2(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g570(.A1(new_n768_), .A2(new_n494_), .A3(new_n357_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n687_), .A2(new_n357_), .A3(new_n757_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774_));
  AND3_X1   g573(.A1(new_n773_), .A2(new_n774_), .A3(G106gat), .ZN(new_n775_));
  AOI21_X1  g574(.A(new_n774_), .B1(new_n773_), .B2(G106gat), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n772_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND4_X1  g577(.A1(new_n566_), .A2(new_n475_), .A3(new_n623_), .A4(new_n589_), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT54), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n779_), .B(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT55), .B1(new_n607_), .B2(KEYINPUT115), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784_));
  AND3_X1   g583(.A1(new_n601_), .A2(KEYINPUT68), .A3(new_n602_), .ZN(new_n785_));
  AOI21_X1  g584(.A(KEYINPUT68), .B1(new_n601_), .B2(new_n602_), .ZN(new_n786_));
  NOR2_X1   g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(new_n783_), .B(new_n784_), .C1(new_n787_), .C2(new_n600_), .ZN(new_n788_));
  INV_X1    g587(.A(new_n601_), .ZN(new_n789_));
  OAI211_X1 g588(.A(G230gat), .B(G233gat), .C1(new_n600_), .C2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n782_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n791_));
  AND3_X1   g590(.A1(new_n791_), .A2(KEYINPUT56), .A3(new_n616_), .ZN(new_n792_));
  AOI21_X1  g591(.A(KEYINPUT56), .B1(new_n791_), .B2(new_n616_), .ZN(new_n793_));
  OR2_X1    g592(.A1(new_n792_), .A2(new_n793_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n460_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n443_), .A2(new_n459_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n455_), .B1(new_n795_), .B2(new_n796_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n469_), .B1(new_n797_), .B2(new_n461_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT117), .B1(new_n798_), .B2(new_n466_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n462_), .B1(new_n470_), .B2(new_n471_), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801_));
  INV_X1    g600(.A(new_n466_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n801_), .A3(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n456_), .A2(new_n461_), .A3(new_n469_), .ZN(new_n804_));
  NAND3_X1  g603(.A1(new_n799_), .A2(new_n803_), .A3(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n463_), .A2(new_n466_), .A3(new_n472_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT118), .ZN(new_n808_));
  XNOR2_X1  g607(.A(new_n807_), .B(new_n808_), .ZN(new_n809_));
  NAND3_X1  g608(.A1(new_n794_), .A2(new_n615_), .A3(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT58), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  NAND4_X1  g611(.A1(new_n794_), .A2(KEYINPUT58), .A3(new_n615_), .A4(new_n809_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n812_), .A2(new_n680_), .A3(new_n813_), .ZN(new_n814_));
  NOR2_X1   g613(.A1(KEYINPUT119), .A2(KEYINPUT57), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n475_), .B1(new_n610_), .B2(new_n614_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(new_n792_), .B2(new_n793_), .ZN(new_n818_));
  AOI22_X1  g617(.A1(new_n818_), .A2(KEYINPUT116), .B1(new_n618_), .B2(new_n809_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n817_), .B(new_n820_), .C1(new_n792_), .C2(new_n793_), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n631_), .B(new_n816_), .C1(new_n819_), .C2(new_n821_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n818_), .A2(KEYINPUT116), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n809_), .A2(new_n618_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n821_), .A3(new_n824_), .ZN(new_n825_));
  AOI21_X1  g624(.A(new_n815_), .B1(new_n825_), .B2(new_n630_), .ZN(new_n826_));
  OAI21_X1  g625(.A(new_n814_), .B1(new_n822_), .B2(new_n826_), .ZN(new_n827_));
  AOI21_X1  g626(.A(new_n781_), .B1(new_n827_), .B2(new_n588_), .ZN(new_n828_));
  NOR2_X1   g627(.A1(new_n327_), .A2(new_n357_), .ZN(new_n829_));
  NAND3_X1  g628(.A1(new_n829_), .A2(new_n391_), .A3(new_n373_), .ZN(new_n830_));
  OAI21_X1  g629(.A(KEYINPUT59), .B1(new_n828_), .B2(new_n830_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n831_), .A2(KEYINPUT120), .ZN(new_n832_));
  INV_X1    g631(.A(KEYINPUT120), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n833_), .B(KEYINPUT59), .C1(new_n828_), .C2(new_n830_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n832_), .A2(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n781_), .B1(new_n827_), .B2(new_n673_), .ZN(new_n836_));
  NOR3_X1   g635(.A1(new_n836_), .A2(KEYINPUT59), .A3(new_n830_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n835_), .A2(new_n838_), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n839_), .A2(KEYINPUT121), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n835_), .A2(new_n841_), .A3(new_n838_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n840_), .A2(new_n842_), .ZN(new_n843_));
  OAI21_X1  g642(.A(G113gat), .B1(new_n843_), .B2(new_n475_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n828_), .ZN(new_n845_));
  INV_X1    g644(.A(new_n830_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  INV_X1    g647(.A(G113gat), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n633_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n844_), .A2(new_n850_), .ZN(G1340gat));
  OAI21_X1  g650(.A(G120gat), .B1(new_n839_), .B2(new_n623_), .ZN(new_n852_));
  INV_X1    g651(.A(G120gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n853_), .B1(new_n623_), .B2(KEYINPUT60), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n854_), .B1(KEYINPUT60), .B2(new_n853_), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n852_), .B1(new_n847_), .B2(new_n855_), .ZN(G1341gat));
  INV_X1    g655(.A(KEYINPUT122), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n841_), .B1(new_n835_), .B2(new_n838_), .ZN(new_n858_));
  AOI211_X1 g657(.A(KEYINPUT121), .B(new_n837_), .C1(new_n832_), .C2(new_n834_), .ZN(new_n859_));
  INV_X1    g658(.A(new_n588_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n860_), .A2(G127gat), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n858_), .A2(new_n859_), .A3(new_n861_), .ZN(new_n862_));
  AOI21_X1  g661(.A(G127gat), .B1(new_n848_), .B2(new_n589_), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n857_), .B1(new_n862_), .B2(new_n863_), .ZN(new_n864_));
  INV_X1    g663(.A(new_n863_), .ZN(new_n865_));
  OAI211_X1 g664(.A(KEYINPUT122), .B(new_n865_), .C1(new_n843_), .C2(new_n861_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n864_), .A2(new_n866_), .ZN(G1342gat));
  OAI21_X1  g666(.A(G134gat), .B1(new_n843_), .B2(new_n566_), .ZN(new_n868_));
  OR3_X1    g667(.A1(new_n847_), .A2(G134gat), .A3(new_n630_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1343gat));
  NAND4_X1  g669(.A1(new_n641_), .A2(new_n391_), .A3(new_n357_), .A4(new_n435_), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n871_), .B(KEYINPUT123), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n828_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n873_), .A2(new_n874_), .ZN(new_n875_));
  NOR3_X1   g674(.A1(new_n828_), .A2(KEYINPUT124), .A3(new_n872_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n875_), .A2(new_n876_), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n877_), .A2(new_n475_), .ZN(new_n878_));
  XNOR2_X1  g677(.A(KEYINPUT125), .B(G141gat), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n878_), .B(new_n879_), .ZN(G1344gat));
  OR2_X1    g679(.A1(new_n875_), .A2(new_n876_), .ZN(new_n881_));
  NAND2_X1  g680(.A1(new_n881_), .A2(new_n624_), .ZN(new_n882_));
  XNOR2_X1  g681(.A(new_n882_), .B(G148gat), .ZN(G1345gat));
  NOR2_X1   g682(.A1(new_n877_), .A2(new_n673_), .ZN(new_n884_));
  XOR2_X1   g683(.A(KEYINPUT61), .B(G155gat), .Z(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(G1346gat));
  INV_X1    g685(.A(G162gat), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n881_), .A2(new_n887_), .A3(new_n631_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n877_), .A2(new_n566_), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n888_), .B1(new_n887_), .B2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT126), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n892_));
  OAI211_X1 g691(.A(new_n888_), .B(new_n892_), .C1(new_n887_), .C2(new_n889_), .ZN(new_n893_));
  AND2_X1   g692(.A1(new_n891_), .A2(new_n893_), .ZN(G1347gat));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n895_));
  NOR2_X1   g694(.A1(new_n641_), .A2(new_n393_), .ZN(new_n896_));
  INV_X1    g695(.A(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n357_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  NOR2_X1   g698(.A1(new_n836_), .A2(new_n899_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n633_), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n895_), .B1(new_n902_), .B2(new_n243_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n901_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n904_));
  OAI211_X1 g703(.A(new_n903_), .B(new_n904_), .C1(new_n233_), .C2(new_n901_), .ZN(G1348gat));
  AOI21_X1  g704(.A(G176gat), .B1(new_n900_), .B2(new_n624_), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n828_), .A2(new_n357_), .ZN(new_n907_));
  NOR3_X1   g706(.A1(new_n897_), .A2(new_n244_), .A3(new_n623_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n906_), .B1(new_n907_), .B2(new_n908_), .ZN(G1349gat));
  NAND3_X1  g708(.A1(new_n907_), .A2(new_n589_), .A3(new_n896_), .ZN(new_n910_));
  NOR2_X1   g709(.A1(new_n588_), .A2(new_n256_), .ZN(new_n911_));
  AOI22_X1  g710(.A1(new_n910_), .A2(new_n263_), .B1(new_n900_), .B2(new_n911_), .ZN(G1350gat));
  NAND3_X1  g711(.A1(new_n900_), .A2(new_n255_), .A3(new_n631_), .ZN(new_n913_));
  NOR3_X1   g712(.A1(new_n836_), .A2(new_n566_), .A3(new_n899_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n913_), .B1(new_n914_), .B2(new_n264_), .ZN(G1351gat));
  NAND2_X1  g714(.A1(new_n357_), .A2(new_n392_), .ZN(new_n916_));
  NOR4_X1   g715(.A1(new_n828_), .A2(new_n916_), .A3(new_n641_), .A4(new_n373_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n917_), .A2(new_n633_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(new_n918_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g718(.A1(new_n917_), .A2(new_n624_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(G204gat), .ZN(G1353gat));
  NAND2_X1  g720(.A1(new_n917_), .A2(new_n860_), .ZN(new_n922_));
  NOR2_X1   g721(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n923_));
  AND2_X1   g722(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n924_));
  NOR3_X1   g723(.A1(new_n922_), .A2(new_n923_), .A3(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(new_n925_), .B1(new_n922_), .B2(new_n923_), .ZN(G1354gat));
  AOI21_X1  g725(.A(G218gat), .B1(new_n917_), .B2(new_n631_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n680_), .A2(G218gat), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n928_), .B(KEYINPUT127), .Z(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n917_), .B2(new_n929_), .ZN(G1355gat));
endmodule


