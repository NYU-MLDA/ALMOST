//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n862_, new_n863_, new_n865_, new_n866_, new_n867_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n877_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n929_,
    new_n930_, new_n931_, new_n932_, new_n933_, new_n935_, new_n936_,
    new_n937_, new_n938_, new_n939_, new_n941_, new_n942_, new_n943_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n951_, new_n952_;
  XOR2_X1   g000(.A(G1gat), .B(G8gat), .Z(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT75), .B(G15gat), .Z(new_n203_));
  NAND2_X1  g002(.A1(new_n203_), .A2(G22gat), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT75), .B(G15gat), .ZN(new_n205_));
  INV_X1    g004(.A(G22gat), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n204_), .A2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G1gat), .ZN(new_n209_));
  INV_X1    g008(.A(G8gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(KEYINPUT14), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n208_), .A2(new_n211_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n212_), .A2(KEYINPUT76), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n214_));
  NAND3_X1  g013(.A1(new_n208_), .A2(new_n214_), .A3(new_n211_), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n202_), .B1(new_n213_), .B2(new_n215_), .ZN(new_n216_));
  AOI21_X1  g015(.A(new_n214_), .B1(new_n208_), .B2(new_n211_), .ZN(new_n217_));
  INV_X1    g016(.A(new_n211_), .ZN(new_n218_));
  AOI211_X1 g017(.A(KEYINPUT76), .B(new_n218_), .C1(new_n204_), .C2(new_n207_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n202_), .ZN(new_n220_));
  NOR3_X1   g019(.A1(new_n217_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n216_), .A2(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(G231gat), .A2(G233gat), .ZN(new_n223_));
  AND2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NOR2_X1   g023(.A1(new_n222_), .A2(new_n223_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G71gat), .B(G78gat), .Z(new_n226_));
  XNOR2_X1  g025(.A(G57gat), .B(G64gat), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n226_), .B1(KEYINPUT11), .B2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n227_), .A2(new_n229_), .A3(KEYINPUT11), .ZN(new_n230_));
  INV_X1    g029(.A(new_n230_), .ZN(new_n231_));
  AOI21_X1  g030(.A(new_n229_), .B1(new_n227_), .B2(KEYINPUT11), .ZN(new_n232_));
  OAI21_X1  g031(.A(new_n228_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n227_), .A2(KEYINPUT11), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n234_), .A2(KEYINPUT68), .ZN(new_n235_));
  OR2_X1    g034(.A1(new_n227_), .A2(KEYINPUT11), .ZN(new_n236_));
  NAND4_X1  g035(.A1(new_n235_), .A2(new_n236_), .A3(new_n226_), .A4(new_n230_), .ZN(new_n237_));
  AOI21_X1  g036(.A(KEYINPUT69), .B1(new_n233_), .B2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  NAND3_X1  g038(.A1(new_n233_), .A2(new_n237_), .A3(KEYINPUT69), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  OR3_X1    g040(.A1(new_n224_), .A2(new_n225_), .A3(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n241_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G127gat), .B(G155gat), .Z(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT16), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G183gat), .B(G211gat), .ZN(new_n246_));
  XNOR2_X1  g045(.A(new_n245_), .B(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n247_), .B(KEYINPUT17), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n242_), .A2(new_n243_), .A3(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n233_), .A2(new_n237_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT77), .ZN(new_n251_));
  OR3_X1    g050(.A1(new_n224_), .A2(new_n225_), .A3(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n253_));
  NOR2_X1   g052(.A1(new_n247_), .A2(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n251_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n252_), .A2(new_n254_), .A3(new_n255_), .ZN(new_n256_));
  AND2_X1   g055(.A1(new_n249_), .A2(new_n256_), .ZN(new_n257_));
  XOR2_X1   g056(.A(G8gat), .B(G36gat), .Z(new_n258_));
  XNOR2_X1  g057(.A(KEYINPUT88), .B(KEYINPUT18), .ZN(new_n259_));
  XNOR2_X1  g058(.A(new_n258_), .B(new_n259_), .ZN(new_n260_));
  XNOR2_X1  g059(.A(G64gat), .B(G92gat), .ZN(new_n261_));
  XNOR2_X1  g060(.A(new_n260_), .B(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT21), .ZN(new_n264_));
  INV_X1    g063(.A(G204gat), .ZN(new_n265_));
  OAI21_X1  g064(.A(KEYINPUT85), .B1(new_n265_), .B2(G197gat), .ZN(new_n266_));
  AND2_X1   g065(.A1(KEYINPUT84), .A2(G204gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(KEYINPUT84), .A2(G204gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(new_n267_), .A2(new_n268_), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n266_), .B1(new_n269_), .B2(G197gat), .ZN(new_n270_));
  INV_X1    g069(.A(G197gat), .ZN(new_n271_));
  NOR4_X1   g070(.A1(new_n267_), .A2(new_n268_), .A3(KEYINPUT85), .A4(new_n271_), .ZN(new_n272_));
  OAI21_X1  g071(.A(new_n264_), .B1(new_n270_), .B2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274_));
  NOR3_X1   g073(.A1(new_n267_), .A2(new_n268_), .A3(G197gat), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n264_), .B1(G197gat), .B2(G204gat), .ZN(new_n276_));
  INV_X1    g075(.A(new_n276_), .ZN(new_n277_));
  OAI21_X1  g076(.A(new_n274_), .B1(new_n275_), .B2(new_n277_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n278_), .ZN(new_n279_));
  NOR2_X1   g078(.A1(new_n270_), .A2(new_n272_), .ZN(new_n280_));
  NOR2_X1   g079(.A1(new_n274_), .A2(new_n264_), .ZN(new_n281_));
  AOI22_X1  g080(.A1(new_n273_), .A2(new_n279_), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  NOR2_X1   g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283_));
  INV_X1    g082(.A(new_n283_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G169gat), .A2(G176gat), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n284_), .A2(KEYINPUT24), .A3(new_n285_), .ZN(new_n286_));
  INV_X1    g085(.A(G190gat), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n287_), .A2(KEYINPUT78), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT78), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(G190gat), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n288_), .A2(new_n290_), .A3(KEYINPUT26), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT26), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n292_), .A2(G190gat), .ZN(new_n293_));
  INV_X1    g092(.A(G183gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(KEYINPUT25), .ZN(new_n295_));
  INV_X1    g094(.A(KEYINPUT25), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(G183gat), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n293_), .A2(new_n295_), .A3(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n286_), .B1(new_n291_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT79), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  OAI211_X1 g100(.A(KEYINPUT79), .B(new_n286_), .C1(new_n291_), .C2(new_n298_), .ZN(new_n302_));
  NAND2_X1  g101(.A1(G183gat), .A2(G190gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT23), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND3_X1  g104(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  INV_X1    g106(.A(new_n307_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT24), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n283_), .A2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n308_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n301_), .A2(new_n302_), .A3(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n288_), .A2(new_n290_), .A3(new_n294_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n308_), .A2(new_n314_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n316_), .B(G169gat), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n315_), .A2(new_n317_), .ZN(new_n318_));
  NAND3_X1  g117(.A1(new_n282_), .A2(new_n313_), .A3(new_n318_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT20), .ZN(new_n320_));
  OR2_X1    g119(.A1(KEYINPUT84), .A2(G204gat), .ZN(new_n321_));
  NAND2_X1  g120(.A1(KEYINPUT84), .A2(G204gat), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n321_), .A2(G197gat), .A3(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(new_n266_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(KEYINPUT85), .ZN(new_n326_));
  NAND4_X1  g125(.A1(new_n321_), .A2(new_n326_), .A3(G197gat), .A4(new_n322_), .ZN(new_n327_));
  NAND3_X1  g126(.A1(new_n325_), .A2(new_n281_), .A3(new_n327_), .ZN(new_n328_));
  AOI21_X1  g127(.A(KEYINPUT21), .B1(new_n325_), .B2(new_n327_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n328_), .B1(new_n329_), .B2(new_n278_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n287_), .A2(KEYINPUT26), .ZN(new_n331_));
  NAND4_X1  g130(.A1(new_n293_), .A2(new_n295_), .A3(new_n297_), .A4(new_n331_), .ZN(new_n332_));
  NAND4_X1  g131(.A1(new_n308_), .A2(new_n332_), .A3(new_n286_), .A4(new_n310_), .ZN(new_n333_));
  OAI211_X1 g132(.A(new_n305_), .B(new_n306_), .C1(G183gat), .C2(G190gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n317_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n333_), .A2(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n320_), .B1(new_n330_), .B2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n319_), .A2(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n339_), .B(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n338_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n313_), .A2(new_n318_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n344_), .A2(new_n330_), .ZN(new_n345_));
  AND2_X1   g144(.A1(new_n333_), .A2(new_n335_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n320_), .B1(new_n282_), .B2(new_n346_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n345_), .A2(new_n341_), .A3(new_n347_), .ZN(new_n348_));
  NAND3_X1  g147(.A1(new_n343_), .A2(new_n348_), .A3(KEYINPUT87), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT87), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n345_), .A2(new_n350_), .A3(new_n347_), .A4(new_n341_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n263_), .B1(new_n349_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(new_n263_), .A3(new_n351_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT27), .B1(new_n353_), .B2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT27), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n273_), .A2(new_n279_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n346_), .A2(new_n357_), .A3(new_n328_), .ZN(new_n358_));
  AOI21_X1  g157(.A(new_n311_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n359_));
  AOI22_X1  g158(.A1(new_n359_), .A2(new_n302_), .B1(new_n317_), .B2(new_n315_), .ZN(new_n360_));
  OAI211_X1 g159(.A(new_n358_), .B(KEYINPUT20), .C1(new_n360_), .C2(new_n282_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT87), .B1(new_n361_), .B2(new_n342_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n341_), .B1(new_n319_), .B2(new_n337_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n351_), .B1(new_n362_), .B2(new_n363_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n356_), .B1(new_n364_), .B2(new_n262_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n319_), .A2(new_n341_), .A3(new_n337_), .ZN(new_n366_));
  INV_X1    g165(.A(KEYINPUT91), .ZN(new_n367_));
  NAND2_X1  g166(.A1(new_n366_), .A2(new_n367_), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n319_), .A2(new_n337_), .A3(KEYINPUT91), .A4(new_n341_), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n282_), .B1(new_n318_), .B2(new_n313_), .ZN(new_n370_));
  OAI21_X1  g169(.A(KEYINPUT20), .B1(new_n330_), .B2(new_n336_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n342_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n368_), .A2(new_n369_), .A3(new_n372_), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n373_), .A2(new_n263_), .ZN(new_n374_));
  INV_X1    g173(.A(KEYINPUT92), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n373_), .A2(KEYINPUT92), .A3(new_n263_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n365_), .A2(new_n376_), .A3(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n378_), .A2(KEYINPUT93), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT93), .ZN(new_n380_));
  NAND4_X1  g179(.A1(new_n365_), .A2(new_n376_), .A3(new_n380_), .A4(new_n377_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n355_), .B1(new_n379_), .B2(new_n381_), .ZN(new_n382_));
  XNOR2_X1  g181(.A(G78gat), .B(G106gat), .ZN(new_n383_));
  INV_X1    g182(.A(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G155gat), .A2(G162gat), .ZN(new_n385_));
  INV_X1    g184(.A(new_n385_), .ZN(new_n386_));
  NOR2_X1   g185(.A1(G155gat), .A2(G162gat), .ZN(new_n387_));
  NOR2_X1   g186(.A1(new_n386_), .A2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n390_));
  XNOR2_X1  g189(.A(new_n390_), .B(KEYINPUT81), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT3), .ZN(new_n392_));
  INV_X1    g191(.A(G141gat), .ZN(new_n393_));
  INV_X1    g192(.A(G148gat), .ZN(new_n394_));
  NAND3_X1  g193(.A1(new_n392_), .A2(new_n393_), .A3(new_n394_), .ZN(new_n395_));
  OAI21_X1  g194(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n396_));
  NAND3_X1  g195(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n397_));
  AND3_X1   g196(.A1(new_n395_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n389_), .B1(new_n391_), .B2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n393_), .A2(new_n394_), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G141gat), .A2(G148gat), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n387_), .B1(KEYINPUT1), .B2(new_n385_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n385_), .A2(KEYINPUT1), .ZN(new_n404_));
  AOI21_X1  g203(.A(new_n402_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT29), .B1(new_n399_), .B2(new_n405_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(KEYINPUT83), .A2(G233gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NOR2_X1   g207(.A1(KEYINPUT83), .A2(G233gat), .ZN(new_n409_));
  OAI21_X1  g208(.A(G228gat), .B1(new_n408_), .B2(new_n409_), .ZN(new_n410_));
  AND3_X1   g209(.A1(new_n406_), .A2(new_n330_), .A3(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n410_), .B1(new_n406_), .B2(new_n330_), .ZN(new_n412_));
  OAI21_X1  g211(.A(new_n384_), .B1(new_n411_), .B2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n410_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT29), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT81), .ZN(new_n416_));
  XNOR2_X1  g215(.A(new_n390_), .B(new_n416_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n395_), .A2(new_n396_), .A3(new_n397_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n388_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n405_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n415_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  OAI21_X1  g220(.A(new_n414_), .B1(new_n282_), .B2(new_n421_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n406_), .A2(new_n330_), .A3(new_n410_), .ZN(new_n423_));
  NAND3_X1  g222(.A1(new_n422_), .A2(new_n383_), .A3(new_n423_), .ZN(new_n424_));
  NAND3_X1  g223(.A1(new_n413_), .A2(new_n424_), .A3(KEYINPUT82), .ZN(new_n425_));
  NAND3_X1  g224(.A1(new_n419_), .A2(new_n415_), .A3(new_n420_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n426_), .B(KEYINPUT28), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n425_), .A2(new_n428_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(G22gat), .B(G50gat), .ZN(new_n430_));
  NAND4_X1  g229(.A1(new_n413_), .A2(new_n424_), .A3(KEYINPUT82), .A4(new_n427_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n429_), .A2(new_n430_), .A3(new_n431_), .ZN(new_n432_));
  AOI21_X1  g231(.A(new_n430_), .B1(new_n429_), .B2(new_n431_), .ZN(new_n433_));
  NOR2_X1   g232(.A1(new_n432_), .A2(new_n433_), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G71gat), .B(G99gat), .ZN(new_n435_));
  INV_X1    g234(.A(G43gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n360_), .B(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(KEYINPUT80), .B(KEYINPUT31), .Z(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G127gat), .B(G134gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(G113gat), .B(G120gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n441_), .B(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  NAND2_X1  g243(.A1(G227gat), .A2(G233gat), .ZN(new_n445_));
  INV_X1    g244(.A(G15gat), .ZN(new_n446_));
  XNOR2_X1  g245(.A(new_n445_), .B(new_n446_), .ZN(new_n447_));
  XNOR2_X1  g246(.A(new_n447_), .B(KEYINPUT30), .ZN(new_n448_));
  XNOR2_X1  g247(.A(new_n444_), .B(new_n448_), .ZN(new_n449_));
  XNOR2_X1  g248(.A(new_n440_), .B(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G225gat), .A2(G233gat), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n419_), .A2(new_n420_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n444_), .ZN(new_n454_));
  NAND3_X1  g253(.A1(new_n419_), .A2(new_n420_), .A3(new_n443_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n452_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n454_), .A2(KEYINPUT4), .A3(new_n455_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT4), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n453_), .A2(new_n458_), .A3(new_n444_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT89), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT89), .ZN(new_n461_));
  NAND4_X1  g260(.A1(new_n453_), .A2(new_n461_), .A3(new_n458_), .A4(new_n444_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n457_), .A2(new_n460_), .A3(new_n462_), .ZN(new_n463_));
  AOI21_X1  g262(.A(new_n456_), .B1(new_n463_), .B2(new_n452_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G1gat), .B(G29gat), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n465_), .B(G85gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(KEYINPUT0), .B(G57gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n464_), .B(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n450_), .A2(new_n469_), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n382_), .A2(new_n434_), .A3(new_n470_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n379_), .A2(new_n381_), .ZN(new_n472_));
  AND2_X1   g271(.A1(new_n464_), .A2(new_n468_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n463_), .A2(new_n452_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n456_), .ZN(new_n475_));
  AOI21_X1  g274(.A(new_n468_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  NOR2_X1   g275(.A1(new_n473_), .A2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n477_), .B1(new_n432_), .B2(new_n433_), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n478_), .A2(new_n355_), .ZN(new_n479_));
  INV_X1    g278(.A(KEYINPUT32), .ZN(new_n480_));
  OAI21_X1  g279(.A(new_n364_), .B1(new_n480_), .B2(new_n263_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n373_), .A2(KEYINPUT32), .A3(new_n262_), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n469_), .A2(new_n481_), .A3(new_n482_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n476_), .A2(KEYINPUT33), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n454_), .A2(new_n452_), .A3(new_n455_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n468_), .B(new_n485_), .C1(new_n463_), .C2(new_n452_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n353_), .A2(new_n484_), .A3(new_n354_), .A4(new_n486_), .ZN(new_n487_));
  OAI21_X1  g286(.A(KEYINPUT90), .B1(new_n476_), .B2(KEYINPUT33), .ZN(new_n488_));
  INV_X1    g287(.A(KEYINPUT90), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT33), .ZN(new_n490_));
  OAI211_X1 g289(.A(new_n489_), .B(new_n490_), .C1(new_n464_), .C2(new_n468_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n488_), .A2(new_n491_), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n483_), .B1(new_n487_), .B2(new_n492_), .ZN(new_n493_));
  AOI22_X1  g292(.A1(new_n472_), .A2(new_n479_), .B1(new_n493_), .B2(new_n434_), .ZN(new_n494_));
  INV_X1    g293(.A(new_n450_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n471_), .B1(new_n494_), .B2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G229gat), .A2(G233gat), .ZN(new_n497_));
  INV_X1    g296(.A(new_n497_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n213_), .A2(new_n202_), .A3(new_n215_), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n220_), .B1(new_n217_), .B2(new_n219_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G29gat), .B(G36gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(G43gat), .B(G50gat), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n501_), .B(new_n502_), .ZN(new_n503_));
  AND3_X1   g302(.A1(new_n499_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n503_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n505_));
  OAI21_X1  g304(.A(new_n498_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n499_), .A2(new_n500_), .A3(new_n503_), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n503_), .B(KEYINPUT15), .ZN(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  OAI211_X1 g308(.A(new_n507_), .B(new_n497_), .C1(new_n222_), .C2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n506_), .A2(new_n510_), .ZN(new_n511_));
  XNOR2_X1  g310(.A(G113gat), .B(G141gat), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G169gat), .B(G197gat), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n512_), .B(new_n513_), .Z(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n511_), .A2(new_n515_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n506_), .A2(new_n510_), .A3(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n496_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(G230gat), .A2(G233gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(KEYINPUT64), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  XOR2_X1   g321(.A(G85gat), .B(G92gat), .Z(new_n523_));
  INV_X1    g322(.A(G99gat), .ZN(new_n524_));
  INV_X1    g323(.A(G106gat), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n524_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT7), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n527_), .A2(KEYINPUT66), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(KEYINPUT66), .B(KEYINPUT7), .ZN(new_n530_));
  OAI21_X1  g329(.A(new_n529_), .B1(new_n530_), .B2(new_n526_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G99gat), .A2(G106gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n532_), .A2(KEYINPUT6), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT6), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n534_), .A2(G99gat), .A3(G106gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n533_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(new_n536_), .ZN(new_n537_));
  OAI21_X1  g336(.A(new_n523_), .B1(new_n531_), .B2(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT67), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(new_n539_), .A3(KEYINPUT8), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  AOI21_X1  g340(.A(new_n539_), .B1(new_n538_), .B2(KEYINPUT8), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n536_), .B(KEYINPUT65), .ZN(new_n543_));
  NOR2_X1   g342(.A1(new_n543_), .A2(new_n531_), .ZN(new_n544_));
  INV_X1    g343(.A(KEYINPUT8), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n523_), .A2(new_n545_), .ZN(new_n546_));
  OAI22_X1  g345(.A1(new_n541_), .A2(new_n542_), .B1(new_n544_), .B2(new_n546_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(KEYINPUT10), .B(G99gat), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n548_), .A2(G106gat), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT9), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n550_), .A2(G85gat), .A3(G92gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n523_), .A2(KEYINPUT9), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n549_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT65), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n536_), .B(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND4_X1  g356(.A1(new_n547_), .A2(new_n240_), .A3(new_n557_), .A4(new_n239_), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n547_), .A2(new_n557_), .B1(new_n240_), .B2(new_n239_), .ZN(new_n560_));
  OAI21_X1  g359(.A(new_n522_), .B1(new_n559_), .B2(new_n560_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n531_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n546_), .B1(new_n556_), .B2(new_n562_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n538_), .A2(KEYINPUT8), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT67), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n563_), .B1(new_n565_), .B2(new_n540_), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT70), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n554_), .A2(new_n556_), .A3(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(KEYINPUT70), .B1(new_n553_), .B2(new_n543_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n568_), .A2(new_n569_), .ZN(new_n570_));
  OAI211_X1 g369(.A(KEYINPUT12), .B(new_n250_), .C1(new_n566_), .C2(new_n570_), .ZN(new_n571_));
  XNOR2_X1  g370(.A(KEYINPUT71), .B(KEYINPUT12), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  OAI211_X1 g372(.A(new_n558_), .B(new_n571_), .C1(new_n560_), .C2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n561_), .B1(new_n574_), .B2(new_n522_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G120gat), .B(G148gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT5), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G176gat), .B(G204gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n577_), .B(new_n578_), .Z(new_n579_));
  NAND2_X1  g378(.A1(new_n575_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n579_), .ZN(new_n581_));
  OAI211_X1 g380(.A(new_n561_), .B(new_n581_), .C1(new_n574_), .C2(new_n522_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(KEYINPUT13), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NOR2_X1   g385(.A1(new_n583_), .A2(new_n584_), .ZN(new_n587_));
  NOR2_X1   g386(.A1(new_n586_), .A2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT37), .ZN(new_n589_));
  OAI21_X1  g388(.A(new_n508_), .B1(new_n566_), .B2(new_n570_), .ZN(new_n590_));
  NAND3_X1  g389(.A1(new_n547_), .A2(new_n503_), .A3(new_n557_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT73), .ZN(new_n592_));
  NAND2_X1  g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  XNOR2_X1  g392(.A(new_n593_), .B(KEYINPUT34), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT35), .Z(new_n595_));
  NAND4_X1  g394(.A1(new_n590_), .A2(new_n591_), .A3(new_n592_), .A4(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n590_), .A2(new_n591_), .A3(new_n595_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n597_), .A2(KEYINPUT73), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n594_), .A2(KEYINPUT35), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n599_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n600_));
  OAI211_X1 g399(.A(KEYINPUT36), .B(new_n596_), .C1(new_n598_), .C2(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G190gat), .B(G218gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT72), .ZN(new_n603_));
  XOR2_X1   g402(.A(G134gat), .B(G162gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n601_), .A2(new_n605_), .ZN(new_n606_));
  AND2_X1   g405(.A1(new_n590_), .A2(new_n591_), .ZN(new_n607_));
  OAI211_X1 g406(.A(KEYINPUT73), .B(new_n597_), .C1(new_n607_), .C2(new_n599_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(KEYINPUT74), .A3(new_n596_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n605_), .A2(new_n610_), .ZN(new_n611_));
  AND3_X1   g410(.A1(new_n606_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n612_));
  AOI21_X1  g411(.A(new_n609_), .B1(new_n606_), .B2(new_n611_), .ZN(new_n613_));
  OAI21_X1  g412(.A(new_n589_), .B1(new_n612_), .B2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n606_), .A2(new_n611_), .ZN(new_n615_));
  INV_X1    g414(.A(new_n609_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND3_X1  g416(.A1(new_n606_), .A2(new_n609_), .A3(new_n611_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n617_), .A2(KEYINPUT37), .A3(new_n618_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n614_), .A2(new_n619_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n620_), .ZN(new_n621_));
  AND4_X1   g420(.A1(new_n257_), .A2(new_n519_), .A3(new_n588_), .A4(new_n621_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n622_), .A2(new_n209_), .A3(new_n469_), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n623_), .B(KEYINPUT38), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n612_), .A2(new_n613_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  AND2_X1   g425(.A1(new_n496_), .A2(new_n626_), .ZN(new_n627_));
  NAND4_X1  g426(.A1(new_n627_), .A2(new_n257_), .A3(new_n518_), .A4(new_n588_), .ZN(new_n628_));
  XOR2_X1   g427(.A(new_n628_), .B(KEYINPUT94), .Z(new_n629_));
  AND2_X1   g428(.A1(new_n629_), .A2(new_n469_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n624_), .B1(new_n630_), .B2(new_n209_), .ZN(G1324gat));
  OR2_X1    g430(.A1(new_n628_), .A2(new_n382_), .ZN(new_n632_));
  AND2_X1   g431(.A1(new_n632_), .A2(KEYINPUT96), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n632_), .A2(KEYINPUT96), .ZN(new_n634_));
  NOR3_X1   g433(.A1(new_n633_), .A2(new_n634_), .A3(new_n210_), .ZN(new_n635_));
  OR2_X1    g434(.A1(KEYINPUT97), .A2(KEYINPUT39), .ZN(new_n636_));
  NAND2_X1  g435(.A1(KEYINPUT97), .A2(KEYINPUT39), .ZN(new_n637_));
  NAND3_X1  g436(.A1(new_n635_), .A2(new_n636_), .A3(new_n637_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n382_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n622_), .A2(new_n210_), .A3(new_n639_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT95), .Z(new_n641_));
  OAI211_X1 g440(.A(new_n638_), .B(new_n641_), .C1(new_n635_), .C2(new_n636_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT40), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  OR2_X1    g443(.A1(new_n635_), .A2(new_n636_), .ZN(new_n645_));
  NAND4_X1  g444(.A1(new_n645_), .A2(KEYINPUT40), .A3(new_n638_), .A4(new_n641_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(G1325gat));
  AOI21_X1  g446(.A(new_n446_), .B1(new_n629_), .B2(new_n495_), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n648_), .B(KEYINPUT41), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n622_), .A2(new_n446_), .A3(new_n495_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n649_), .A2(new_n650_), .ZN(G1326gat));
  INV_X1    g450(.A(new_n434_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n206_), .B1(new_n629_), .B2(new_n652_), .ZN(new_n653_));
  XOR2_X1   g452(.A(new_n653_), .B(KEYINPUT42), .Z(new_n654_));
  NAND3_X1  g453(.A1(new_n622_), .A2(new_n206_), .A3(new_n652_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1327gat));
  INV_X1    g455(.A(new_n588_), .ZN(new_n657_));
  NOR3_X1   g456(.A1(new_n657_), .A2(new_n626_), .A3(new_n257_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n519_), .A2(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(G29gat), .B1(new_n660_), .B2(new_n469_), .ZN(new_n661_));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n662_));
  INV_X1    g461(.A(new_n257_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n588_), .A2(new_n663_), .A3(new_n518_), .ZN(new_n664_));
  AOI21_X1  g463(.A(KEYINPUT92), .B1(new_n373_), .B2(new_n263_), .ZN(new_n665_));
  NOR3_X1   g464(.A1(new_n665_), .A2(new_n352_), .A3(new_n356_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n380_), .B1(new_n666_), .B2(new_n377_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n381_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n479_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n493_), .A2(new_n434_), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n495_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n355_), .ZN(new_n672_));
  AND4_X1   g471(.A1(new_n434_), .A2(new_n472_), .A3(new_n672_), .A4(new_n470_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n620_), .B1(new_n671_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT43), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT43), .ZN(new_n676_));
  NAND3_X1  g475(.A1(new_n496_), .A2(new_n676_), .A3(new_n620_), .ZN(new_n677_));
  AOI21_X1  g476(.A(new_n664_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n678_));
  OAI21_X1  g477(.A(new_n662_), .B1(new_n678_), .B2(KEYINPUT44), .ZN(new_n679_));
  INV_X1    g478(.A(new_n664_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n496_), .A2(new_n676_), .A3(new_n620_), .ZN(new_n681_));
  AOI21_X1  g480(.A(new_n676_), .B1(new_n496_), .B2(new_n620_), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n680_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n683_), .A2(KEYINPUT98), .A3(new_n684_), .ZN(new_n685_));
  NAND2_X1  g484(.A1(new_n679_), .A2(new_n685_), .ZN(new_n686_));
  OAI211_X1 g485(.A(KEYINPUT44), .B(new_n680_), .C1(new_n681_), .C2(new_n682_), .ZN(new_n687_));
  AND2_X1   g486(.A1(new_n686_), .A2(new_n687_), .ZN(new_n688_));
  AND2_X1   g487(.A1(new_n469_), .A2(G29gat), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n661_), .B1(new_n688_), .B2(new_n689_), .ZN(G1328gat));
  INV_X1    g489(.A(G36gat), .ZN(new_n691_));
  NAND3_X1  g490(.A1(new_n660_), .A2(new_n691_), .A3(new_n639_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT45), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n382_), .B1(new_n678_), .B2(KEYINPUT44), .ZN(new_n694_));
  NOR3_X1   g493(.A1(new_n678_), .A2(new_n662_), .A3(KEYINPUT44), .ZN(new_n695_));
  AOI21_X1  g494(.A(KEYINPUT98), .B1(new_n683_), .B2(new_n684_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n694_), .B(KEYINPUT99), .C1(new_n695_), .C2(new_n696_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n697_), .A2(G36gat), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT99), .B1(new_n686_), .B2(new_n694_), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT100), .ZN(new_n700_));
  NOR3_X1   g499(.A1(new_n698_), .A2(new_n699_), .A3(new_n700_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n687_), .A2(new_n639_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n702_), .B1(new_n679_), .B2(new_n685_), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n691_), .B1(new_n703_), .B2(KEYINPUT99), .ZN(new_n704_));
  OAI21_X1  g503(.A(new_n694_), .B1(new_n695_), .B2(new_n696_), .ZN(new_n705_));
  INV_X1    g504(.A(KEYINPUT99), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n705_), .A2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(KEYINPUT100), .B1(new_n704_), .B2(new_n707_), .ZN(new_n708_));
  OAI21_X1  g507(.A(new_n693_), .B1(new_n701_), .B2(new_n708_), .ZN(new_n709_));
  NOR2_X1   g508(.A1(KEYINPUT101), .A2(KEYINPUT46), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(new_n711_));
  OAI221_X1 g510(.A(new_n693_), .B1(KEYINPUT101), .B2(KEYINPUT46), .C1(new_n701_), .C2(new_n708_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1329gat));
  NAND4_X1  g512(.A1(new_n686_), .A2(G43gat), .A3(new_n495_), .A4(new_n687_), .ZN(new_n714_));
  OR2_X1    g513(.A1(new_n714_), .A2(KEYINPUT102), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n436_), .B1(new_n659_), .B2(new_n450_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n714_), .A2(KEYINPUT102), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n715_), .A2(new_n716_), .A3(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n718_), .B(new_n720_), .ZN(G1330gat));
  AOI21_X1  g520(.A(G50gat), .B1(new_n660_), .B2(new_n652_), .ZN(new_n722_));
  AND2_X1   g521(.A1(new_n652_), .A2(G50gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n722_), .B1(new_n688_), .B2(new_n723_), .ZN(G1331gat));
  INV_X1    g523(.A(new_n518_), .ZN(new_n725_));
  AND2_X1   g524(.A1(new_n496_), .A2(new_n725_), .ZN(new_n726_));
  AND4_X1   g525(.A1(new_n257_), .A2(new_n726_), .A3(new_n657_), .A4(new_n621_), .ZN(new_n727_));
  AOI21_X1  g526(.A(G57gat), .B1(new_n727_), .B2(new_n469_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT104), .ZN(new_n729_));
  AND4_X1   g528(.A1(new_n627_), .A2(new_n257_), .A3(new_n725_), .A4(new_n657_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n469_), .A2(G57gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n729_), .B1(new_n730_), .B2(new_n731_), .ZN(G1332gat));
  INV_X1    g531(.A(G64gat), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n733_), .B1(new_n730_), .B2(new_n639_), .ZN(new_n734_));
  XOR2_X1   g533(.A(new_n734_), .B(KEYINPUT48), .Z(new_n735_));
  NAND3_X1  g534(.A1(new_n727_), .A2(new_n733_), .A3(new_n639_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(G1333gat));
  INV_X1    g536(.A(G71gat), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n738_), .B1(new_n730_), .B2(new_n495_), .ZN(new_n739_));
  XOR2_X1   g538(.A(new_n739_), .B(KEYINPUT49), .Z(new_n740_));
  NAND3_X1  g539(.A1(new_n727_), .A2(new_n738_), .A3(new_n495_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1334gat));
  INV_X1    g541(.A(G78gat), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n730_), .B2(new_n652_), .ZN(new_n744_));
  XOR2_X1   g543(.A(KEYINPUT105), .B(KEYINPUT50), .Z(new_n745_));
  XNOR2_X1  g544(.A(new_n744_), .B(new_n745_), .ZN(new_n746_));
  NAND3_X1  g545(.A1(new_n727_), .A2(new_n743_), .A3(new_n652_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1335gat));
  AND4_X1   g547(.A1(new_n625_), .A2(new_n726_), .A3(new_n663_), .A4(new_n657_), .ZN(new_n749_));
  AOI21_X1  g548(.A(G85gat), .B1(new_n749_), .B2(new_n469_), .ZN(new_n750_));
  XOR2_X1   g549(.A(new_n750_), .B(KEYINPUT106), .Z(new_n751_));
  NAND3_X1  g550(.A1(new_n657_), .A2(new_n663_), .A3(new_n725_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n675_), .B2(new_n677_), .ZN(new_n753_));
  AND2_X1   g552(.A1(new_n469_), .A2(G85gat), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n751_), .B1(new_n753_), .B2(new_n754_), .ZN(G1336gat));
  AOI21_X1  g554(.A(G92gat), .B1(new_n749_), .B2(new_n639_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n639_), .A2(G92gat), .ZN(new_n757_));
  XOR2_X1   g556(.A(new_n757_), .B(KEYINPUT107), .Z(new_n758_));
  AOI21_X1  g557(.A(new_n756_), .B1(new_n753_), .B2(new_n758_), .ZN(G1337gat));
  AOI21_X1  g558(.A(new_n524_), .B1(new_n753_), .B2(new_n495_), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n450_), .A2(new_n548_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n749_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n763_));
  XNOR2_X1  g562(.A(new_n762_), .B(new_n763_), .ZN(G1338gat));
  NAND3_X1  g563(.A1(new_n749_), .A2(new_n525_), .A3(new_n652_), .ZN(new_n765_));
  XOR2_X1   g564(.A(new_n765_), .B(KEYINPUT109), .Z(new_n766_));
  AOI21_X1  g565(.A(new_n525_), .B1(new_n753_), .B2(new_n652_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n767_), .A2(KEYINPUT52), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(KEYINPUT52), .ZN(new_n769_));
  NAND3_X1  g568(.A1(new_n766_), .A2(new_n768_), .A3(new_n769_), .ZN(new_n770_));
  XNOR2_X1  g569(.A(new_n770_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND2_X1  g570(.A1(new_n257_), .A2(new_n725_), .ZN(new_n772_));
  XNOR2_X1  g571(.A(new_n772_), .B(KEYINPUT110), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n621_), .A2(new_n588_), .A3(new_n773_), .ZN(new_n774_));
  XNOR2_X1  g573(.A(new_n774_), .B(KEYINPUT54), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT57), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT55), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n777_), .B1(new_n574_), .B2(new_n522_), .ZN(new_n778_));
  AND2_X1   g577(.A1(new_n571_), .A2(new_n558_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n547_), .A2(new_n557_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n241_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n781_), .A2(new_n572_), .ZN(new_n782_));
  NAND4_X1  g581(.A1(new_n779_), .A2(new_n782_), .A3(KEYINPUT55), .A4(new_n521_), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n574_), .A2(new_n522_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n778_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n579_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(KEYINPUT56), .A3(new_n579_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n518_), .A2(new_n582_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT111), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n518_), .A2(new_n582_), .A3(new_n793_), .ZN(new_n794_));
  AND2_X1   g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n517_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n507_), .A2(new_n498_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n509_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n798_));
  NOR2_X1   g597(.A1(new_n797_), .A2(new_n798_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n497_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n800_), .A2(new_n515_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n799_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(KEYINPUT112), .A3(new_n515_), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n796_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  AOI22_X1  g604(.A1(new_n790_), .A2(new_n795_), .B1(new_n583_), .B2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(new_n776_), .B1(new_n806_), .B2(new_n625_), .ZN(new_n807_));
  AND3_X1   g606(.A1(new_n785_), .A2(KEYINPUT56), .A3(new_n579_), .ZN(new_n808_));
  AOI21_X1  g607(.A(KEYINPUT56), .B1(new_n785_), .B2(new_n579_), .ZN(new_n809_));
  INV_X1    g608(.A(KEYINPUT113), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n810_), .B1(new_n805_), .B2(new_n582_), .ZN(new_n811_));
  INV_X1    g610(.A(new_n503_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n216_), .B2(new_n221_), .ZN(new_n813_));
  AOI21_X1  g612(.A(new_n498_), .B1(new_n813_), .B2(new_n507_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n802_), .B1(new_n814_), .B2(new_n514_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n799_), .ZN(new_n816_));
  NAND3_X1  g615(.A1(new_n815_), .A2(new_n804_), .A3(new_n816_), .ZN(new_n817_));
  AND4_X1   g616(.A1(new_n810_), .A2(new_n582_), .A3(new_n817_), .A4(new_n517_), .ZN(new_n818_));
  OAI22_X1  g617(.A1(new_n808_), .A2(new_n809_), .B1(new_n811_), .B2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n819_), .A2(new_n820_), .ZN(new_n821_));
  OAI211_X1 g620(.A(new_n790_), .B(KEYINPUT58), .C1(new_n811_), .C2(new_n818_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n620_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n807_), .A2(new_n823_), .ZN(new_n824_));
  OAI211_X1 g623(.A(new_n792_), .B(new_n794_), .C1(new_n808_), .C2(new_n809_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n583_), .A2(new_n805_), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n625_), .B1(new_n825_), .B2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n827_), .A2(KEYINPUT57), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n827_), .A2(KEYINPUT114), .A3(KEYINPUT57), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n824_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n775_), .B1(new_n832_), .B2(new_n257_), .ZN(new_n833_));
  NOR2_X1   g632(.A1(new_n639_), .A2(new_n652_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n834_), .A2(new_n469_), .A3(new_n495_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n833_), .A2(new_n836_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(G113gat), .B1(new_n838_), .B2(new_n518_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(KEYINPUT115), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n841_));
  XNOR2_X1  g640(.A(new_n774_), .B(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n830_), .A2(new_n831_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n824_), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n257_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n845_), .A2(KEYINPUT116), .ZN(new_n846_));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847_));
  OAI21_X1  g646(.A(new_n847_), .B1(new_n832_), .B2(new_n257_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n842_), .B1(new_n846_), .B2(new_n848_), .ZN(new_n849_));
  OR3_X1    g648(.A1(new_n849_), .A2(KEYINPUT59), .A3(new_n835_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n837_), .A2(KEYINPUT59), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  INV_X1    g651(.A(new_n852_), .ZN(new_n853_));
  XOR2_X1   g652(.A(KEYINPUT117), .B(G113gat), .Z(new_n854_));
  NOR2_X1   g653(.A1(new_n725_), .A2(new_n854_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n840_), .B1(new_n853_), .B2(new_n855_), .ZN(G1340gat));
  OAI21_X1  g655(.A(G120gat), .B1(new_n852_), .B2(new_n588_), .ZN(new_n857_));
  INV_X1    g656(.A(G120gat), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n858_), .B1(new_n588_), .B2(KEYINPUT60), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n859_), .B1(KEYINPUT60), .B2(new_n858_), .ZN(new_n860_));
  OAI21_X1  g659(.A(new_n857_), .B1(new_n837_), .B2(new_n860_), .ZN(G1341gat));
  OAI21_X1  g660(.A(G127gat), .B1(new_n852_), .B2(new_n663_), .ZN(new_n862_));
  OR2_X1    g661(.A1(new_n663_), .A2(G127gat), .ZN(new_n863_));
  OAI21_X1  g662(.A(new_n862_), .B1(new_n837_), .B2(new_n863_), .ZN(G1342gat));
  AOI21_X1  g663(.A(G134gat), .B1(new_n838_), .B2(new_n625_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT118), .B(G134gat), .ZN(new_n866_));
  NOR2_X1   g665(.A1(new_n621_), .A2(new_n866_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n865_), .B1(new_n853_), .B2(new_n867_), .ZN(G1343gat));
  NOR3_X1   g667(.A1(new_n639_), .A2(new_n477_), .A3(new_n434_), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n450_), .B(new_n869_), .C1(new_n845_), .C2(new_n842_), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n871_));
  NAND2_X1  g670(.A1(new_n870_), .A2(new_n871_), .ZN(new_n872_));
  NAND4_X1  g671(.A1(new_n833_), .A2(KEYINPUT119), .A3(new_n450_), .A4(new_n869_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n872_), .A2(new_n873_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n874_), .A2(new_n518_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n657_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(new_n877_), .B(G148gat), .ZN(G1345gat));
  XNOR2_X1  g677(.A(KEYINPUT61), .B(G155gat), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880_));
  AOI21_X1  g679(.A(new_n880_), .B1(new_n874_), .B2(new_n257_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n881_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n874_), .A2(new_n880_), .A3(new_n257_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n879_), .B1(new_n882_), .B2(new_n883_), .ZN(new_n884_));
  AOI211_X1 g683(.A(KEYINPUT120), .B(new_n663_), .C1(new_n872_), .C2(new_n873_), .ZN(new_n885_));
  INV_X1    g684(.A(new_n879_), .ZN(new_n886_));
  NOR3_X1   g685(.A1(new_n881_), .A2(new_n885_), .A3(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(new_n884_), .A2(new_n887_), .ZN(G1346gat));
  AND3_X1   g687(.A1(new_n874_), .A2(G162gat), .A3(new_n620_), .ZN(new_n889_));
  AOI21_X1  g688(.A(G162gat), .B1(new_n874_), .B2(new_n625_), .ZN(new_n890_));
  OR2_X1    g689(.A1(new_n890_), .A2(KEYINPUT121), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(KEYINPUT121), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n889_), .B1(new_n891_), .B2(new_n892_), .ZN(G1347gat));
  INV_X1    g692(.A(KEYINPUT62), .ZN(new_n894_));
  NOR3_X1   g693(.A1(new_n832_), .A2(new_n847_), .A3(new_n257_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n831_), .ZN(new_n896_));
  AOI21_X1  g695(.A(KEYINPUT114), .B1(new_n827_), .B2(KEYINPUT57), .ZN(new_n897_));
  OAI211_X1 g696(.A(new_n807_), .B(new_n823_), .C1(new_n896_), .C2(new_n897_), .ZN(new_n898_));
  AOI21_X1  g697(.A(KEYINPUT116), .B1(new_n898_), .B2(new_n663_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n775_), .B1(new_n895_), .B2(new_n899_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n382_), .A2(new_n469_), .A3(new_n450_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n518_), .ZN(new_n902_));
  XNOR2_X1  g701(.A(new_n902_), .B(KEYINPUT122), .ZN(new_n903_));
  NOR2_X1   g702(.A1(new_n903_), .A2(new_n652_), .ZN(new_n904_));
  NAND3_X1  g703(.A1(new_n900_), .A2(KEYINPUT123), .A3(new_n904_), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n905_), .A2(G169gat), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907_));
  INV_X1    g706(.A(new_n904_), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n907_), .B1(new_n849_), .B2(new_n908_), .ZN(new_n909_));
  AOI21_X1  g708(.A(new_n894_), .B1(new_n906_), .B2(new_n909_), .ZN(new_n910_));
  AND4_X1   g709(.A1(new_n894_), .A2(new_n909_), .A3(G169gat), .A4(new_n905_), .ZN(new_n911_));
  INV_X1    g710(.A(new_n901_), .ZN(new_n912_));
  NOR2_X1   g711(.A1(new_n912_), .A2(new_n652_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  OAI21_X1  g713(.A(KEYINPUT124), .B1(new_n849_), .B2(new_n914_), .ZN(new_n915_));
  INV_X1    g714(.A(KEYINPUT124), .ZN(new_n916_));
  NAND3_X1  g715(.A1(new_n900_), .A2(new_n916_), .A3(new_n913_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n915_), .A2(new_n917_), .ZN(new_n918_));
  XNOR2_X1  g717(.A(KEYINPUT22), .B(G169gat), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n518_), .A2(new_n919_), .ZN(new_n920_));
  XOR2_X1   g719(.A(new_n920_), .B(KEYINPUT125), .Z(new_n921_));
  OAI22_X1  g720(.A1(new_n910_), .A2(new_n911_), .B1(new_n918_), .B2(new_n921_), .ZN(G1348gat));
  INV_X1    g721(.A(new_n918_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(new_n657_), .ZN(new_n924_));
  INV_X1    g723(.A(G176gat), .ZN(new_n925_));
  AND2_X1   g724(.A1(new_n833_), .A2(new_n434_), .ZN(new_n926_));
  NOR3_X1   g725(.A1(new_n912_), .A2(new_n925_), .A3(new_n588_), .ZN(new_n927_));
  AOI22_X1  g726(.A1(new_n924_), .A2(new_n925_), .B1(new_n926_), .B2(new_n927_), .ZN(G1349gat));
  NAND3_X1  g727(.A1(new_n926_), .A2(new_n257_), .A3(new_n901_), .ZN(new_n929_));
  NOR2_X1   g728(.A1(new_n929_), .A2(KEYINPUT126), .ZN(new_n930_));
  NOR2_X1   g729(.A1(new_n930_), .A2(G183gat), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n929_), .A2(KEYINPUT126), .ZN(new_n932_));
  AOI21_X1  g731(.A(new_n663_), .B1(new_n295_), .B2(new_n297_), .ZN(new_n933_));
  AOI22_X1  g732(.A1(new_n931_), .A2(new_n932_), .B1(new_n923_), .B2(new_n933_), .ZN(G1350gat));
  NAND3_X1  g733(.A1(new_n915_), .A2(new_n620_), .A3(new_n917_), .ZN(new_n935_));
  INV_X1    g734(.A(KEYINPUT127), .ZN(new_n936_));
  AND3_X1   g735(.A1(new_n935_), .A2(new_n936_), .A3(G190gat), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n936_), .B1(new_n935_), .B2(G190gat), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n625_), .A2(new_n293_), .A3(new_n331_), .ZN(new_n939_));
  OAI22_X1  g738(.A1(new_n937_), .A2(new_n938_), .B1(new_n918_), .B2(new_n939_), .ZN(G1351gat));
  NOR2_X1   g739(.A1(new_n382_), .A2(new_n478_), .ZN(new_n941_));
  OAI211_X1 g740(.A(new_n450_), .B(new_n941_), .C1(new_n845_), .C2(new_n842_), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n942_), .A2(new_n725_), .ZN(new_n943_));
  XNOR2_X1  g742(.A(new_n943_), .B(new_n271_), .ZN(G1352gat));
  NOR2_X1   g743(.A1(new_n942_), .A2(new_n588_), .ZN(new_n945_));
  MUX2_X1   g744(.A(G204gat), .B(new_n269_), .S(new_n945_), .Z(G1353gat));
  NOR2_X1   g745(.A1(new_n942_), .A2(new_n663_), .ZN(new_n947_));
  NOR3_X1   g746(.A1(new_n947_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n948_));
  XOR2_X1   g747(.A(KEYINPUT63), .B(G211gat), .Z(new_n949_));
  AOI21_X1  g748(.A(new_n948_), .B1(new_n947_), .B2(new_n949_), .ZN(G1354gat));
  OAI21_X1  g749(.A(G218gat), .B1(new_n942_), .B2(new_n621_), .ZN(new_n951_));
  OR2_X1    g750(.A1(new_n626_), .A2(G218gat), .ZN(new_n952_));
  OAI21_X1  g751(.A(new_n951_), .B1(new_n942_), .B2(new_n952_), .ZN(G1355gat));
endmodule


