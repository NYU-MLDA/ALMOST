//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:33:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n663_, new_n664_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n742_, new_n743_, new_n744_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n851_, new_n852_, new_n853_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n862_, new_n863_,
    new_n864_, new_n865_, new_n866_, new_n868_, new_n870_, new_n871_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n903_, new_n904_, new_n905_, new_n907_,
    new_n908_, new_n910_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n917_, new_n918_, new_n919_, new_n920_;
  XNOR2_X1  g000(.A(G127gat), .B(G134gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G120gat), .ZN(new_n203_));
  OR2_X1    g002(.A1(new_n202_), .A2(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n202_), .A2(new_n203_), .ZN(new_n205_));
  NAND3_X1  g004(.A1(new_n204_), .A2(KEYINPUT84), .A3(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT84), .ZN(new_n207_));
  NAND3_X1  g006(.A1(new_n202_), .A2(new_n203_), .A3(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n206_), .A2(new_n208_), .ZN(new_n209_));
  XNOR2_X1  g008(.A(new_n209_), .B(KEYINPUT31), .ZN(new_n210_));
  OR2_X1    g009(.A1(new_n210_), .A2(KEYINPUT83), .ZN(new_n211_));
  XOR2_X1   g010(.A(new_n211_), .B(G99gat), .Z(new_n212_));
  INV_X1    g011(.A(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(G169gat), .ZN(new_n214_));
  OR3_X1    g013(.A1(new_n214_), .A2(KEYINPUT22), .A3(G176gat), .ZN(new_n215_));
  OAI21_X1  g014(.A(new_n214_), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NOR2_X1   g016(.A1(G183gat), .A2(G190gat), .ZN(new_n218_));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT23), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NAND3_X1  g020(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n221_), .A2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n217_), .B1(new_n218_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n223_), .ZN(new_n226_));
  INV_X1    g025(.A(G176gat), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n214_), .A2(new_n227_), .ZN(new_n228_));
  OAI21_X1  g027(.A(new_n226_), .B1(KEYINPUT24), .B2(new_n228_), .ZN(new_n229_));
  NAND2_X1  g028(.A1(G169gat), .A2(G176gat), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n228_), .A2(KEYINPUT24), .A3(new_n230_), .ZN(new_n231_));
  XNOR2_X1  g030(.A(KEYINPUT26), .B(G190gat), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT78), .ZN(new_n233_));
  INV_X1    g032(.A(G183gat), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n233_), .A2(new_n234_), .A3(KEYINPUT25), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT25), .ZN(new_n236_));
  OAI21_X1  g035(.A(KEYINPUT78), .B1(new_n236_), .B2(G183gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n232_), .A2(new_n235_), .A3(new_n237_), .ZN(new_n238_));
  OAI21_X1  g037(.A(KEYINPUT79), .B1(new_n234_), .B2(KEYINPUT25), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT79), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(new_n236_), .A3(G183gat), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n231_), .B1(new_n238_), .B2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(new_n229_), .B1(new_n243_), .B2(KEYINPUT80), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n245_));
  OAI211_X1 g044(.A(new_n245_), .B(new_n231_), .C1(new_n238_), .C2(new_n242_), .ZN(new_n246_));
  AOI21_X1  g045(.A(new_n225_), .B1(new_n244_), .B2(new_n246_), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G15gat), .B(G43gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n248_), .B(KEYINPUT82), .ZN(new_n249_));
  XOR2_X1   g048(.A(new_n247_), .B(new_n249_), .Z(new_n250_));
  XNOR2_X1  g049(.A(KEYINPUT81), .B(KEYINPUT30), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  XNOR2_X1  g052(.A(new_n247_), .B(new_n249_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n251_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(G227gat), .A2(G233gat), .ZN(new_n256_));
  INV_X1    g055(.A(G71gat), .ZN(new_n257_));
  XNOR2_X1  g056(.A(new_n256_), .B(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n253_), .A2(new_n255_), .A3(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n259_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n213_), .B1(new_n261_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n262_), .ZN(new_n264_));
  NAND3_X1  g063(.A1(new_n264_), .A2(new_n212_), .A3(new_n260_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n263_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(G155gat), .A2(G162gat), .ZN(new_n267_));
  OR2_X1    g066(.A1(G155gat), .A2(G162gat), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G141gat), .A2(G148gat), .ZN(new_n269_));
  XOR2_X1   g068(.A(new_n269_), .B(KEYINPUT3), .Z(new_n270_));
  NAND2_X1  g069(.A1(G141gat), .A2(G148gat), .ZN(new_n271_));
  XOR2_X1   g070(.A(new_n271_), .B(KEYINPUT2), .Z(new_n272_));
  OAI211_X1 g071(.A(new_n267_), .B(new_n268_), .C1(new_n270_), .C2(new_n272_), .ZN(new_n273_));
  OAI21_X1  g072(.A(KEYINPUT85), .B1(new_n267_), .B2(KEYINPUT1), .ZN(new_n274_));
  INV_X1    g073(.A(KEYINPUT85), .ZN(new_n275_));
  INV_X1    g074(.A(KEYINPUT1), .ZN(new_n276_));
  NAND4_X1  g075(.A1(new_n275_), .A2(new_n276_), .A3(G155gat), .A4(G162gat), .ZN(new_n277_));
  NAND2_X1  g076(.A1(new_n267_), .A2(KEYINPUT1), .ZN(new_n278_));
  NAND4_X1  g077(.A1(new_n274_), .A2(new_n277_), .A3(new_n278_), .A4(new_n268_), .ZN(new_n279_));
  XOR2_X1   g078(.A(G141gat), .B(G148gat), .Z(new_n280_));
  AND3_X1   g079(.A1(new_n279_), .A2(KEYINPUT86), .A3(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(KEYINPUT86), .B1(new_n279_), .B2(new_n280_), .ZN(new_n282_));
  OAI21_X1  g081(.A(new_n273_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT29), .ZN(new_n284_));
  NOR2_X1   g083(.A1(G197gat), .A2(G204gat), .ZN(new_n285_));
  INV_X1    g084(.A(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G197gat), .A2(G204gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(KEYINPUT21), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT21), .ZN(new_n289_));
  INV_X1    g088(.A(new_n287_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n289_), .B1(new_n290_), .B2(new_n285_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G211gat), .B(G218gat), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n288_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT87), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT87), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n288_), .A2(new_n291_), .A3(new_n295_), .A4(new_n292_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n292_), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n297_), .A2(KEYINPUT88), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n288_), .B1(new_n297_), .B2(KEYINPUT88), .ZN(new_n299_));
  AOI22_X1  g098(.A1(new_n294_), .A2(new_n296_), .B1(new_n298_), .B2(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G228gat), .ZN(new_n301_));
  INV_X1    g100(.A(G233gat), .ZN(new_n302_));
  NOR2_X1   g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NOR2_X1   g102(.A1(new_n300_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n284_), .A2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n303_), .ZN(new_n306_));
  XOR2_X1   g105(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n307_));
  AOI21_X1  g106(.A(new_n300_), .B1(new_n283_), .B2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n305_), .B1(new_n306_), .B2(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G78gat), .B(G106gat), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n309_), .A2(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(new_n310_), .ZN(new_n312_));
  OAI211_X1 g111(.A(new_n305_), .B(new_n312_), .C1(new_n306_), .C2(new_n308_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n311_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n313_), .ZN(new_n315_));
  NOR2_X1   g114(.A1(new_n315_), .A2(KEYINPUT90), .ZN(new_n316_));
  OR2_X1    g115(.A1(new_n283_), .A2(KEYINPUT29), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G22gat), .B(G50gat), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n318_), .B(KEYINPUT28), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n317_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n320_), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n314_), .B1(new_n316_), .B2(new_n321_), .ZN(new_n322_));
  NAND4_X1  g121(.A1(new_n311_), .A2(new_n320_), .A3(KEYINPUT90), .A4(new_n313_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(G226gat), .A2(G233gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(new_n325_), .B(KEYINPUT19), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n243_), .A2(KEYINPUT80), .ZN(new_n327_));
  INV_X1    g126(.A(new_n229_), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n327_), .A2(new_n246_), .A3(new_n328_), .ZN(new_n329_));
  NAND3_X1  g128(.A1(new_n329_), .A2(new_n300_), .A3(new_n224_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n330_), .A2(KEYINPUT91), .A3(KEYINPUT20), .ZN(new_n331_));
  XOR2_X1   g130(.A(KEYINPUT92), .B(KEYINPUT24), .Z(new_n332_));
  OAI21_X1  g131(.A(new_n226_), .B1(new_n332_), .B2(new_n228_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n332_), .A2(new_n228_), .A3(new_n230_), .ZN(new_n335_));
  XNOR2_X1  g134(.A(KEYINPUT25), .B(G183gat), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(new_n232_), .ZN(new_n337_));
  NAND4_X1  g136(.A1(new_n334_), .A2(KEYINPUT93), .A3(new_n335_), .A4(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT93), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n335_), .A2(new_n337_), .ZN(new_n340_));
  OAI21_X1  g139(.A(new_n339_), .B1(new_n340_), .B2(new_n333_), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n225_), .A2(KEYINPUT94), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT94), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n224_), .A2(new_n343_), .ZN(new_n344_));
  OAI211_X1 g143(.A(new_n338_), .B(new_n341_), .C1(new_n342_), .C2(new_n344_), .ZN(new_n345_));
  INV_X1    g144(.A(new_n300_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n345_), .A2(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n331_), .A2(new_n347_), .ZN(new_n348_));
  AOI21_X1  g147(.A(KEYINPUT91), .B1(new_n330_), .B2(KEYINPUT20), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n326_), .B1(new_n348_), .B2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G8gat), .B(G36gat), .Z(new_n351_));
  XNOR2_X1  g150(.A(KEYINPUT95), .B(KEYINPUT18), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n351_), .B(new_n352_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(G64gat), .B(G92gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n353_), .B(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n326_), .ZN(new_n357_));
  OAI211_X1 g156(.A(KEYINPUT20), .B(new_n357_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n358_));
  NOR2_X1   g157(.A1(new_n247_), .A2(new_n300_), .ZN(new_n359_));
  OR2_X1    g158(.A1(new_n358_), .A2(new_n359_), .ZN(new_n360_));
  AND3_X1   g159(.A1(new_n350_), .A2(new_n356_), .A3(new_n360_), .ZN(new_n361_));
  AOI21_X1  g160(.A(new_n356_), .B1(new_n350_), .B2(new_n360_), .ZN(new_n362_));
  OAI21_X1  g161(.A(KEYINPUT96), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  INV_X1    g162(.A(KEYINPUT20), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n364_), .B1(new_n247_), .B2(new_n300_), .ZN(new_n365_));
  AOI22_X1  g164(.A1(new_n365_), .A2(KEYINPUT91), .B1(new_n346_), .B2(new_n345_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n349_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n357_), .B1(new_n366_), .B2(new_n367_), .ZN(new_n368_));
  NOR2_X1   g167(.A1(new_n358_), .A2(new_n359_), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n355_), .B1(new_n368_), .B2(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT96), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n350_), .A2(new_n360_), .A3(new_n356_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n370_), .A2(new_n371_), .A3(new_n372_), .ZN(new_n373_));
  XOR2_X1   g172(.A(G1gat), .B(G29gat), .Z(new_n374_));
  XNOR2_X1  g173(.A(G57gat), .B(G85gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(new_n374_), .B(new_n375_), .ZN(new_n376_));
  XNOR2_X1  g175(.A(KEYINPUT97), .B(KEYINPUT0), .ZN(new_n377_));
  XNOR2_X1  g176(.A(new_n376_), .B(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT4), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n283_), .A2(new_n209_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n204_), .A2(new_n205_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n273_), .B(new_n382_), .C1(new_n281_), .C2(new_n282_), .ZN(new_n383_));
  AOI21_X1  g182(.A(new_n380_), .B1(new_n381_), .B2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT4), .B1(new_n283_), .B2(new_n209_), .ZN(new_n386_));
  NOR3_X1   g185(.A1(new_n384_), .A2(new_n385_), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n381_), .A2(new_n383_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n388_), .A2(new_n385_), .ZN(new_n389_));
  INV_X1    g188(.A(new_n389_), .ZN(new_n390_));
  OAI211_X1 g189(.A(KEYINPUT33), .B(new_n379_), .C1(new_n387_), .C2(new_n390_), .ZN(new_n391_));
  AOI21_X1  g190(.A(new_n386_), .B1(new_n388_), .B2(KEYINPUT4), .ZN(new_n392_));
  INV_X1    g191(.A(new_n385_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(new_n378_), .B1(new_n394_), .B2(new_n389_), .ZN(new_n395_));
  INV_X1    g194(.A(KEYINPUT33), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n385_), .B1(new_n384_), .B2(new_n386_), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n381_), .A2(new_n383_), .A3(new_n393_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n398_), .A2(new_n378_), .ZN(new_n399_));
  AOI21_X1  g198(.A(new_n396_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n400_));
  OAI21_X1  g199(.A(new_n391_), .B1(new_n395_), .B2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n363_), .A2(new_n373_), .A3(new_n402_), .ZN(new_n403_));
  NAND3_X1  g202(.A1(new_n366_), .A2(new_n357_), .A3(new_n367_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n224_), .B1(new_n340_), .B2(new_n333_), .ZN(new_n405_));
  OAI21_X1  g204(.A(KEYINPUT20), .B1(new_n346_), .B2(new_n405_), .ZN(new_n406_));
  OAI21_X1  g205(.A(new_n326_), .B1(new_n359_), .B2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT99), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  OAI211_X1 g208(.A(KEYINPUT99), .B(new_n326_), .C1(new_n359_), .C2(new_n406_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n404_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n356_), .A2(KEYINPUT32), .ZN(new_n412_));
  INV_X1    g211(.A(new_n412_), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n379_), .B1(new_n387_), .B2(new_n390_), .ZN(new_n414_));
  NAND3_X1  g213(.A1(new_n394_), .A2(new_n378_), .A3(new_n389_), .ZN(new_n415_));
  AOI22_X1  g214(.A1(new_n411_), .A2(new_n413_), .B1(new_n414_), .B2(new_n415_), .ZN(new_n416_));
  NAND3_X1  g215(.A1(new_n350_), .A2(new_n360_), .A3(new_n412_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT98), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n417_), .A2(new_n418_), .ZN(new_n419_));
  NOR2_X1   g218(.A1(new_n417_), .A2(new_n418_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n416_), .B1(new_n419_), .B2(new_n420_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n324_), .B1(new_n403_), .B2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n370_), .A2(new_n372_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(KEYINPUT100), .B(KEYINPUT27), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n423_), .A2(new_n424_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n415_), .A2(new_n414_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n322_), .B2(new_n323_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n411_), .A2(new_n355_), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n428_), .A2(KEYINPUT27), .A3(new_n372_), .ZN(new_n429_));
  AND3_X1   g228(.A1(new_n425_), .A2(new_n427_), .A3(new_n429_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n266_), .B1(new_n422_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n425_), .A2(new_n429_), .ZN(new_n432_));
  NOR2_X1   g231(.A1(new_n432_), .A2(new_n324_), .ZN(new_n433_));
  INV_X1    g232(.A(new_n426_), .ZN(new_n434_));
  INV_X1    g233(.A(new_n266_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n433_), .A2(new_n434_), .A3(new_n435_), .ZN(new_n436_));
  AND2_X1   g235(.A1(new_n431_), .A2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(KEYINPUT77), .ZN(new_n438_));
  NAND2_X1  g237(.A1(G229gat), .A2(G233gat), .ZN(new_n439_));
  INV_X1    g238(.A(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G15gat), .B(G22gat), .ZN(new_n441_));
  INV_X1    g240(.A(G1gat), .ZN(new_n442_));
  INV_X1    g241(.A(G8gat), .ZN(new_n443_));
  OAI21_X1  g242(.A(KEYINPUT14), .B1(new_n442_), .B2(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(new_n441_), .B1(new_n444_), .B2(KEYINPUT74), .ZN(new_n445_));
  AND2_X1   g244(.A1(new_n444_), .A2(KEYINPUT74), .ZN(new_n446_));
  XNOR2_X1  g245(.A(G1gat), .B(G8gat), .ZN(new_n447_));
  OR3_X1    g246(.A1(new_n445_), .A2(new_n446_), .A3(new_n447_), .ZN(new_n448_));
  OAI21_X1  g247(.A(new_n447_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n449_));
  AND2_X1   g248(.A1(new_n448_), .A2(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G29gat), .B(G36gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(G43gat), .B(G50gat), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n451_), .B(new_n452_), .ZN(new_n453_));
  AND2_X1   g252(.A1(new_n450_), .A2(new_n453_), .ZN(new_n454_));
  NOR2_X1   g253(.A1(new_n450_), .A2(new_n453_), .ZN(new_n455_));
  OAI21_X1  g254(.A(new_n440_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n453_), .B(KEYINPUT15), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n448_), .A2(new_n449_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n450_), .A2(new_n453_), .ZN(new_n460_));
  NAND3_X1  g259(.A1(new_n459_), .A2(new_n460_), .A3(new_n439_), .ZN(new_n461_));
  XNOR2_X1  g260(.A(G113gat), .B(G141gat), .ZN(new_n462_));
  XNOR2_X1  g261(.A(new_n462_), .B(KEYINPUT76), .ZN(new_n463_));
  XNOR2_X1  g262(.A(G169gat), .B(G197gat), .ZN(new_n464_));
  XNOR2_X1  g263(.A(new_n463_), .B(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n456_), .A2(new_n461_), .A3(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(new_n467_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n466_), .B1(new_n456_), .B2(new_n461_), .ZN(new_n469_));
  OAI21_X1  g268(.A(new_n438_), .B1(new_n468_), .B2(new_n469_), .ZN(new_n470_));
  INV_X1    g269(.A(new_n469_), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n471_), .A2(KEYINPUT77), .A3(new_n467_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n470_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT13), .ZN(new_n475_));
  XNOR2_X1  g274(.A(G120gat), .B(G148gat), .ZN(new_n476_));
  XNOR2_X1  g275(.A(new_n476_), .B(KEYINPUT5), .ZN(new_n477_));
  XNOR2_X1  g276(.A(G176gat), .B(G204gat), .ZN(new_n478_));
  XOR2_X1   g277(.A(new_n477_), .B(new_n478_), .Z(new_n479_));
  NAND2_X1  g278(.A1(G230gat), .A2(G233gat), .ZN(new_n480_));
  INV_X1    g279(.A(G64gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(G57gat), .ZN(new_n482_));
  INV_X1    g281(.A(G57gat), .ZN(new_n483_));
  NAND2_X1  g282(.A1(new_n483_), .A2(G64gat), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n482_), .A2(new_n484_), .A3(KEYINPUT11), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n257_), .A2(KEYINPUT68), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT68), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(G71gat), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n487_), .A2(new_n489_), .ZN(new_n490_));
  NOR2_X1   g289(.A1(new_n490_), .A2(G78gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(KEYINPUT68), .B(G71gat), .ZN(new_n492_));
  INV_X1    g291(.A(G78gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  OAI21_X1  g293(.A(new_n486_), .B1(new_n491_), .B2(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n490_), .A2(G78gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n492_), .A2(new_n493_), .ZN(new_n497_));
  AOI21_X1  g296(.A(KEYINPUT11), .B1(new_n482_), .B2(new_n484_), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n496_), .B(new_n497_), .C1(new_n485_), .C2(new_n498_), .ZN(new_n499_));
  AND2_X1   g298(.A1(new_n495_), .A2(new_n499_), .ZN(new_n500_));
  OR3_X1    g299(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n502_));
  NAND2_X1  g301(.A1(G99gat), .A2(G106gat), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n503_), .A2(KEYINPUT6), .ZN(new_n504_));
  NOR2_X1   g303(.A1(new_n503_), .A2(KEYINPUT6), .ZN(new_n505_));
  OAI211_X1 g304(.A(new_n501_), .B(new_n502_), .C1(new_n504_), .C2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT8), .ZN(new_n507_));
  XNOR2_X1  g306(.A(G85gat), .B(G92gat), .ZN(new_n508_));
  OAI21_X1  g307(.A(new_n507_), .B1(new_n508_), .B2(KEYINPUT67), .ZN(new_n509_));
  INV_X1    g308(.A(new_n508_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n506_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n511_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n509_), .B1(new_n506_), .B2(new_n510_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n504_), .A2(new_n505_), .ZN(new_n515_));
  INV_X1    g314(.A(G106gat), .ZN(new_n516_));
  XOR2_X1   g315(.A(KEYINPUT10), .B(G99gat), .Z(new_n517_));
  AOI21_X1  g316(.A(new_n515_), .B1(new_n516_), .B2(new_n517_), .ZN(new_n518_));
  NAND3_X1  g317(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n519_));
  XNOR2_X1  g318(.A(new_n519_), .B(KEYINPUT65), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT9), .ZN(new_n521_));
  AOI22_X1  g320(.A1(new_n521_), .A2(KEYINPUT64), .B1(G85gat), .B2(G92gat), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT64), .ZN(new_n523_));
  NAND2_X1  g322(.A1(new_n523_), .A2(KEYINPUT9), .ZN(new_n524_));
  INV_X1    g323(.A(G85gat), .ZN(new_n525_));
  INV_X1    g324(.A(G92gat), .ZN(new_n526_));
  AOI22_X1  g325(.A1(new_n522_), .A2(new_n524_), .B1(new_n525_), .B2(new_n526_), .ZN(new_n527_));
  AND3_X1   g326(.A1(new_n520_), .A2(new_n527_), .A3(KEYINPUT66), .ZN(new_n528_));
  AOI21_X1  g327(.A(KEYINPUT66), .B1(new_n520_), .B2(new_n527_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n518_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  AOI21_X1  g329(.A(new_n500_), .B1(new_n514_), .B2(new_n530_), .ZN(new_n531_));
  AOI21_X1  g330(.A(new_n480_), .B1(new_n531_), .B2(KEYINPUT69), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n495_), .A2(new_n499_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(new_n517_), .A2(new_n516_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n534_), .B1(new_n504_), .B2(new_n505_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n520_), .A2(new_n527_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT66), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n520_), .A2(new_n527_), .A3(KEYINPUT66), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n535_), .B1(new_n538_), .B2(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n506_), .A2(new_n510_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n509_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n543_), .A2(new_n511_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n533_), .B1(new_n540_), .B2(new_n544_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT69), .ZN(new_n546_));
  NAND3_X1  g345(.A1(new_n514_), .A2(new_n530_), .A3(new_n500_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n545_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n532_), .A2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  INV_X1    g349(.A(new_n480_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n545_), .A2(KEYINPUT12), .A3(new_n547_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n514_), .A2(new_n530_), .ZN(new_n553_));
  INV_X1    g352(.A(KEYINPUT12), .ZN(new_n554_));
  NAND3_X1  g353(.A1(new_n553_), .A2(new_n554_), .A3(new_n533_), .ZN(new_n555_));
  AOI21_X1  g354(.A(new_n551_), .B1(new_n552_), .B2(new_n555_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n479_), .B1(new_n550_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n552_), .A2(new_n555_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n558_), .A2(new_n480_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n479_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n559_), .A2(new_n549_), .A3(new_n560_), .ZN(new_n561_));
  AND3_X1   g360(.A1(new_n557_), .A2(new_n561_), .A3(KEYINPUT70), .ZN(new_n562_));
  AOI21_X1  g361(.A(KEYINPUT70), .B1(new_n557_), .B2(new_n561_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n475_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n557_), .A2(new_n561_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT70), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n565_), .A2(new_n566_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n557_), .A2(new_n561_), .A3(KEYINPUT70), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(KEYINPUT13), .A3(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n564_), .A2(new_n569_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n553_), .A2(new_n457_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(G232gat), .A2(G233gat), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT34), .ZN(new_n573_));
  INV_X1    g372(.A(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT35), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n514_), .A2(new_n530_), .A3(new_n453_), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n571_), .A2(new_n576_), .A3(new_n577_), .ZN(new_n578_));
  NOR2_X1   g377(.A1(new_n574_), .A2(new_n575_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n579_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n571_), .A2(new_n581_), .A3(new_n576_), .A4(new_n577_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(new_n580_), .A2(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(G190gat), .B(G218gat), .Z(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(KEYINPUT71), .ZN(new_n585_));
  XNOR2_X1  g384(.A(G134gat), .B(G162gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n587_), .A2(KEYINPUT36), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n587_), .A2(KEYINPUT36), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n588_), .A2(new_n589_), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n583_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(KEYINPUT73), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT37), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n583_), .A2(new_n590_), .ZN(new_n594_));
  INV_X1    g393(.A(KEYINPUT73), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n580_), .A2(new_n589_), .A3(new_n582_), .ZN(new_n597_));
  NAND4_X1  g396(.A1(new_n592_), .A2(new_n593_), .A3(new_n596_), .A4(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT72), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  NAND4_X1  g399(.A1(new_n580_), .A2(KEYINPUT72), .A3(new_n589_), .A4(new_n582_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n600_), .A2(new_n594_), .A3(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n602_), .A2(KEYINPUT37), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n598_), .A2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n458_), .B(new_n605_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n606_), .A2(new_n533_), .ZN(new_n607_));
  NOR2_X1   g406(.A1(new_n450_), .A2(new_n605_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n458_), .B1(G231gat), .B2(G233gat), .ZN(new_n609_));
  OAI21_X1  g408(.A(new_n500_), .B1(new_n608_), .B2(new_n609_), .ZN(new_n610_));
  XOR2_X1   g409(.A(G127gat), .B(G155gat), .Z(new_n611_));
  XNOR2_X1  g410(.A(new_n611_), .B(KEYINPUT16), .ZN(new_n612_));
  XNOR2_X1  g411(.A(G183gat), .B(G211gat), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(KEYINPUT17), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n614_), .B(new_n615_), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n607_), .A2(new_n610_), .A3(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n614_), .A2(new_n615_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n619_), .B1(new_n607_), .B2(new_n610_), .ZN(new_n620_));
  OAI21_X1  g419(.A(KEYINPUT75), .B1(new_n618_), .B2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n620_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT75), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n622_), .A2(new_n623_), .A3(new_n617_), .ZN(new_n624_));
  NAND2_X1  g423(.A1(new_n621_), .A2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n604_), .A2(new_n626_), .ZN(new_n627_));
  NOR4_X1   g426(.A1(new_n437_), .A2(new_n474_), .A3(new_n570_), .A4(new_n627_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n628_), .A2(new_n442_), .A3(new_n426_), .ZN(new_n629_));
  INV_X1    g428(.A(KEYINPUT38), .ZN(new_n630_));
  OR2_X1    g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n596_), .A2(new_n597_), .ZN(new_n632_));
  NOR2_X1   g431(.A1(new_n594_), .A2(new_n595_), .ZN(new_n633_));
  OAI21_X1  g432(.A(KEYINPUT102), .B1(new_n632_), .B2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT102), .ZN(new_n635_));
  NAND4_X1  g434(.A1(new_n592_), .A2(new_n635_), .A3(new_n596_), .A4(new_n597_), .ZN(new_n636_));
  AND2_X1   g435(.A1(new_n634_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NOR2_X1   g437(.A1(new_n437_), .A2(new_n638_), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n564_), .A2(new_n569_), .A3(new_n473_), .ZN(new_n640_));
  OR2_X1    g439(.A1(new_n640_), .A2(KEYINPUT101), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(KEYINPUT101), .ZN(new_n642_));
  AND3_X1   g441(.A1(new_n641_), .A2(new_n626_), .A3(new_n642_), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n639_), .A2(new_n426_), .A3(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n644_), .A2(G1gat), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n629_), .A2(new_n630_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n631_), .A2(new_n645_), .A3(new_n646_), .ZN(G1324gat));
  NAND3_X1  g446(.A1(new_n639_), .A2(new_n432_), .A3(new_n643_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n648_), .A2(G8gat), .ZN(new_n649_));
  XNOR2_X1  g448(.A(new_n649_), .B(KEYINPUT39), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n628_), .A2(new_n443_), .A3(new_n432_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n650_), .A2(new_n651_), .A3(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n652_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(G1325gat));
  INV_X1    g455(.A(G15gat), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n628_), .A2(new_n657_), .A3(new_n435_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n639_), .A2(new_n435_), .A3(new_n643_), .ZN(new_n659_));
  AND3_X1   g458(.A1(new_n659_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n660_));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(new_n659_), .B2(G15gat), .ZN(new_n661_));
  OAI21_X1  g460(.A(new_n658_), .B1(new_n660_), .B2(new_n661_), .ZN(G1326gat));
  INV_X1    g461(.A(G22gat), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n628_), .A2(new_n663_), .A3(new_n324_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n639_), .A2(new_n324_), .A3(new_n643_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT42), .ZN(new_n666_));
  AND3_X1   g465(.A1(new_n665_), .A2(new_n666_), .A3(G22gat), .ZN(new_n667_));
  AOI21_X1  g466(.A(new_n666_), .B1(new_n665_), .B2(G22gat), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n664_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  XOR2_X1   g468(.A(new_n669_), .B(KEYINPUT104), .Z(G1327gat));
  NAND2_X1  g469(.A1(new_n431_), .A2(new_n436_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n570_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n637_), .A2(new_n626_), .ZN(new_n673_));
  AND4_X1   g472(.A1(new_n671_), .A2(new_n473_), .A3(new_n672_), .A4(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n426_), .ZN(new_n675_));
  INV_X1    g474(.A(new_n604_), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT43), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n676_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n671_), .A2(new_n679_), .ZN(new_n680_));
  OR2_X1    g479(.A1(new_n604_), .A2(KEYINPUT105), .ZN(new_n681_));
  NAND2_X1  g480(.A1(new_n604_), .A2(KEYINPUT105), .ZN(new_n682_));
  AOI22_X1  g481(.A1(new_n431_), .A2(new_n436_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  OAI21_X1  g482(.A(new_n680_), .B1(new_n683_), .B2(new_n677_), .ZN(new_n684_));
  NAND3_X1  g483(.A1(new_n641_), .A2(new_n625_), .A3(new_n642_), .ZN(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n684_), .A2(KEYINPUT44), .A3(new_n686_), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n681_), .A2(new_n682_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n677_), .B1(new_n671_), .B2(new_n688_), .ZN(new_n689_));
  AOI21_X1  g488(.A(new_n678_), .B1(new_n431_), .B2(new_n436_), .ZN(new_n690_));
  OAI21_X1  g489(.A(new_n686_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  AOI21_X1  g490(.A(KEYINPUT44), .B1(new_n691_), .B2(KEYINPUT106), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT106), .ZN(new_n693_));
  NAND3_X1  g492(.A1(new_n684_), .A2(new_n693_), .A3(new_n686_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n687_), .B1(new_n692_), .B2(new_n694_), .ZN(new_n695_));
  AND2_X1   g494(.A1(new_n426_), .A2(G29gat), .ZN(new_n696_));
  AOI21_X1  g495(.A(new_n675_), .B1(new_n695_), .B2(new_n696_), .ZN(G1328gat));
  INV_X1    g496(.A(KEYINPUT46), .ZN(new_n698_));
  INV_X1    g497(.A(G36gat), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n699_), .B1(new_n695_), .B2(new_n432_), .ZN(new_n700_));
  NAND3_X1  g499(.A1(new_n674_), .A2(new_n699_), .A3(new_n432_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n702_));
  OR2_X1    g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n701_), .A2(new_n702_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n698_), .B1(new_n700_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n705_), .ZN(new_n707_));
  INV_X1    g506(.A(new_n432_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n671_), .A2(new_n688_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n709_), .A2(KEYINPUT43), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n685_), .B1(new_n710_), .B2(new_n680_), .ZN(new_n711_));
  AOI221_X4 g510(.A(new_n708_), .B1(new_n711_), .B2(KEYINPUT44), .C1(new_n692_), .C2(new_n694_), .ZN(new_n712_));
  OAI211_X1 g511(.A(new_n707_), .B(KEYINPUT46), .C1(new_n712_), .C2(new_n699_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n706_), .A2(new_n713_), .ZN(G1329gat));
  AND2_X1   g513(.A1(new_n674_), .A2(new_n435_), .ZN(new_n715_));
  NOR2_X1   g514(.A1(new_n715_), .A2(G43gat), .ZN(new_n716_));
  AND2_X1   g515(.A1(new_n435_), .A2(G43gat), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n716_), .B1(new_n695_), .B2(new_n717_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n719_));
  NOR2_X1   g518(.A1(new_n718_), .A2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n719_), .ZN(new_n721_));
  AOI211_X1 g520(.A(new_n716_), .B(new_n721_), .C1(new_n695_), .C2(new_n717_), .ZN(new_n722_));
  NOR2_X1   g521(.A1(new_n720_), .A2(new_n722_), .ZN(G1330gat));
  INV_X1    g522(.A(G50gat), .ZN(new_n724_));
  NAND3_X1  g523(.A1(new_n674_), .A2(new_n724_), .A3(new_n324_), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n695_), .A2(KEYINPUT109), .A3(new_n324_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(G50gat), .ZN(new_n727_));
  AOI21_X1  g526(.A(KEYINPUT109), .B1(new_n695_), .B2(new_n324_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n725_), .B1(new_n727_), .B2(new_n728_), .ZN(G1331gat));
  NOR4_X1   g528(.A1(new_n437_), .A2(new_n473_), .A3(new_n672_), .A4(new_n627_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(new_n483_), .A3(new_n426_), .ZN(new_n731_));
  AND4_X1   g530(.A1(new_n470_), .A2(new_n621_), .A3(new_n624_), .A4(new_n472_), .ZN(new_n732_));
  AND3_X1   g531(.A1(new_n639_), .A2(new_n570_), .A3(new_n732_), .ZN(new_n733_));
  AND2_X1   g532(.A1(new_n733_), .A2(new_n426_), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n731_), .B1(new_n734_), .B2(new_n483_), .ZN(G1332gat));
  AOI21_X1  g534(.A(new_n481_), .B1(new_n733_), .B2(new_n432_), .ZN(new_n736_));
  XOR2_X1   g535(.A(new_n736_), .B(KEYINPUT48), .Z(new_n737_));
  NAND2_X1  g536(.A1(new_n432_), .A2(new_n481_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT110), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n730_), .A2(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n737_), .A2(new_n740_), .ZN(G1333gat));
  AOI21_X1  g540(.A(new_n257_), .B1(new_n733_), .B2(new_n435_), .ZN(new_n742_));
  XOR2_X1   g541(.A(new_n742_), .B(KEYINPUT49), .Z(new_n743_));
  NAND3_X1  g542(.A1(new_n730_), .A2(new_n257_), .A3(new_n435_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(G1334gat));
  AOI21_X1  g544(.A(new_n493_), .B1(new_n733_), .B2(new_n324_), .ZN(new_n746_));
  XOR2_X1   g545(.A(new_n746_), .B(KEYINPUT50), .Z(new_n747_));
  NAND3_X1  g546(.A1(new_n730_), .A2(new_n493_), .A3(new_n324_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1335gat));
  NOR3_X1   g548(.A1(new_n672_), .A2(new_n473_), .A3(new_n626_), .ZN(new_n750_));
  AND2_X1   g549(.A1(new_n684_), .A2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n434_), .ZN(new_n753_));
  AND4_X1   g552(.A1(new_n671_), .A2(new_n474_), .A3(new_n570_), .A4(new_n673_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n754_), .A2(new_n525_), .A3(new_n426_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(G1336gat));
  OAI21_X1  g555(.A(G92gat), .B1(new_n752_), .B2(new_n708_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n754_), .A2(new_n526_), .A3(new_n432_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n757_), .A2(new_n758_), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n752_), .B2(new_n266_), .ZN(new_n760_));
  NAND3_X1  g559(.A1(new_n754_), .A2(new_n435_), .A3(new_n517_), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  XNOR2_X1  g561(.A(new_n762_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g562(.A1(new_n754_), .A2(new_n516_), .A3(new_n324_), .ZN(new_n764_));
  NAND3_X1  g563(.A1(new_n684_), .A2(new_n324_), .A3(new_n750_), .ZN(new_n765_));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766_));
  AND3_X1   g565(.A1(new_n765_), .A2(new_n766_), .A3(G106gat), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n766_), .B1(new_n765_), .B2(G106gat), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  XNOR2_X1  g568(.A(new_n769_), .B(KEYINPUT53), .ZN(G1339gat));
  XNOR2_X1  g569(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n771_));
  INV_X1    g570(.A(new_n771_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n564_), .A2(new_n569_), .A3(new_n732_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n773_), .A2(KEYINPUT111), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT111), .ZN(new_n775_));
  NAND4_X1  g574(.A1(new_n564_), .A2(new_n569_), .A3(new_n732_), .A4(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n774_), .A2(new_n776_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n772_), .B1(new_n777_), .B2(new_n604_), .ZN(new_n778_));
  AOI211_X1 g577(.A(new_n676_), .B(new_n771_), .C1(new_n774_), .C2(new_n776_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n552_), .A2(new_n551_), .A3(new_n555_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n559_), .A2(KEYINPUT55), .A3(new_n781_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n783_));
  AOI21_X1  g582(.A(new_n560_), .B1(new_n556_), .B2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(KEYINPUT56), .A3(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(new_n785_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT56), .B1(new_n782_), .B2(new_n784_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789_));
  NOR3_X1   g588(.A1(new_n550_), .A2(new_n556_), .A3(new_n479_), .ZN(new_n790_));
  OAI21_X1  g589(.A(new_n439_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n459_), .A2(new_n460_), .A3(new_n440_), .ZN(new_n792_));
  NAND3_X1  g591(.A1(new_n791_), .A2(new_n465_), .A3(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n467_), .A2(new_n793_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n789_), .B1(new_n790_), .B2(new_n794_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n467_), .A2(new_n793_), .ZN(new_n796_));
  NAND3_X1  g595(.A1(new_n796_), .A2(KEYINPUT115), .A3(new_n561_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n795_), .A2(new_n797_), .ZN(new_n798_));
  OAI21_X1  g597(.A(KEYINPUT116), .B1(new_n788_), .B2(new_n798_), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n799_), .A2(KEYINPUT58), .ZN(new_n800_));
  INV_X1    g599(.A(KEYINPUT58), .ZN(new_n801_));
  OAI211_X1 g600(.A(KEYINPUT116), .B(new_n801_), .C1(new_n788_), .C2(new_n798_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n800_), .A2(new_n676_), .A3(new_n802_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n796_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT113), .ZN(new_n805_));
  AND3_X1   g604(.A1(new_n552_), .A2(new_n551_), .A3(new_n555_), .ZN(new_n806_));
  NOR3_X1   g605(.A1(new_n806_), .A2(new_n556_), .A3(new_n783_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n558_), .A2(new_n783_), .A3(new_n480_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n479_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n805_), .B1(new_n807_), .B2(new_n809_), .ZN(new_n810_));
  INV_X1    g609(.A(KEYINPUT114), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT56), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n782_), .A2(KEYINPUT113), .A3(new_n784_), .ZN(new_n813_));
  NAND4_X1  g612(.A1(new_n810_), .A2(new_n811_), .A3(new_n812_), .A4(new_n813_), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n790_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n814_), .A2(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n785_), .A2(KEYINPUT114), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n782_), .A2(new_n784_), .ZN(new_n818_));
  AOI21_X1  g617(.A(KEYINPUT56), .B1(new_n818_), .B2(new_n805_), .ZN(new_n819_));
  AOI21_X1  g618(.A(new_n817_), .B1(new_n819_), .B2(new_n813_), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n804_), .B1(new_n816_), .B2(new_n820_), .ZN(new_n821_));
  AND3_X1   g620(.A1(new_n634_), .A2(KEYINPUT57), .A3(new_n636_), .ZN(new_n822_));
  NAND2_X1  g621(.A1(new_n821_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n803_), .A2(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT57), .B1(new_n821_), .B2(new_n637_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n625_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n780_), .A2(new_n826_), .ZN(new_n827_));
  NOR4_X1   g626(.A1(new_n432_), .A2(new_n266_), .A3(new_n324_), .A4(new_n434_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT59), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n829_), .A2(KEYINPUT117), .ZN(new_n830_));
  INV_X1    g629(.A(new_n830_), .ZN(new_n831_));
  NAND3_X1  g630(.A1(new_n827_), .A2(new_n828_), .A3(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n832_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n834_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT118), .B1(new_n833_), .B2(new_n835_), .ZN(new_n836_));
  INV_X1    g635(.A(KEYINPUT118), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n827_), .A2(new_n828_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  OAI211_X1 g638(.A(new_n832_), .B(new_n837_), .C1(new_n839_), .C2(new_n834_), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n836_), .A2(new_n840_), .A3(new_n473_), .ZN(new_n841_));
  NAND2_X1  g640(.A1(new_n841_), .A2(G113gat), .ZN(new_n842_));
  OR3_X1    g641(.A1(new_n838_), .A2(G113gat), .A3(new_n474_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(G1340gat));
  INV_X1    g643(.A(G120gat), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n845_), .B1(new_n672_), .B2(KEYINPUT60), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n839_), .B(new_n846_), .C1(KEYINPUT60), .C2(new_n845_), .ZN(new_n847_));
  OAI211_X1 g646(.A(new_n570_), .B(new_n832_), .C1(new_n839_), .C2(new_n834_), .ZN(new_n848_));
  INV_X1    g647(.A(new_n848_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n847_), .B1(new_n849_), .B2(new_n845_), .ZN(G1341gat));
  NAND3_X1  g649(.A1(new_n836_), .A2(new_n840_), .A3(new_n626_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(G127gat), .ZN(new_n852_));
  OR3_X1    g651(.A1(new_n838_), .A2(G127gat), .A3(new_n625_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n852_), .A2(new_n853_), .ZN(G1342gat));
  INV_X1    g653(.A(G134gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n838_), .B2(new_n637_), .ZN(new_n856_));
  XNOR2_X1  g655(.A(new_n856_), .B(KEYINPUT119), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n676_), .A2(G134gat), .ZN(new_n858_));
  XNOR2_X1  g657(.A(new_n858_), .B(KEYINPUT120), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n836_), .A2(new_n840_), .A3(new_n859_), .ZN(new_n860_));
  AND2_X1   g659(.A1(new_n857_), .A2(new_n860_), .ZN(G1343gat));
  AND4_X1   g660(.A1(new_n324_), .A2(new_n708_), .A3(new_n426_), .A4(new_n266_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n827_), .A2(new_n862_), .ZN(new_n863_));
  AND2_X1   g662(.A1(new_n863_), .A2(KEYINPUT121), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n863_), .A2(KEYINPUT121), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n473_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n866_), .B(G141gat), .ZN(G1344gat));
  OAI21_X1  g666(.A(new_n570_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n868_));
  XNOR2_X1  g667(.A(new_n868_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g668(.A(new_n626_), .B1(new_n864_), .B2(new_n865_), .ZN(new_n870_));
  XNOR2_X1  g669(.A(KEYINPUT61), .B(G155gat), .ZN(new_n871_));
  XNOR2_X1  g670(.A(new_n870_), .B(new_n871_), .ZN(G1346gat));
  OR2_X1    g671(.A1(new_n864_), .A2(new_n865_), .ZN(new_n873_));
  NAND2_X1  g672(.A1(new_n873_), .A2(new_n638_), .ZN(new_n874_));
  INV_X1    g673(.A(G162gat), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n875_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n874_), .A2(new_n875_), .B1(new_n873_), .B2(new_n876_), .ZN(G1347gat));
  NOR3_X1   g676(.A1(new_n266_), .A2(new_n324_), .A3(new_n426_), .ZN(new_n878_));
  NAND4_X1  g677(.A1(new_n827_), .A2(new_n432_), .A3(new_n473_), .A4(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(KEYINPUT62), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n879_), .A2(new_n880_), .A3(G169gat), .ZN(new_n881_));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n882_));
  AND2_X1   g681(.A1(new_n881_), .A2(new_n882_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n881_), .A2(new_n882_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n879_), .A2(G169gat), .ZN(new_n885_));
  AOI21_X1  g684(.A(KEYINPUT123), .B1(new_n885_), .B2(KEYINPUT62), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887_));
  AOI211_X1 g686(.A(new_n887_), .B(new_n880_), .C1(new_n879_), .C2(G169gat), .ZN(new_n888_));
  OAI22_X1  g687(.A1(new_n883_), .A2(new_n884_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n889_));
  AND3_X1   g688(.A1(new_n827_), .A2(new_n432_), .A3(new_n878_), .ZN(new_n890_));
  XNOR2_X1  g689(.A(KEYINPUT22), .B(G169gat), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n473_), .A2(new_n891_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(new_n892_), .B(KEYINPUT124), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n890_), .A2(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n889_), .A2(new_n894_), .ZN(G1348gat));
  AOI21_X1  g694(.A(new_n672_), .B1(KEYINPUT125), .B2(new_n227_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n890_), .A2(new_n896_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n227_), .A2(KEYINPUT125), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n897_), .B(new_n898_), .ZN(G1349gat));
  NAND2_X1  g698(.A1(new_n890_), .A2(new_n626_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n900_), .A2(new_n336_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n901_), .B1(new_n234_), .B2(new_n900_), .ZN(G1350gat));
  NAND3_X1  g701(.A1(new_n890_), .A2(new_n232_), .A3(new_n638_), .ZN(new_n903_));
  AND2_X1   g702(.A1(new_n890_), .A2(new_n676_), .ZN(new_n904_));
  INV_X1    g703(.A(G190gat), .ZN(new_n905_));
  OAI21_X1  g704(.A(new_n903_), .B1(new_n904_), .B2(new_n905_), .ZN(G1351gat));
  NAND4_X1  g705(.A1(new_n827_), .A2(new_n427_), .A3(new_n432_), .A4(new_n266_), .ZN(new_n907_));
  NOR2_X1   g706(.A1(new_n907_), .A2(new_n474_), .ZN(new_n908_));
  XOR2_X1   g707(.A(new_n908_), .B(G197gat), .Z(G1352gat));
  NOR2_X1   g708(.A1(new_n907_), .A2(new_n672_), .ZN(new_n910_));
  XOR2_X1   g709(.A(new_n910_), .B(G204gat), .Z(G1353gat));
  NOR2_X1   g710(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n912_));
  AND2_X1   g711(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n913_));
  NOR4_X1   g712(.A1(new_n907_), .A2(new_n625_), .A3(new_n912_), .A4(new_n913_), .ZN(new_n914_));
  OR2_X1    g713(.A1(new_n907_), .A2(new_n625_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n914_), .B1(new_n915_), .B2(new_n912_), .ZN(G1354gat));
  OAI21_X1  g715(.A(G218gat), .B1(new_n907_), .B2(new_n604_), .ZN(new_n917_));
  OR2_X1    g716(.A1(new_n637_), .A2(G218gat), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n917_), .B1(new_n907_), .B2(new_n918_), .ZN(new_n919_));
  INV_X1    g718(.A(KEYINPUT126), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n919_), .B(new_n920_), .ZN(G1355gat));
endmodule


