//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 0 1 0 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n662_, new_n663_, new_n664_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n671_, new_n672_,
    new_n673_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n735_, new_n736_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n778_, new_n779_,
    new_n780_, new_n781_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n875_, new_n876_, new_n877_, new_n879_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n927_, new_n928_, new_n929_,
    new_n931_, new_n932_, new_n934_, new_n935_, new_n936_, new_n937_,
    new_n938_, new_n939_, new_n941_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n948_, new_n949_, new_n950_;
  INV_X1    g000(.A(KEYINPUT71), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G120gat), .B(G148gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT5), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G176gat), .B(G204gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  XNOR2_X1  g005(.A(G57gat), .B(G64gat), .ZN(new_n207_));
  OR2_X1    g006(.A1(new_n207_), .A2(KEYINPUT11), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(KEYINPUT11), .ZN(new_n209_));
  XOR2_X1   g008(.A(G71gat), .B(G78gat), .Z(new_n210_));
  NAND3_X1  g009(.A1(new_n208_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n211_));
  OR2_X1    g010(.A1(new_n209_), .A2(new_n210_), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  INV_X1    g012(.A(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(KEYINPUT6), .ZN(new_n215_));
  AOI21_X1  g014(.A(new_n215_), .B1(G99gat), .B2(G106gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(G99gat), .A2(G106gat), .ZN(new_n217_));
  NOR2_X1   g016(.A1(new_n217_), .A2(KEYINPUT6), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT68), .B1(new_n216_), .B2(new_n218_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n217_), .A2(KEYINPUT6), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n215_), .A2(G99gat), .A3(G106gat), .ZN(new_n221_));
  INV_X1    g020(.A(KEYINPUT68), .ZN(new_n222_));
  NAND3_X1  g021(.A1(new_n220_), .A2(new_n221_), .A3(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(G99gat), .ZN(new_n224_));
  INV_X1    g023(.A(G106gat), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n224_), .A2(new_n225_), .A3(KEYINPUT66), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT7), .ZN(new_n227_));
  INV_X1    g026(.A(KEYINPUT7), .ZN(new_n228_));
  NAND4_X1  g027(.A1(new_n228_), .A2(new_n224_), .A3(new_n225_), .A4(KEYINPUT66), .ZN(new_n229_));
  NAND4_X1  g028(.A1(new_n219_), .A2(new_n223_), .A3(new_n227_), .A4(new_n229_), .ZN(new_n230_));
  XOR2_X1   g029(.A(G85gat), .B(G92gat), .Z(new_n231_));
  NAND2_X1  g030(.A1(new_n230_), .A2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT8), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n220_), .A2(new_n221_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n227_), .A2(new_n235_), .A3(new_n229_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT67), .ZN(new_n237_));
  AOI21_X1  g036(.A(new_n234_), .B1(new_n236_), .B2(new_n237_), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n227_), .A2(new_n235_), .A3(KEYINPUT67), .A4(new_n229_), .ZN(new_n239_));
  AOI22_X1  g038(.A1(new_n232_), .A2(KEYINPUT8), .B1(new_n238_), .B2(new_n239_), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT10), .B(G99gat), .ZN(new_n241_));
  OAI21_X1  g040(.A(new_n235_), .B1(new_n241_), .B2(G106gat), .ZN(new_n242_));
  NAND3_X1  g041(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(new_n243_), .B(KEYINPUT65), .Z(new_n244_));
  OAI21_X1  g043(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(KEYINPUT64), .B(G85gat), .ZN(new_n246_));
  INV_X1    g045(.A(G92gat), .ZN(new_n247_));
  OAI21_X1  g046(.A(new_n245_), .B1(new_n246_), .B2(new_n247_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n242_), .B1(new_n244_), .B2(new_n248_), .ZN(new_n249_));
  OAI211_X1 g048(.A(KEYINPUT69), .B(new_n214_), .C1(new_n240_), .C2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G230gat), .A2(G233gat), .ZN(new_n251_));
  INV_X1    g050(.A(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n250_), .A2(new_n252_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(new_n238_), .A2(new_n239_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n231_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n227_), .A2(new_n229_), .ZN(new_n256_));
  AOI21_X1  g055(.A(new_n222_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n257_));
  NOR2_X1   g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n255_), .B1(new_n258_), .B2(new_n223_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n254_), .B1(new_n259_), .B2(new_n233_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n249_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n213_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n262_), .A2(KEYINPUT69), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n236_), .A2(new_n237_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n234_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n264_), .A2(new_n239_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n233_), .B1(new_n230_), .B2(new_n231_), .ZN(new_n267_));
  OAI211_X1 g066(.A(new_n213_), .B(new_n261_), .C1(new_n266_), .C2(new_n267_), .ZN(new_n268_));
  AOI21_X1  g067(.A(new_n253_), .B1(new_n263_), .B2(new_n268_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n214_), .B1(new_n240_), .B2(new_n249_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n270_), .A2(KEYINPUT12), .A3(new_n268_), .ZN(new_n271_));
  OAI21_X1  g070(.A(new_n261_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n272_));
  INV_X1    g071(.A(KEYINPUT12), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n272_), .A2(new_n273_), .A3(new_n214_), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n252_), .B1(new_n271_), .B2(new_n274_), .ZN(new_n275_));
  OAI21_X1  g074(.A(new_n206_), .B1(new_n269_), .B2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n268_), .A2(KEYINPUT12), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(new_n262_), .ZN(new_n278_));
  INV_X1    g077(.A(new_n274_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n251_), .B1(new_n278_), .B2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT69), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n270_), .A2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(new_n268_), .ZN(new_n283_));
  OAI211_X1 g082(.A(new_n252_), .B(new_n250_), .C1(new_n282_), .C2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(new_n206_), .ZN(new_n285_));
  NAND3_X1  g084(.A1(new_n280_), .A2(new_n284_), .A3(new_n285_), .ZN(new_n286_));
  AND3_X1   g085(.A1(new_n276_), .A2(new_n286_), .A3(KEYINPUT70), .ZN(new_n287_));
  AOI21_X1  g086(.A(KEYINPUT70), .B1(new_n276_), .B2(new_n286_), .ZN(new_n288_));
  INV_X1    g087(.A(KEYINPUT13), .ZN(new_n289_));
  NOR3_X1   g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n291_));
  NOR3_X1   g090(.A1(new_n269_), .A2(new_n275_), .A3(new_n206_), .ZN(new_n292_));
  AOI21_X1  g091(.A(new_n285_), .B1(new_n280_), .B2(new_n284_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n291_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n276_), .A2(new_n286_), .A3(KEYINPUT70), .ZN(new_n295_));
  AOI21_X1  g094(.A(KEYINPUT13), .B1(new_n294_), .B2(new_n295_), .ZN(new_n296_));
  OAI21_X1  g095(.A(new_n202_), .B1(new_n290_), .B2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(KEYINPUT77), .ZN(new_n298_));
  XNOR2_X1  g097(.A(G29gat), .B(G36gat), .ZN(new_n299_));
  INV_X1    g098(.A(new_n299_), .ZN(new_n300_));
  XOR2_X1   g099(.A(G43gat), .B(G50gat), .Z(new_n301_));
  NAND2_X1  g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G43gat), .B(G50gat), .ZN(new_n303_));
  NAND2_X1  g102(.A1(new_n299_), .A2(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n302_), .A2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(KEYINPUT15), .ZN(new_n306_));
  XNOR2_X1  g105(.A(G15gat), .B(G22gat), .ZN(new_n307_));
  INV_X1    g106(.A(G1gat), .ZN(new_n308_));
  INV_X1    g107(.A(G8gat), .ZN(new_n309_));
  OAI21_X1  g108(.A(KEYINPUT14), .B1(new_n308_), .B2(new_n309_), .ZN(new_n310_));
  NAND2_X1  g109(.A1(new_n307_), .A2(new_n310_), .ZN(new_n311_));
  XNOR2_X1  g110(.A(G1gat), .B(G8gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n306_), .A2(new_n313_), .ZN(new_n314_));
  INV_X1    g113(.A(new_n305_), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n314_), .A2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(G229gat), .A2(G233gat), .ZN(new_n318_));
  INV_X1    g117(.A(new_n318_), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n298_), .B1(new_n317_), .B2(new_n319_), .ZN(new_n320_));
  NAND4_X1  g119(.A1(new_n314_), .A2(KEYINPUT77), .A3(new_n318_), .A4(new_n316_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT76), .ZN(new_n322_));
  XNOR2_X1  g121(.A(new_n313_), .B(new_n315_), .ZN(new_n323_));
  AOI21_X1  g122(.A(new_n322_), .B1(new_n323_), .B2(new_n319_), .ZN(new_n324_));
  AND3_X1   g123(.A1(new_n323_), .A2(new_n322_), .A3(new_n319_), .ZN(new_n325_));
  OAI211_X1 g124(.A(new_n320_), .B(new_n321_), .C1(new_n324_), .C2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(G113gat), .B(G141gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n327_), .B(KEYINPUT78), .ZN(new_n328_));
  XNOR2_X1  g127(.A(G169gat), .B(G197gat), .ZN(new_n329_));
  XNOR2_X1  g128(.A(new_n328_), .B(new_n329_), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n326_), .B(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n289_), .B1(new_n287_), .B2(new_n288_), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n294_), .A2(KEYINPUT13), .A3(new_n295_), .ZN(new_n333_));
  NAND3_X1  g132(.A1(new_n332_), .A2(new_n333_), .A3(KEYINPUT71), .ZN(new_n334_));
  XOR2_X1   g133(.A(G127gat), .B(G134gat), .Z(new_n335_));
  XOR2_X1   g134(.A(G113gat), .B(G120gat), .Z(new_n336_));
  XNOR2_X1  g135(.A(new_n335_), .B(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XNOR2_X1  g137(.A(G155gat), .B(G162gat), .ZN(new_n339_));
  NOR2_X1   g138(.A1(new_n339_), .A2(KEYINPUT1), .ZN(new_n340_));
  INV_X1    g139(.A(G141gat), .ZN(new_n341_));
  INV_X1    g140(.A(G148gat), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(G141gat), .A2(G148gat), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT1), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G155gat), .A2(G162gat), .ZN(new_n346_));
  OAI211_X1 g145(.A(new_n343_), .B(new_n344_), .C1(new_n345_), .C2(new_n346_), .ZN(new_n347_));
  OR2_X1    g146(.A1(new_n340_), .A2(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT84), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n339_), .A2(new_n349_), .ZN(new_n350_));
  OR2_X1    g149(.A1(G155gat), .A2(G162gat), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n351_), .A2(KEYINPUT84), .A3(new_n346_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT2), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n344_), .A2(new_n353_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n355_));
  NOR3_X1   g154(.A1(KEYINPUT83), .A2(G141gat), .A3(G148gat), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n357_));
  OAI211_X1 g156(.A(new_n354_), .B(new_n355_), .C1(new_n356_), .C2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT83), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n359_), .A2(new_n341_), .A3(new_n342_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(new_n360_), .A2(KEYINPUT3), .ZN(new_n361_));
  OAI211_X1 g160(.A(new_n350_), .B(new_n352_), .C1(new_n358_), .C2(new_n361_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n348_), .A2(new_n362_), .ZN(new_n363_));
  NAND2_X1  g162(.A1(new_n338_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n337_), .A2(new_n348_), .A3(new_n362_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(KEYINPUT4), .A3(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G225gat), .A2(G233gat), .ZN(new_n367_));
  INV_X1    g166(.A(new_n367_), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n338_), .A2(new_n363_), .A3(new_n369_), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n366_), .A2(new_n368_), .A3(new_n370_), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n364_), .A2(new_n365_), .A3(new_n367_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n371_), .A2(new_n372_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G1gat), .B(G29gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(G85gat), .ZN(new_n375_));
  XNOR2_X1  g174(.A(KEYINPUT0), .B(G57gat), .ZN(new_n376_));
  XOR2_X1   g175(.A(new_n375_), .B(new_n376_), .Z(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n373_), .A2(new_n378_), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n371_), .A2(new_n372_), .A3(new_n377_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G226gat), .A2(G233gat), .ZN(new_n382_));
  XNOR2_X1  g181(.A(new_n382_), .B(KEYINPUT19), .ZN(new_n383_));
  NOR2_X1   g182(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(new_n384_), .B(G169gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G183gat), .A2(G190gat), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n386_), .A2(KEYINPUT23), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT23), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n388_), .A2(G183gat), .A3(G190gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n389_), .A3(KEYINPUT81), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n386_), .A2(new_n391_), .A3(KEYINPUT23), .ZN(new_n392_));
  NAND2_X1  g191(.A1(new_n390_), .A2(new_n392_), .ZN(new_n393_));
  NOR2_X1   g192(.A1(G183gat), .A2(G190gat), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n385_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(G183gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n396_), .A2(KEYINPUT25), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT25), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n398_), .A2(G183gat), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT91), .ZN(new_n400_));
  AND3_X1   g199(.A1(new_n397_), .A2(new_n399_), .A3(new_n400_), .ZN(new_n401_));
  AOI21_X1  g200(.A(new_n400_), .B1(new_n397_), .B2(new_n399_), .ZN(new_n402_));
  XOR2_X1   g201(.A(KEYINPUT26), .B(G190gat), .Z(new_n403_));
  NOR3_X1   g202(.A1(new_n401_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n404_));
  INV_X1    g203(.A(KEYINPUT24), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n405_), .B1(G169gat), .B2(G176gat), .ZN(new_n406_));
  NOR2_X1   g205(.A1(G169gat), .A2(G176gat), .ZN(new_n407_));
  INV_X1    g206(.A(KEYINPUT80), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  OAI21_X1  g208(.A(KEYINPUT80), .B1(G169gat), .B2(G176gat), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n406_), .A2(new_n409_), .A3(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(KEYINPUT82), .ZN(new_n412_));
  NAND3_X1  g211(.A1(new_n386_), .A2(new_n412_), .A3(KEYINPUT23), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n387_), .A2(new_n389_), .A3(KEYINPUT82), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n407_), .A2(new_n405_), .ZN(new_n415_));
  NAND4_X1  g214(.A1(new_n411_), .A2(new_n413_), .A3(new_n414_), .A4(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n395_), .B1(new_n404_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(G218gat), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(G211gat), .ZN(new_n419_));
  INV_X1    g218(.A(G211gat), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n420_), .A2(G218gat), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(KEYINPUT21), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G197gat), .B(G204gat), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n422_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT88), .ZN(new_n426_));
  INV_X1    g225(.A(G204gat), .ZN(new_n427_));
  NAND3_X1  g226(.A1(new_n426_), .A2(new_n427_), .A3(G197gat), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(G197gat), .ZN(new_n429_));
  INV_X1    g228(.A(G197gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n430_), .A2(G204gat), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n429_), .A2(new_n431_), .ZN(new_n432_));
  OAI211_X1 g231(.A(KEYINPUT21), .B(new_n428_), .C1(new_n432_), .C2(new_n426_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n425_), .A2(new_n433_), .ZN(new_n434_));
  INV_X1    g233(.A(KEYINPUT89), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n422_), .A2(new_n435_), .ZN(new_n436_));
  NAND3_X1  g235(.A1(new_n419_), .A2(new_n421_), .A3(KEYINPUT89), .ZN(new_n437_));
  NAND4_X1  g236(.A1(new_n436_), .A2(KEYINPUT21), .A3(new_n432_), .A4(new_n437_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n434_), .A2(new_n438_), .ZN(new_n439_));
  OAI21_X1  g238(.A(KEYINPUT20), .B1(new_n417_), .B2(new_n439_), .ZN(new_n440_));
  AND2_X1   g239(.A1(new_n390_), .A2(new_n392_), .ZN(new_n441_));
  INV_X1    g240(.A(KEYINPUT79), .ZN(new_n442_));
  INV_X1    g241(.A(G190gat), .ZN(new_n443_));
  OR3_X1    g242(.A1(new_n442_), .A2(new_n443_), .A3(KEYINPUT26), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT26), .B1(new_n442_), .B2(new_n443_), .ZN(new_n445_));
  NAND4_X1  g244(.A1(new_n444_), .A2(new_n397_), .A3(new_n399_), .A4(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n409_), .A2(new_n410_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n447_), .A2(new_n405_), .ZN(new_n448_));
  NAND4_X1  g247(.A1(new_n441_), .A2(new_n446_), .A3(new_n448_), .A4(new_n411_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n414_), .A2(new_n413_), .ZN(new_n450_));
  OAI21_X1  g249(.A(new_n385_), .B1(new_n450_), .B2(new_n394_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n449_), .A2(new_n451_), .B1(new_n434_), .B2(new_n438_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n383_), .B1(new_n440_), .B2(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G8gat), .B(G36gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT18), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G64gat), .B(G92gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n455_), .B(new_n456_), .ZN(new_n457_));
  AND2_X1   g256(.A1(new_n457_), .A2(KEYINPUT32), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n417_), .A2(new_n439_), .ZN(new_n459_));
  AND3_X1   g258(.A1(new_n437_), .A2(KEYINPUT21), .A3(new_n432_), .ZN(new_n460_));
  AOI22_X1  g259(.A1(new_n436_), .A2(new_n460_), .B1(new_n425_), .B2(new_n433_), .ZN(new_n461_));
  NAND3_X1  g260(.A1(new_n461_), .A2(new_n451_), .A3(new_n449_), .ZN(new_n462_));
  NAND3_X1  g261(.A1(new_n459_), .A2(new_n462_), .A3(KEYINPUT20), .ZN(new_n463_));
  OAI211_X1 g262(.A(new_n453_), .B(new_n458_), .C1(new_n383_), .C2(new_n463_), .ZN(new_n464_));
  NOR3_X1   g263(.A1(new_n440_), .A2(new_n452_), .A3(new_n383_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n383_), .ZN(new_n466_));
  INV_X1    g265(.A(KEYINPUT20), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n467_), .B1(new_n417_), .B2(new_n439_), .ZN(new_n468_));
  AOI21_X1  g267(.A(new_n466_), .B1(new_n468_), .B2(new_n462_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n464_), .B1(new_n470_), .B2(KEYINPUT98), .ZN(new_n471_));
  INV_X1    g270(.A(KEYINPUT98), .ZN(new_n472_));
  AOI21_X1  g271(.A(new_n458_), .B1(new_n470_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n381_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n457_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n475_), .B1(new_n465_), .B2(new_n469_), .ZN(new_n476_));
  NAND2_X1  g275(.A1(new_n463_), .A2(new_n383_), .ZN(new_n477_));
  OAI211_X1 g276(.A(new_n461_), .B(new_n395_), .C1(new_n404_), .C2(new_n416_), .ZN(new_n478_));
  NAND2_X1  g277(.A1(new_n449_), .A2(new_n451_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(new_n439_), .ZN(new_n480_));
  NAND4_X1  g279(.A1(new_n478_), .A2(new_n480_), .A3(KEYINPUT20), .A4(new_n466_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n477_), .A2(new_n457_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT92), .ZN(new_n483_));
  NAND3_X1  g282(.A1(new_n476_), .A2(new_n482_), .A3(new_n483_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n470_), .A2(KEYINPUT92), .A3(new_n457_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n484_), .A2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT94), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n380_), .A2(new_n487_), .ZN(new_n488_));
  NAND4_X1  g287(.A1(new_n371_), .A2(KEYINPUT94), .A3(new_n372_), .A4(new_n377_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT95), .B(KEYINPUT33), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n488_), .A2(new_n489_), .A3(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n486_), .A2(new_n491_), .ZN(new_n492_));
  NAND4_X1  g291(.A1(new_n371_), .A2(KEYINPUT33), .A3(new_n372_), .A4(new_n377_), .ZN(new_n493_));
  OR2_X1    g292(.A1(new_n493_), .A2(KEYINPUT93), .ZN(new_n494_));
  NAND3_X1  g293(.A1(new_n366_), .A2(new_n367_), .A3(new_n370_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n495_), .A2(KEYINPUT97), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n364_), .A2(new_n365_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT96), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n497_), .A2(new_n498_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n364_), .A2(KEYINPUT96), .A3(new_n365_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n499_), .A2(new_n368_), .A3(new_n500_), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT97), .ZN(new_n502_));
  NAND4_X1  g301(.A1(new_n366_), .A2(new_n502_), .A3(new_n367_), .A4(new_n370_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n496_), .A2(new_n501_), .A3(new_n378_), .A4(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n493_), .A2(KEYINPUT93), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n494_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  OAI21_X1  g305(.A(new_n474_), .B1(new_n492_), .B2(new_n506_), .ZN(new_n507_));
  XOR2_X1   g306(.A(KEYINPUT86), .B(KEYINPUT28), .Z(new_n508_));
  INV_X1    g307(.A(KEYINPUT85), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n340_), .A2(new_n347_), .ZN(new_n510_));
  AND2_X1   g309(.A1(new_n350_), .A2(new_n352_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n360_), .A2(KEYINPUT3), .ZN(new_n512_));
  NAND2_X1  g311(.A1(new_n356_), .A2(new_n357_), .ZN(new_n513_));
  NAND4_X1  g312(.A1(new_n512_), .A2(new_n513_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n514_));
  AOI21_X1  g313(.A(new_n510_), .B1(new_n511_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT29), .ZN(new_n516_));
  AOI21_X1  g315(.A(new_n509_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  AND4_X1   g316(.A1(new_n509_), .A2(new_n348_), .A3(new_n362_), .A4(new_n516_), .ZN(new_n518_));
  OAI21_X1  g317(.A(new_n508_), .B1(new_n517_), .B2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NOR2_X1   g320(.A1(KEYINPUT87), .A2(G233gat), .ZN(new_n522_));
  OAI21_X1  g321(.A(G228gat), .B1(new_n521_), .B2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  XNOR2_X1  g323(.A(KEYINPUT90), .B(KEYINPUT29), .ZN(new_n525_));
  AOI21_X1  g324(.A(new_n525_), .B1(new_n348_), .B2(new_n362_), .ZN(new_n526_));
  OAI21_X1  g325(.A(new_n524_), .B1(new_n526_), .B2(new_n461_), .ZN(new_n527_));
  OAI211_X1 g326(.A(new_n439_), .B(new_n523_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  OAI21_X1  g328(.A(KEYINPUT85), .B1(new_n363_), .B2(KEYINPUT29), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n515_), .A2(new_n509_), .A3(new_n516_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n508_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n530_), .A2(new_n531_), .A3(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n519_), .A2(new_n529_), .A3(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n529_), .B1(new_n519_), .B2(new_n533_), .ZN(new_n535_));
  XNOR2_X1  g334(.A(G78gat), .B(G106gat), .ZN(new_n536_));
  XNOR2_X1  g335(.A(G22gat), .B(G50gat), .ZN(new_n537_));
  XNOR2_X1  g336(.A(new_n536_), .B(new_n537_), .ZN(new_n538_));
  INV_X1    g337(.A(new_n538_), .ZN(new_n539_));
  NOR3_X1   g338(.A1(new_n534_), .A2(new_n535_), .A3(new_n539_), .ZN(new_n540_));
  AND2_X1   g339(.A1(new_n527_), .A2(new_n528_), .ZN(new_n541_));
  INV_X1    g340(.A(new_n533_), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n532_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n543_));
  OAI21_X1  g342(.A(new_n541_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n519_), .A2(new_n529_), .A3(new_n533_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n538_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(G71gat), .B(G99gat), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n547_), .B(G43gat), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n449_), .A2(new_n451_), .A3(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  AOI21_X1  g349(.A(new_n548_), .B1(new_n449_), .B2(new_n451_), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n338_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(G227gat), .A2(G233gat), .ZN(new_n553_));
  INV_X1    g352(.A(G15gat), .ZN(new_n554_));
  XNOR2_X1  g353(.A(new_n553_), .B(new_n554_), .ZN(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT30), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n556_), .B(KEYINPUT31), .ZN(new_n557_));
  INV_X1    g356(.A(new_n548_), .ZN(new_n558_));
  NAND2_X1  g357(.A1(new_n479_), .A2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n559_), .A2(new_n337_), .A3(new_n549_), .ZN(new_n560_));
  AND3_X1   g359(.A1(new_n552_), .A2(new_n557_), .A3(new_n560_), .ZN(new_n561_));
  AOI21_X1  g360(.A(new_n557_), .B1(new_n552_), .B2(new_n560_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n561_), .A2(new_n562_), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n540_), .A2(new_n546_), .A3(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n507_), .A2(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n563_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n566_), .B1(new_n540_), .B2(new_n546_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n539_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n544_), .A2(new_n538_), .A3(new_n545_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n568_), .A2(new_n569_), .A3(new_n563_), .ZN(new_n570_));
  NAND2_X1  g369(.A1(new_n567_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT27), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n484_), .A2(new_n572_), .A3(new_n485_), .ZN(new_n573_));
  XOR2_X1   g372(.A(new_n457_), .B(KEYINPUT99), .Z(new_n574_));
  OAI21_X1  g373(.A(new_n453_), .B1(new_n383_), .B2(new_n463_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n574_), .A2(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n576_), .A2(KEYINPUT27), .A3(new_n482_), .ZN(new_n577_));
  AND2_X1   g376(.A1(new_n573_), .A2(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n381_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n571_), .A2(new_n578_), .A3(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n565_), .A2(new_n580_), .ZN(new_n581_));
  NAND4_X1  g380(.A1(new_n297_), .A2(new_n331_), .A3(new_n334_), .A4(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT34), .Z(new_n584_));
  INV_X1    g383(.A(KEYINPUT35), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n584_), .A2(new_n585_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  NAND2_X1  g386(.A1(new_n272_), .A2(new_n306_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT73), .ZN(new_n589_));
  AOI21_X1  g388(.A(new_n587_), .B1(new_n588_), .B2(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n232_), .A2(KEYINPUT8), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n249_), .B1(new_n591_), .B2(new_n254_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n592_), .A2(new_n305_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n584_), .A2(new_n585_), .ZN(new_n594_));
  XOR2_X1   g393(.A(new_n594_), .B(KEYINPUT72), .Z(new_n595_));
  NAND3_X1  g394(.A1(new_n593_), .A2(new_n588_), .A3(new_n595_), .ZN(new_n596_));
  AND2_X1   g395(.A1(new_n590_), .A2(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n590_), .A2(new_n596_), .ZN(new_n598_));
  XNOR2_X1  g397(.A(G190gat), .B(G218gat), .ZN(new_n599_));
  XNOR2_X1  g398(.A(G134gat), .B(G162gat), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n599_), .B(new_n600_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n601_), .A2(KEYINPUT36), .ZN(new_n602_));
  INV_X1    g401(.A(new_n602_), .ZN(new_n603_));
  NOR3_X1   g402(.A1(new_n597_), .A2(new_n598_), .A3(new_n603_), .ZN(new_n604_));
  XOR2_X1   g403(.A(new_n601_), .B(KEYINPUT36), .Z(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  OR2_X1    g405(.A1(new_n590_), .A2(new_n596_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n590_), .A2(new_n596_), .ZN(new_n608_));
  AOI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(KEYINPUT37), .B1(new_n604_), .B2(new_n609_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n605_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT37), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n607_), .A2(new_n608_), .ZN(new_n613_));
  OAI211_X1 g412(.A(new_n611_), .B(new_n612_), .C1(new_n613_), .C2(new_n603_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n610_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n313_), .B(new_n616_), .ZN(new_n617_));
  XNOR2_X1  g416(.A(new_n617_), .B(new_n213_), .ZN(new_n618_));
  XOR2_X1   g417(.A(G127gat), .B(G155gat), .Z(new_n619_));
  XNOR2_X1  g418(.A(new_n619_), .B(KEYINPUT16), .ZN(new_n620_));
  XNOR2_X1  g419(.A(G183gat), .B(G211gat), .ZN(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT17), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n618_), .A2(new_n623_), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n624_), .B(KEYINPUT75), .ZN(new_n625_));
  OR2_X1    g424(.A1(new_n618_), .A2(KEYINPUT74), .ZN(new_n626_));
  NAND2_X1  g425(.A1(new_n618_), .A2(KEYINPUT74), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT17), .ZN(new_n628_));
  NOR2_X1   g427(.A1(new_n622_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n626_), .A2(new_n627_), .A3(new_n629_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n625_), .A2(new_n630_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n615_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n632_), .ZN(new_n633_));
  NOR2_X1   g432(.A1(new_n582_), .A2(new_n633_), .ZN(new_n634_));
  NAND3_X1  g433(.A1(new_n634_), .A2(new_n308_), .A3(new_n381_), .ZN(new_n635_));
  INV_X1    g434(.A(KEYINPUT38), .ZN(new_n636_));
  OR2_X1    g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  AND3_X1   g436(.A1(new_n297_), .A2(new_n331_), .A3(new_n334_), .ZN(new_n638_));
  OAI21_X1  g437(.A(new_n611_), .B1(new_n613_), .B2(new_n603_), .ZN(new_n639_));
  INV_X1    g438(.A(new_n639_), .ZN(new_n640_));
  AOI211_X1 g439(.A(new_n631_), .B(new_n640_), .C1(new_n565_), .C2(new_n580_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n638_), .A2(new_n641_), .ZN(new_n642_));
  OAI21_X1  g441(.A(G1gat), .B1(new_n642_), .B2(new_n579_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n635_), .A2(new_n636_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n637_), .A2(new_n643_), .A3(new_n644_), .ZN(G1324gat));
  NAND2_X1  g444(.A1(new_n573_), .A2(new_n577_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n634_), .A2(new_n309_), .A3(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n638_), .A2(new_n646_), .A3(new_n641_), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT100), .ZN(new_n649_));
  NOR2_X1   g448(.A1(new_n649_), .A2(KEYINPUT39), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n309_), .B1(new_n649_), .B2(KEYINPUT39), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n648_), .A2(new_n650_), .A3(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n650_), .B1(new_n648_), .B2(new_n651_), .ZN(new_n654_));
  OAI21_X1  g453(.A(new_n647_), .B1(new_n653_), .B2(new_n654_), .ZN(new_n655_));
  OR2_X1    g454(.A1(new_n655_), .A2(KEYINPUT102), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(KEYINPUT102), .ZN(new_n657_));
  XNOR2_X1  g456(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n658_));
  AND3_X1   g457(.A1(new_n656_), .A2(new_n657_), .A3(new_n658_), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n658_), .B1(new_n656_), .B2(new_n657_), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n659_), .A2(new_n660_), .ZN(G1325gat));
  OAI21_X1  g460(.A(G15gat), .B1(new_n642_), .B2(new_n566_), .ZN(new_n662_));
  XOR2_X1   g461(.A(new_n662_), .B(KEYINPUT41), .Z(new_n663_));
  NAND3_X1  g462(.A1(new_n634_), .A2(new_n554_), .A3(new_n563_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n663_), .A2(new_n664_), .ZN(G1326gat));
  NOR2_X1   g464(.A1(new_n540_), .A2(new_n546_), .ZN(new_n666_));
  OAI21_X1  g465(.A(G22gat), .B1(new_n642_), .B2(new_n666_), .ZN(new_n667_));
  XNOR2_X1  g466(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n668_));
  XNOR2_X1  g467(.A(new_n667_), .B(new_n668_), .ZN(new_n669_));
  INV_X1    g468(.A(G22gat), .ZN(new_n670_));
  INV_X1    g469(.A(new_n666_), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n634_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n669_), .A2(new_n672_), .ZN(new_n673_));
  XOR2_X1   g472(.A(new_n673_), .B(KEYINPUT104), .Z(G1327gat));
  INV_X1    g473(.A(new_n631_), .ZN(new_n675_));
  NOR2_X1   g474(.A1(new_n675_), .A2(new_n639_), .ZN(new_n676_));
  INV_X1    g475(.A(new_n676_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n582_), .A2(new_n677_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n679_), .A2(G29gat), .A3(new_n579_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681_));
  NAND4_X1  g480(.A1(new_n297_), .A2(new_n631_), .A3(new_n331_), .A4(new_n334_), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT105), .ZN(new_n683_));
  INV_X1    g482(.A(KEYINPUT107), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n610_), .A2(new_n614_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n565_), .B2(new_n580_), .ZN(new_n686_));
  OAI211_X1 g485(.A(new_n684_), .B(KEYINPUT43), .C1(new_n686_), .C2(KEYINPUT106), .ZN(new_n687_));
  AND3_X1   g486(.A1(new_n568_), .A2(new_n563_), .A3(new_n569_), .ZN(new_n688_));
  AOI21_X1  g487(.A(new_n563_), .B1(new_n568_), .B2(new_n569_), .ZN(new_n689_));
  OAI21_X1  g488(.A(new_n579_), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NOR2_X1   g489(.A1(new_n690_), .A2(new_n646_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n666_), .A2(new_n566_), .ZN(new_n692_));
  AND2_X1   g491(.A1(new_n504_), .A2(new_n505_), .ZN(new_n693_));
  NAND4_X1  g492(.A1(new_n693_), .A2(new_n486_), .A3(new_n494_), .A4(new_n491_), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n692_), .B1(new_n694_), .B2(new_n474_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n615_), .B1(new_n691_), .B2(new_n695_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT106), .ZN(new_n697_));
  AOI21_X1  g496(.A(KEYINPUT107), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n699_), .B1(new_n686_), .B2(new_n684_), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n687_), .B1(new_n698_), .B2(new_n700_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n681_), .B1(new_n683_), .B2(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n703_));
  XNOR2_X1  g502(.A(new_n682_), .B(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n701_), .ZN(new_n705_));
  NAND3_X1  g504(.A1(new_n704_), .A2(new_n705_), .A3(KEYINPUT44), .ZN(new_n706_));
  AND2_X1   g505(.A1(new_n702_), .A2(new_n706_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n707_), .A2(KEYINPUT108), .A3(new_n381_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(G29gat), .ZN(new_n709_));
  AOI21_X1  g508(.A(KEYINPUT108), .B1(new_n707_), .B2(new_n381_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n680_), .B1(new_n709_), .B2(new_n710_), .ZN(G1328gat));
  INV_X1    g510(.A(KEYINPUT110), .ZN(new_n712_));
  INV_X1    g511(.A(KEYINPUT46), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n712_), .A2(new_n713_), .ZN(new_n714_));
  NOR2_X1   g513(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n702_), .A2(new_n646_), .A3(new_n706_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n716_), .A2(G36gat), .ZN(new_n717_));
  NOR2_X1   g516(.A1(new_n578_), .A2(G36gat), .ZN(new_n718_));
  NAND4_X1  g517(.A1(new_n638_), .A2(new_n581_), .A3(new_n676_), .A4(new_n718_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT109), .ZN(new_n720_));
  INV_X1    g519(.A(KEYINPUT109), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n678_), .A2(new_n721_), .A3(new_n718_), .ZN(new_n722_));
  AND3_X1   g521(.A1(new_n720_), .A2(KEYINPUT45), .A3(new_n722_), .ZN(new_n723_));
  AOI21_X1  g522(.A(KEYINPUT45), .B1(new_n720_), .B2(new_n722_), .ZN(new_n724_));
  NOR2_X1   g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  AOI211_X1 g524(.A(new_n714_), .B(new_n715_), .C1(new_n717_), .C2(new_n725_), .ZN(new_n726_));
  AND4_X1   g525(.A1(new_n712_), .A2(new_n717_), .A3(new_n713_), .A4(new_n725_), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(new_n727_), .ZN(G1329gat));
  NAND3_X1  g527(.A1(new_n702_), .A2(new_n563_), .A3(new_n706_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n729_), .A2(G43gat), .ZN(new_n730_));
  OR3_X1    g529(.A1(new_n679_), .A2(G43gat), .A3(new_n566_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(new_n732_));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n732_), .B(new_n733_), .ZN(G1330gat));
  AOI21_X1  g533(.A(G50gat), .B1(new_n678_), .B2(new_n671_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n671_), .A2(G50gat), .ZN(new_n736_));
  AOI21_X1  g535(.A(new_n735_), .B1(new_n707_), .B2(new_n736_), .ZN(G1331gat));
  AND2_X1   g536(.A1(new_n297_), .A2(new_n334_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n738_), .A2(new_n331_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n739_), .A2(new_n641_), .ZN(new_n740_));
  INV_X1    g539(.A(G57gat), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n740_), .A2(new_n741_), .A3(new_n579_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n739_), .A2(new_n581_), .ZN(new_n743_));
  OR3_X1    g542(.A1(new_n743_), .A2(KEYINPUT111), .A3(new_n633_), .ZN(new_n744_));
  OAI21_X1  g543(.A(KEYINPUT111), .B1(new_n743_), .B2(new_n633_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n744_), .A2(new_n381_), .A3(new_n745_), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n742_), .B1(new_n746_), .B2(new_n741_), .ZN(G1332gat));
  NOR2_X1   g546(.A1(new_n743_), .A2(new_n633_), .ZN(new_n748_));
  INV_X1    g547(.A(G64gat), .ZN(new_n749_));
  NAND3_X1  g548(.A1(new_n748_), .A2(new_n749_), .A3(new_n646_), .ZN(new_n750_));
  INV_X1    g549(.A(new_n740_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n751_), .A2(new_n646_), .ZN(new_n752_));
  XOR2_X1   g551(.A(KEYINPUT112), .B(KEYINPUT48), .Z(new_n753_));
  AND3_X1   g552(.A1(new_n752_), .A2(G64gat), .A3(new_n753_), .ZN(new_n754_));
  AOI21_X1  g553(.A(new_n753_), .B1(new_n752_), .B2(G64gat), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n750_), .B1(new_n754_), .B2(new_n755_), .ZN(G1333gat));
  INV_X1    g555(.A(G71gat), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n748_), .A2(new_n757_), .A3(new_n563_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G71gat), .B1(new_n740_), .B2(new_n566_), .ZN(new_n759_));
  AND2_X1   g558(.A1(new_n759_), .A2(KEYINPUT49), .ZN(new_n760_));
  NOR2_X1   g559(.A1(new_n759_), .A2(KEYINPUT49), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n758_), .B1(new_n760_), .B2(new_n761_), .ZN(G1334gat));
  INV_X1    g561(.A(G78gat), .ZN(new_n763_));
  NAND3_X1  g562(.A1(new_n748_), .A2(new_n763_), .A3(new_n671_), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n751_), .A2(new_n671_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n765_), .B1(new_n766_), .B2(G78gat), .ZN(new_n767_));
  AOI211_X1 g566(.A(KEYINPUT50), .B(new_n763_), .C1(new_n751_), .C2(new_n671_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n764_), .B1(new_n767_), .B2(new_n768_), .ZN(G1335gat));
  NAND3_X1  g568(.A1(new_n705_), .A2(new_n631_), .A3(new_n739_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n770_), .A2(new_n246_), .A3(new_n579_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n743_), .A2(new_n677_), .ZN(new_n772_));
  AOI21_X1  g571(.A(G85gat), .B1(new_n772_), .B2(new_n381_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n771_), .A2(new_n773_), .ZN(G1336gat));
  OAI21_X1  g573(.A(G92gat), .B1(new_n770_), .B2(new_n578_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n772_), .A2(new_n247_), .A3(new_n646_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n775_), .A2(new_n776_), .ZN(G1337gat));
  OAI21_X1  g576(.A(G99gat), .B1(new_n770_), .B2(new_n566_), .ZN(new_n778_));
  NOR2_X1   g577(.A1(new_n566_), .A2(new_n241_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n772_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  XNOR2_X1  g580(.A(new_n781_), .B(KEYINPUT51), .ZN(G1338gat));
  XNOR2_X1  g581(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT52), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n705_), .A2(new_n631_), .A3(new_n671_), .A4(new_n739_), .ZN(new_n785_));
  AOI21_X1  g584(.A(new_n784_), .B1(new_n785_), .B2(G106gat), .ZN(new_n786_));
  INV_X1    g585(.A(new_n786_), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n785_), .A2(new_n784_), .A3(G106gat), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n772_), .A2(new_n225_), .A3(new_n671_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n783_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n788_), .ZN(new_n792_));
  OAI211_X1 g591(.A(new_n790_), .B(new_n783_), .C1(new_n792_), .C2(new_n786_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NOR2_X1   g593(.A1(new_n791_), .A2(new_n794_), .ZN(G1339gat));
  NAND2_X1  g594(.A1(new_n331_), .A2(G113gat), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n631_), .A2(new_n331_), .ZN(new_n797_));
  NAND3_X1  g596(.A1(new_n332_), .A2(new_n797_), .A3(new_n333_), .ZN(new_n798_));
  OR2_X1    g597(.A1(new_n798_), .A2(KEYINPUT114), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n798_), .A2(KEYINPUT114), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n799_), .A2(new_n685_), .A3(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(KEYINPUT54), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803_));
  NAND4_X1  g602(.A1(new_n799_), .A2(new_n803_), .A3(new_n685_), .A4(new_n800_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n323_), .A2(new_n318_), .ZN(new_n806_));
  OAI211_X1 g605(.A(new_n330_), .B(new_n806_), .C1(new_n317_), .C2(new_n318_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n807_), .B1(new_n326_), .B2(new_n330_), .ZN(new_n808_));
  INV_X1    g607(.A(KEYINPUT116), .ZN(new_n809_));
  OR2_X1    g608(.A1(new_n808_), .A2(new_n809_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n808_), .A2(new_n809_), .ZN(new_n811_));
  AOI21_X1  g610(.A(new_n292_), .B1(new_n810_), .B2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n280_), .A2(KEYINPUT115), .A3(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT115), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n815_), .B1(new_n275_), .B2(KEYINPUT55), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n275_), .A2(KEYINPUT55), .ZN(new_n817_));
  NAND3_X1  g616(.A1(new_n271_), .A2(new_n252_), .A3(new_n274_), .ZN(new_n818_));
  NAND4_X1  g617(.A1(new_n814_), .A2(new_n816_), .A3(new_n817_), .A4(new_n818_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n819_), .A2(KEYINPUT56), .A3(new_n206_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n820_), .ZN(new_n821_));
  AOI21_X1  g620(.A(KEYINPUT56), .B1(new_n819_), .B2(new_n206_), .ZN(new_n822_));
  OAI21_X1  g621(.A(new_n812_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(KEYINPUT58), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n685_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  OAI211_X1 g624(.A(new_n812_), .B(KEYINPUT58), .C1(new_n822_), .C2(new_n821_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n825_), .A2(new_n826_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n331_), .A2(new_n286_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n819_), .A2(new_n206_), .ZN(new_n829_));
  INV_X1    g628(.A(KEYINPUT56), .ZN(new_n830_));
  NAND2_X1  g629(.A1(new_n829_), .A2(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n828_), .B1(new_n831_), .B2(new_n820_), .ZN(new_n832_));
  AOI22_X1  g631(.A1(new_n810_), .A2(new_n811_), .B1(new_n294_), .B2(new_n295_), .ZN(new_n833_));
  OAI211_X1 g632(.A(KEYINPUT57), .B(new_n639_), .C1(new_n832_), .C2(new_n833_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n827_), .A2(new_n834_), .ZN(new_n835_));
  OAI211_X1 g634(.A(new_n331_), .B(new_n286_), .C1(new_n821_), .C2(new_n822_), .ZN(new_n836_));
  INV_X1    g635(.A(new_n833_), .ZN(new_n837_));
  AOI21_X1  g636(.A(new_n640_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n838_));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839_));
  NAND2_X1  g638(.A1(new_n838_), .A2(new_n839_), .ZN(new_n840_));
  XOR2_X1   g639(.A(KEYINPUT118), .B(KEYINPUT57), .Z(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  OAI21_X1  g641(.A(new_n639_), .B1(new_n832_), .B2(new_n833_), .ZN(new_n843_));
  AOI21_X1  g642(.A(new_n842_), .B1(new_n843_), .B2(KEYINPUT117), .ZN(new_n844_));
  AOI21_X1  g643(.A(new_n835_), .B1(new_n840_), .B2(new_n844_), .ZN(new_n845_));
  OAI21_X1  g644(.A(new_n805_), .B1(new_n845_), .B2(new_n675_), .ZN(new_n846_));
  NOR2_X1   g645(.A1(new_n646_), .A2(new_n579_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  NOR2_X1   g647(.A1(new_n848_), .A2(new_n570_), .ZN(new_n849_));
  NAND4_X1  g648(.A1(new_n846_), .A2(KEYINPUT120), .A3(KEYINPUT59), .A4(new_n849_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n844_), .A2(new_n840_), .ZN(new_n851_));
  AOI22_X1  g650(.A1(new_n838_), .A2(KEYINPUT57), .B1(new_n825_), .B2(new_n826_), .ZN(new_n852_));
  AOI21_X1  g651(.A(new_n675_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  AND2_X1   g652(.A1(new_n802_), .A2(new_n804_), .ZN(new_n854_));
  OAI211_X1 g653(.A(KEYINPUT120), .B(new_n849_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n855_));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n796_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n858_));
  OAI211_X1 g657(.A(new_n331_), .B(new_n849_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n859_));
  INV_X1    g658(.A(G113gat), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n859_), .A2(KEYINPUT119), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT119), .B1(new_n859_), .B2(new_n860_), .ZN(new_n862_));
  NOR3_X1   g661(.A1(new_n858_), .A2(new_n861_), .A3(new_n862_), .ZN(G1340gat));
  NOR2_X1   g662(.A1(new_n853_), .A2(new_n854_), .ZN(new_n864_));
  NOR3_X1   g663(.A1(new_n864_), .A2(new_n570_), .A3(new_n848_), .ZN(new_n865_));
  XOR2_X1   g664(.A(KEYINPUT121), .B(G120gat), .Z(new_n866_));
  OAI21_X1  g665(.A(new_n866_), .B1(new_n738_), .B2(KEYINPUT60), .ZN(new_n867_));
  OAI211_X1 g666(.A(new_n865_), .B(new_n867_), .C1(KEYINPUT60), .C2(new_n866_), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n738_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n866_), .ZN(G1341gat));
  INV_X1    g669(.A(G127gat), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n865_), .A2(new_n871_), .A3(new_n675_), .ZN(new_n872_));
  AOI21_X1  g671(.A(new_n631_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n873_), .B2(new_n871_), .ZN(G1342gat));
  INV_X1    g673(.A(G134gat), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n865_), .A2(new_n875_), .A3(new_n640_), .ZN(new_n876_));
  AOI21_X1  g675(.A(new_n685_), .B1(new_n850_), .B2(new_n857_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n876_), .B1(new_n877_), .B2(new_n875_), .ZN(G1343gat));
  NAND2_X1  g677(.A1(new_n847_), .A2(new_n689_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(KEYINPUT122), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n864_), .A2(new_n881_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n882_), .A2(new_n331_), .ZN(new_n883_));
  XNOR2_X1  g682(.A(new_n883_), .B(G141gat), .ZN(G1344gat));
  INV_X1    g683(.A(new_n738_), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n882_), .A2(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(new_n886_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n888_));
  NAND4_X1  g687(.A1(new_n846_), .A2(new_n888_), .A3(new_n675_), .A4(new_n880_), .ZN(new_n889_));
  OAI211_X1 g688(.A(new_n675_), .B(new_n880_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n890_), .A2(KEYINPUT123), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT61), .B(G155gat), .ZN(new_n893_));
  INV_X1    g692(.A(new_n893_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n892_), .A2(new_n894_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n889_), .A2(new_n891_), .A3(new_n893_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n896_), .ZN(G1346gat));
  OAI211_X1 g696(.A(new_n615_), .B(new_n880_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n898_), .A2(G162gat), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n846_), .A2(new_n880_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n639_), .A2(G162gat), .ZN(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n899_), .B1(new_n900_), .B2(new_n902_), .ZN(new_n903_));
  INV_X1    g702(.A(KEYINPUT124), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n903_), .A2(new_n904_), .ZN(new_n905_));
  OAI211_X1 g704(.A(new_n899_), .B(KEYINPUT124), .C1(new_n900_), .C2(new_n902_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n905_), .A2(new_n906_), .ZN(G1347gat));
  INV_X1    g706(.A(KEYINPUT125), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n578_), .A2(new_n381_), .A3(new_n570_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n909_), .ZN(new_n910_));
  OAI21_X1  g709(.A(new_n908_), .B1(new_n864_), .B2(new_n910_), .ZN(new_n911_));
  OAI211_X1 g710(.A(KEYINPUT125), .B(new_n909_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n911_), .A2(new_n912_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT22), .B(G169gat), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n331_), .A2(new_n915_), .ZN(new_n916_));
  OAI211_X1 g715(.A(new_n331_), .B(new_n909_), .C1(new_n853_), .C2(new_n854_), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918_));
  AND3_X1   g717(.A1(new_n917_), .A2(new_n918_), .A3(G169gat), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n918_), .B1(new_n917_), .B2(G169gat), .ZN(new_n920_));
  OAI22_X1  g719(.A1(new_n914_), .A2(new_n916_), .B1(new_n919_), .B2(new_n920_), .ZN(G1348gat));
  NOR2_X1   g720(.A1(new_n864_), .A2(new_n910_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n885_), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n923_), .A2(G176gat), .ZN(new_n924_));
  OR2_X1    g723(.A1(new_n738_), .A2(G176gat), .ZN(new_n925_));
  OAI21_X1  g724(.A(new_n924_), .B1(new_n914_), .B2(new_n925_), .ZN(G1349gat));
  AOI21_X1  g725(.A(G183gat), .B1(new_n922_), .B2(new_n675_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n401_), .A2(new_n402_), .ZN(new_n928_));
  NOR2_X1   g727(.A1(new_n631_), .A2(new_n928_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n927_), .B1(new_n913_), .B2(new_n929_), .ZN(G1350gat));
  OR2_X1    g729(.A1(new_n639_), .A2(new_n403_), .ZN(new_n931_));
  AOI21_X1  g730(.A(new_n685_), .B1(new_n911_), .B2(new_n912_), .ZN(new_n932_));
  OAI22_X1  g731(.A1(new_n914_), .A2(new_n931_), .B1(new_n932_), .B2(new_n443_), .ZN(G1351gat));
  NAND2_X1  g732(.A1(new_n689_), .A2(new_n579_), .ZN(new_n934_));
  INV_X1    g733(.A(new_n934_), .ZN(new_n935_));
  AOI21_X1  g734(.A(new_n578_), .B1(new_n935_), .B2(KEYINPUT126), .ZN(new_n936_));
  OAI21_X1  g735(.A(new_n936_), .B1(KEYINPUT126), .B2(new_n935_), .ZN(new_n937_));
  NOR2_X1   g736(.A1(new_n864_), .A2(new_n937_), .ZN(new_n938_));
  NAND2_X1  g737(.A1(new_n938_), .A2(new_n331_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(new_n939_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g739(.A1(new_n938_), .A2(new_n885_), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n941_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g741(.A(KEYINPUT63), .B(G211gat), .ZN(new_n943_));
  NOR4_X1   g742(.A1(new_n864_), .A2(new_n631_), .A3(new_n937_), .A4(new_n943_), .ZN(new_n944_));
  NAND2_X1  g743(.A1(new_n938_), .A2(new_n675_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n946_));
  AOI21_X1  g745(.A(new_n944_), .B1(new_n945_), .B2(new_n946_), .ZN(G1354gat));
  AOI21_X1  g746(.A(G218gat), .B1(new_n938_), .B2(new_n640_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n685_), .A2(new_n418_), .ZN(new_n949_));
  XNOR2_X1  g748(.A(new_n949_), .B(KEYINPUT127), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n948_), .B1(new_n938_), .B2(new_n950_), .ZN(G1355gat));
endmodule


