//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n751_,
    new_n752_, new_n753_, new_n755_, new_n756_, new_n757_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n770_, new_n771_, new_n773_,
    new_n774_, new_n775_, new_n776_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n871_, new_n873_,
    new_n874_, new_n876_, new_n877_, new_n878_, new_n880_, new_n881_,
    new_n882_, new_n883_, new_n884_, new_n885_, new_n887_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n895_, new_n896_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n917_,
    new_n918_, new_n919_, new_n920_, new_n922_, new_n923_, new_n924_,
    new_n925_, new_n926_, new_n927_, new_n928_, new_n930_, new_n931_,
    new_n932_, new_n933_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_;
  INV_X1    g000(.A(KEYINPUT7), .ZN(new_n202_));
  INV_X1    g001(.A(G99gat), .ZN(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n202_), .A2(new_n203_), .A3(new_n204_), .ZN(new_n205_));
  NAND2_X1  g004(.A1(G99gat), .A2(G106gat), .ZN(new_n206_));
  INV_X1    g005(.A(KEYINPUT6), .ZN(new_n207_));
  NAND2_X1  g006(.A1(new_n206_), .A2(new_n207_), .ZN(new_n208_));
  NAND3_X1  g007(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n209_));
  OAI21_X1  g008(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n210_));
  NAND4_X1  g009(.A1(new_n205_), .A2(new_n208_), .A3(new_n209_), .A4(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(G85gat), .ZN(new_n212_));
  INV_X1    g011(.A(G92gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(G85gat), .A2(G92gat), .ZN(new_n215_));
  AND2_X1   g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n211_), .A2(new_n216_), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT8), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AND2_X1   g018(.A1(new_n203_), .A2(KEYINPUT10), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n203_), .A2(KEYINPUT10), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n204_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n222_));
  AND2_X1   g021(.A1(new_n208_), .A2(new_n209_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n214_), .A2(KEYINPUT9), .A3(new_n215_), .ZN(new_n224_));
  OR2_X1    g023(.A1(new_n215_), .A2(KEYINPUT9), .ZN(new_n225_));
  NAND4_X1  g024(.A1(new_n222_), .A2(new_n223_), .A3(new_n224_), .A4(new_n225_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n211_), .A2(KEYINPUT8), .A3(new_n216_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n219_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  XOR2_X1   g027(.A(G71gat), .B(G78gat), .Z(new_n229_));
  AND2_X1   g028(.A1(G57gat), .A2(G64gat), .ZN(new_n230_));
  NOR2_X1   g029(.A1(G57gat), .A2(G64gat), .ZN(new_n231_));
  OAI21_X1  g030(.A(KEYINPUT11), .B1(new_n230_), .B2(new_n231_), .ZN(new_n232_));
  INV_X1    g031(.A(G57gat), .ZN(new_n233_));
  INV_X1    g032(.A(G64gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT11), .ZN(new_n236_));
  NAND2_X1  g035(.A1(G57gat), .A2(G64gat), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n235_), .A2(new_n236_), .A3(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n229_), .A2(new_n232_), .A3(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G71gat), .B(G78gat), .ZN(new_n240_));
  OAI211_X1 g039(.A(new_n240_), .B(KEYINPUT11), .C1(new_n231_), .C2(new_n230_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n239_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(new_n242_), .ZN(new_n243_));
  XNOR2_X1  g042(.A(KEYINPUT67), .B(KEYINPUT12), .ZN(new_n244_));
  AND3_X1   g043(.A1(new_n228_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n245_));
  AOI22_X1  g044(.A1(new_n228_), .A2(new_n243_), .B1(KEYINPUT67), .B2(KEYINPUT12), .ZN(new_n246_));
  NOR2_X1   g045(.A1(new_n245_), .A2(new_n246_), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT68), .ZN(new_n248_));
  NAND4_X1  g047(.A1(new_n219_), .A2(new_n242_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(G230gat), .A2(G233gat), .ZN(new_n250_));
  XNOR2_X1  g049(.A(new_n250_), .B(KEYINPUT64), .ZN(new_n251_));
  NAND4_X1  g050(.A1(new_n247_), .A2(new_n248_), .A3(new_n249_), .A4(new_n251_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n228_), .A2(new_n243_), .ZN(new_n253_));
  NAND2_X1  g052(.A1(KEYINPUT67), .A2(KEYINPUT12), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n253_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n228_), .A2(new_n243_), .A3(new_n244_), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n255_), .A2(new_n249_), .A3(new_n251_), .A4(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT68), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n252_), .A2(new_n258_), .ZN(new_n259_));
  INV_X1    g058(.A(new_n251_), .ZN(new_n260_));
  INV_X1    g059(.A(new_n227_), .ZN(new_n261_));
  AOI21_X1  g060(.A(KEYINPUT8), .B1(new_n211_), .B2(new_n216_), .ZN(new_n262_));
  NOR2_X1   g061(.A1(new_n261_), .A2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT65), .ZN(new_n264_));
  NAND4_X1  g063(.A1(new_n263_), .A2(new_n264_), .A3(new_n226_), .A4(new_n242_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n249_), .A2(KEYINPUT65), .ZN(new_n266_));
  NAND3_X1  g065(.A1(new_n265_), .A2(new_n266_), .A3(KEYINPUT66), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n253_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT66), .B1(new_n265_), .B2(new_n266_), .ZN(new_n269_));
  OAI21_X1  g068(.A(new_n260_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n259_), .A2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(G120gat), .B(G148gat), .ZN(new_n272_));
  XNOR2_X1  g071(.A(new_n272_), .B(G204gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT5), .B(G176gat), .ZN(new_n274_));
  XOR2_X1   g073(.A(new_n273_), .B(new_n274_), .Z(new_n275_));
  NAND2_X1  g074(.A1(new_n271_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(new_n275_), .ZN(new_n277_));
  NAND3_X1  g076(.A1(new_n259_), .A2(new_n270_), .A3(new_n277_), .ZN(new_n278_));
  NAND2_X1  g077(.A1(new_n276_), .A2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT13), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n276_), .A2(KEYINPUT13), .A3(new_n278_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n281_), .A2(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(KEYINPUT97), .ZN(new_n284_));
  NAND2_X1  g083(.A1(G141gat), .A2(G148gat), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT2), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT3), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n288_), .B1(G141gat), .B2(G148gat), .ZN(new_n289_));
  NOR2_X1   g088(.A1(G141gat), .A2(G148gat), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n290_), .A2(KEYINPUT3), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n287_), .B1(new_n289_), .B2(new_n291_), .ZN(new_n292_));
  NAND2_X1  g091(.A1(new_n285_), .A2(KEYINPUT81), .ZN(new_n293_));
  INV_X1    g092(.A(KEYINPUT81), .ZN(new_n294_));
  NAND3_X1  g093(.A1(new_n294_), .A2(G141gat), .A3(G148gat), .ZN(new_n295_));
  AND2_X1   g094(.A1(new_n286_), .A2(KEYINPUT84), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n286_), .A2(KEYINPUT84), .ZN(new_n297_));
  OAI211_X1 g096(.A(new_n293_), .B(new_n295_), .C1(new_n296_), .C2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n292_), .A2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(KEYINPUT85), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n299_), .A2(new_n300_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n292_), .A2(new_n298_), .A3(KEYINPUT85), .ZN(new_n302_));
  INV_X1    g101(.A(G155gat), .ZN(new_n303_));
  INV_X1    g102(.A(G162gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND2_X1  g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n307_), .B(KEYINPUT86), .ZN(new_n308_));
  NAND3_X1  g107(.A1(new_n301_), .A2(new_n302_), .A3(new_n308_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n293_), .A2(new_n295_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT1), .ZN(new_n311_));
  NAND3_X1  g110(.A1(new_n305_), .A2(new_n311_), .A3(new_n306_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  XOR2_X1   g113(.A(new_n290_), .B(KEYINPUT82), .Z(new_n315_));
  OAI21_X1  g114(.A(KEYINPUT83), .B1(new_n314_), .B2(new_n315_), .ZN(new_n316_));
  AND2_X1   g115(.A1(new_n312_), .A2(new_n313_), .ZN(new_n317_));
  INV_X1    g116(.A(KEYINPUT83), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n290_), .B(KEYINPUT82), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n317_), .A2(new_n318_), .A3(new_n310_), .A4(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n316_), .A2(new_n320_), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n309_), .A2(new_n321_), .A3(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n323_), .A2(G50gat), .ZN(new_n324_));
  INV_X1    g123(.A(G50gat), .ZN(new_n325_));
  NAND4_X1  g124(.A1(new_n309_), .A2(new_n321_), .A3(new_n322_), .A4(new_n325_), .ZN(new_n326_));
  NAND2_X1  g125(.A1(new_n324_), .A2(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT28), .B(G22gat), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NAND3_X1  g129(.A1(new_n324_), .A2(new_n328_), .A3(new_n326_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  XOR2_X1   g131(.A(G78gat), .B(G106gat), .Z(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G228gat), .A2(G233gat), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n309_), .A2(new_n321_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT29), .ZN(new_n337_));
  XNOR2_X1  g136(.A(G197gat), .B(G204gat), .ZN(new_n338_));
  INV_X1    g137(.A(KEYINPUT21), .ZN(new_n339_));
  NAND2_X1  g138(.A1(new_n338_), .A2(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(G197gat), .ZN(new_n341_));
  NOR2_X1   g140(.A1(new_n341_), .A2(G204gat), .ZN(new_n342_));
  INV_X1    g141(.A(G204gat), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n343_), .A2(G197gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT21), .B1(new_n342_), .B2(new_n344_), .ZN(new_n345_));
  XNOR2_X1  g144(.A(G211gat), .B(G218gat), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n340_), .A2(new_n345_), .A3(new_n346_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n347_), .A2(KEYINPUT87), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n345_), .A2(new_n346_), .ZN(new_n349_));
  INV_X1    g148(.A(KEYINPUT87), .ZN(new_n350_));
  NAND4_X1  g149(.A1(new_n340_), .A2(new_n345_), .A3(new_n350_), .A4(new_n346_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n348_), .A2(new_n349_), .A3(new_n351_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n335_), .B1(new_n337_), .B2(new_n352_), .ZN(new_n353_));
  AOI21_X1  g152(.A(new_n322_), .B1(new_n309_), .B2(new_n321_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n352_), .ZN(new_n355_));
  INV_X1    g154(.A(new_n335_), .ZN(new_n356_));
  NOR3_X1   g155(.A1(new_n354_), .A2(new_n355_), .A3(new_n356_), .ZN(new_n357_));
  OAI21_X1  g156(.A(new_n334_), .B1(new_n353_), .B2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT88), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n337_), .A2(new_n352_), .A3(new_n335_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n356_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n360_), .A2(new_n361_), .A3(new_n333_), .ZN(new_n362_));
  NAND4_X1  g161(.A1(new_n332_), .A2(new_n358_), .A3(new_n359_), .A4(new_n362_), .ZN(new_n363_));
  AND3_X1   g162(.A1(new_n324_), .A2(new_n328_), .A3(new_n326_), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n328_), .B1(new_n324_), .B2(new_n326_), .ZN(new_n365_));
  NOR2_X1   g164(.A1(new_n364_), .A2(new_n365_), .ZN(new_n366_));
  NOR3_X1   g165(.A1(new_n353_), .A2(new_n357_), .A3(new_n334_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n333_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n368_));
  OAI21_X1  g167(.A(new_n366_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n367_), .A2(KEYINPUT88), .ZN(new_n370_));
  NAND3_X1  g169(.A1(new_n363_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n371_));
  XNOR2_X1  g170(.A(G71gat), .B(G99gat), .ZN(new_n372_));
  NAND2_X1  g171(.A1(G227gat), .A2(G233gat), .ZN(new_n373_));
  XOR2_X1   g172(.A(new_n372_), .B(new_n373_), .Z(new_n374_));
  INV_X1    g173(.A(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(G183gat), .ZN(new_n376_));
  INV_X1    g175(.A(G190gat), .ZN(new_n377_));
  OAI21_X1  g176(.A(KEYINPUT23), .B1(new_n376_), .B2(new_n377_), .ZN(new_n378_));
  INV_X1    g177(.A(KEYINPUT23), .ZN(new_n379_));
  NAND3_X1  g178(.A1(new_n379_), .A2(G183gat), .A3(G190gat), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n378_), .A2(new_n380_), .ZN(new_n381_));
  OR3_X1    g180(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n382_));
  INV_X1    g181(.A(G169gat), .ZN(new_n383_));
  INV_X1    g182(.A(G176gat), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n383_), .A2(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(G169gat), .A2(G176gat), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(KEYINPUT24), .A3(new_n386_), .ZN(new_n387_));
  AND3_X1   g186(.A1(new_n381_), .A2(new_n382_), .A3(new_n387_), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT26), .B(G190gat), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n390_));
  OAI21_X1  g189(.A(new_n390_), .B1(new_n376_), .B2(KEYINPUT25), .ZN(new_n391_));
  XNOR2_X1  g190(.A(KEYINPUT25), .B(G183gat), .ZN(new_n392_));
  OAI211_X1 g191(.A(new_n389_), .B(new_n391_), .C1(new_n392_), .C2(new_n390_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n388_), .A2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n386_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n376_), .A2(new_n377_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n395_), .B1(new_n381_), .B2(new_n396_), .ZN(new_n397_));
  OR2_X1    g196(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n398_));
  NAND2_X1  g197(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n399_));
  AOI21_X1  g198(.A(G176gat), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  INV_X1    g199(.A(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n397_), .A2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n394_), .A2(new_n402_), .ZN(new_n403_));
  XNOR2_X1  g202(.A(new_n403_), .B(KEYINPUT30), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G127gat), .B(G134gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(G113gat), .B(G120gat), .ZN(new_n406_));
  XNOR2_X1  g205(.A(new_n405_), .B(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n404_), .A2(new_n408_), .ZN(new_n409_));
  AOI22_X1  g208(.A1(new_n388_), .A2(new_n393_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n410_), .B(KEYINPUT30), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n407_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(G15gat), .B(G43gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n413_), .B(KEYINPUT31), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n409_), .A2(new_n412_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n416_), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n415_), .B1(new_n409_), .B2(new_n412_), .ZN(new_n418_));
  OAI21_X1  g217(.A(new_n375_), .B1(new_n417_), .B2(new_n418_), .ZN(new_n419_));
  INV_X1    g218(.A(new_n418_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n420_), .A2(new_n374_), .A3(new_n416_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n419_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n371_), .A2(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT27), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n392_), .A2(new_n389_), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n388_), .A2(new_n425_), .ZN(new_n426_));
  AOI21_X1  g225(.A(KEYINPUT89), .B1(new_n397_), .B2(new_n401_), .ZN(new_n427_));
  AOI22_X1  g226(.A1(new_n378_), .A2(new_n380_), .B1(new_n376_), .B2(new_n377_), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT89), .ZN(new_n429_));
  NOR4_X1   g228(.A1(new_n428_), .A2(new_n400_), .A3(new_n429_), .A4(new_n395_), .ZN(new_n430_));
  OAI21_X1  g229(.A(new_n426_), .B1(new_n427_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n431_), .A2(new_n352_), .ZN(new_n432_));
  NAND4_X1  g231(.A1(new_n410_), .A2(new_n349_), .A3(new_n351_), .A4(new_n348_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n432_), .A2(KEYINPUT20), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(G226gat), .A2(G233gat), .ZN(new_n435_));
  XNOR2_X1  g234(.A(new_n435_), .B(KEYINPUT19), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n437_));
  AOI211_X1 g236(.A(new_n437_), .B(new_n436_), .C1(new_n352_), .C2(new_n403_), .ZN(new_n438_));
  OR2_X1    g237(.A1(new_n431_), .A2(new_n352_), .ZN(new_n439_));
  AOI22_X1  g238(.A1(new_n434_), .A2(new_n436_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n440_));
  XNOR2_X1  g239(.A(G8gat), .B(G36gat), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(G92gat), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT18), .B(G64gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n442_), .B(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  AOI21_X1  g244(.A(new_n424_), .B1(new_n440_), .B2(new_n445_), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT95), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n437_), .B1(new_n352_), .B2(new_n403_), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n388_), .A2(new_n425_), .B1(new_n397_), .B2(new_n401_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n449_), .A2(new_n349_), .A3(new_n351_), .A4(new_n348_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  AOI21_X1  g250(.A(new_n447_), .B1(new_n451_), .B2(new_n436_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n436_), .ZN(new_n453_));
  AOI211_X1 g252(.A(KEYINPUT95), .B(new_n453_), .C1(new_n448_), .C2(new_n450_), .ZN(new_n454_));
  AND4_X1   g253(.A1(KEYINPUT20), .A2(new_n432_), .A3(new_n453_), .A4(new_n433_), .ZN(new_n455_));
  NOR3_X1   g254(.A1(new_n452_), .A2(new_n454_), .A3(new_n455_), .ZN(new_n456_));
  OAI21_X1  g255(.A(new_n446_), .B1(new_n456_), .B2(new_n445_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n336_), .A2(new_n408_), .ZN(new_n458_));
  NAND3_X1  g257(.A1(new_n309_), .A2(new_n321_), .A3(new_n407_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(KEYINPUT4), .A3(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(G225gat), .A2(G233gat), .ZN(new_n461_));
  XNOR2_X1  g260(.A(new_n461_), .B(KEYINPUT90), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n462_), .B(KEYINPUT91), .Z(new_n463_));
  AOI21_X1  g262(.A(new_n407_), .B1(new_n309_), .B2(new_n321_), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT4), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n463_), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n460_), .A2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT92), .ZN(new_n468_));
  AND3_X1   g267(.A1(new_n309_), .A2(new_n321_), .A3(new_n407_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n469_), .A2(new_n464_), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n468_), .B1(new_n470_), .B2(new_n462_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n458_), .A2(new_n468_), .A3(new_n462_), .A4(new_n459_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n467_), .B1(new_n471_), .B2(new_n473_), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G1gat), .B(G29gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(new_n212_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(KEYINPUT0), .B(G57gat), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n476_), .B(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n474_), .A2(new_n479_), .ZN(new_n480_));
  NAND2_X1  g279(.A1(new_n434_), .A2(new_n436_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n438_), .A2(new_n439_), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n481_), .A2(new_n445_), .A3(new_n482_), .ZN(new_n483_));
  AOI21_X1  g282(.A(new_n445_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n424_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  OAI211_X1 g284(.A(new_n467_), .B(new_n478_), .C1(new_n471_), .C2(new_n473_), .ZN(new_n486_));
  NAND4_X1  g285(.A1(new_n457_), .A2(new_n480_), .A3(new_n485_), .A4(new_n486_), .ZN(new_n487_));
  NOR2_X1   g286(.A1(new_n423_), .A2(new_n487_), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n363_), .A2(new_n369_), .A3(new_n370_), .ZN(new_n489_));
  AOI21_X1  g288(.A(new_n422_), .B1(new_n487_), .B2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(KEYINPUT33), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n486_), .A2(new_n491_), .ZN(new_n492_));
  NOR3_X1   g291(.A1(new_n469_), .A2(new_n464_), .A3(new_n463_), .ZN(new_n493_));
  OR3_X1    g292(.A1(new_n493_), .A2(KEYINPUT93), .A3(new_n478_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n464_), .A2(new_n465_), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n460_), .A2(new_n462_), .A3(new_n495_), .ZN(new_n496_));
  INV_X1    g295(.A(KEYINPUT94), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  OAI21_X1  g297(.A(KEYINPUT93), .B1(new_n493_), .B2(new_n478_), .ZN(new_n499_));
  NAND4_X1  g298(.A1(new_n460_), .A2(KEYINPUT94), .A3(new_n462_), .A4(new_n495_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n494_), .A2(new_n498_), .A3(new_n499_), .A4(new_n500_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n458_), .A2(new_n462_), .A3(new_n459_), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n502_), .A2(KEYINPUT92), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(new_n472_), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n504_), .A2(KEYINPUT33), .A3(new_n467_), .A4(new_n478_), .ZN(new_n505_));
  NOR2_X1   g304(.A1(new_n483_), .A2(new_n484_), .ZN(new_n506_));
  NAND4_X1  g305(.A1(new_n492_), .A2(new_n501_), .A3(new_n505_), .A4(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n451_), .A2(new_n436_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT95), .ZN(new_n509_));
  NAND3_X1  g308(.A1(new_n451_), .A2(new_n447_), .A3(new_n436_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n509_), .A2(new_n510_), .ZN(new_n511_));
  OAI211_X1 g310(.A(KEYINPUT32), .B(new_n445_), .C1(new_n511_), .C2(new_n455_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT32), .ZN(new_n513_));
  OAI21_X1  g312(.A(new_n440_), .B1(new_n513_), .B2(new_n444_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n486_), .ZN(new_n515_));
  AOI21_X1  g314(.A(new_n478_), .B1(new_n504_), .B2(new_n467_), .ZN(new_n516_));
  OAI211_X1 g315(.A(new_n512_), .B(new_n514_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n517_));
  NAND3_X1  g316(.A1(new_n507_), .A2(new_n517_), .A3(new_n371_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n490_), .A2(new_n518_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n519_), .A2(KEYINPUT96), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT96), .ZN(new_n521_));
  NAND3_X1  g320(.A1(new_n490_), .A2(new_n518_), .A3(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n488_), .B1(new_n520_), .B2(new_n522_), .ZN(new_n523_));
  XNOR2_X1  g322(.A(G1gat), .B(G8gat), .ZN(new_n524_));
  XNOR2_X1  g323(.A(new_n524_), .B(KEYINPUT77), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526_));
  INV_X1    g325(.A(G1gat), .ZN(new_n527_));
  INV_X1    g326(.A(G8gat), .ZN(new_n528_));
  OAI21_X1  g327(.A(KEYINPUT14), .B1(new_n527_), .B2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n526_), .A2(new_n529_), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n525_), .B(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT79), .ZN(new_n532_));
  INV_X1    g331(.A(G29gat), .ZN(new_n533_));
  INV_X1    g332(.A(G36gat), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n533_), .A2(new_n534_), .ZN(new_n535_));
  NAND2_X1  g334(.A1(G29gat), .A2(G36gat), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n535_), .A2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(G43gat), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n538_), .A2(G50gat), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n325_), .A2(G43gat), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n537_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  XNOR2_X1  g340(.A(G43gat), .B(G50gat), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n542_), .A2(new_n535_), .A3(new_n536_), .ZN(new_n543_));
  AND3_X1   g342(.A1(new_n541_), .A2(new_n543_), .A3(KEYINPUT15), .ZN(new_n544_));
  AOI21_X1  g343(.A(KEYINPUT15), .B1(new_n541_), .B2(new_n543_), .ZN(new_n545_));
  OAI211_X1 g344(.A(new_n531_), .B(new_n532_), .C1(new_n544_), .C2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n530_), .ZN(new_n547_));
  XNOR2_X1  g346(.A(new_n525_), .B(new_n547_), .ZN(new_n548_));
  NOR2_X1   g347(.A1(new_n544_), .A2(new_n545_), .ZN(new_n549_));
  OAI21_X1  g348(.A(KEYINPUT79), .B1(new_n548_), .B2(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(G229gat), .A2(G233gat), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n541_), .A2(new_n543_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n552_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n548_), .A2(new_n553_), .ZN(new_n554_));
  NAND4_X1  g353(.A1(new_n546_), .A2(new_n550_), .A3(new_n551_), .A4(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(new_n551_), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n548_), .A2(new_n553_), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n531_), .A2(new_n552_), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n556_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  XNOR2_X1  g358(.A(G113gat), .B(G141gat), .ZN(new_n560_));
  XNOR2_X1  g359(.A(G169gat), .B(G197gat), .ZN(new_n561_));
  XNOR2_X1  g360(.A(new_n560_), .B(new_n561_), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  AND3_X1   g362(.A1(new_n555_), .A2(new_n559_), .A3(new_n563_), .ZN(new_n564_));
  AOI21_X1  g363(.A(new_n563_), .B1(new_n555_), .B2(new_n559_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n564_), .A2(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n284_), .B1(new_n523_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n488_), .ZN(new_n568_));
  AND3_X1   g367(.A1(new_n490_), .A2(new_n518_), .A3(new_n521_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n521_), .B1(new_n490_), .B2(new_n518_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n568_), .B1(new_n569_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n566_), .ZN(new_n572_));
  NAND3_X1  g371(.A1(new_n571_), .A2(KEYINPUT97), .A3(new_n572_), .ZN(new_n573_));
  AOI21_X1  g372(.A(new_n283_), .B1(new_n567_), .B2(new_n573_), .ZN(new_n574_));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575_));
  XNOR2_X1  g374(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n575_), .B(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(G127gat), .B(G155gat), .ZN(new_n578_));
  XOR2_X1   g377(.A(new_n577_), .B(new_n578_), .Z(new_n579_));
  XOR2_X1   g378(.A(new_n579_), .B(KEYINPUT17), .Z(new_n580_));
  INV_X1    g379(.A(new_n579_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n581_), .A2(KEYINPUT17), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n242_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n548_), .ZN(new_n585_));
  MUX2_X1   g384(.A(new_n580_), .B(new_n582_), .S(new_n585_), .Z(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT71), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n549_), .A2(new_n228_), .ZN(new_n589_));
  NAND4_X1  g388(.A1(new_n219_), .A2(new_n552_), .A3(new_n226_), .A4(new_n227_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n589_), .A2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(KEYINPUT69), .B(KEYINPUT34), .ZN(new_n592_));
  AND2_X1   g391(.A1(G232gat), .A2(G233gat), .ZN(new_n593_));
  OR2_X1    g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n592_), .A2(new_n593_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT35), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT35), .ZN(new_n598_));
  NAND3_X1  g397(.A1(new_n594_), .A2(new_n598_), .A3(new_n595_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n597_), .A2(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AOI21_X1  g400(.A(new_n588_), .B1(new_n591_), .B2(new_n601_), .ZN(new_n602_));
  AOI211_X1 g401(.A(KEYINPUT71), .B(new_n600_), .C1(new_n589_), .C2(new_n590_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n591_), .A2(new_n597_), .ZN(new_n604_));
  NOR3_X1   g403(.A1(new_n602_), .A2(new_n603_), .A3(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(G218gat), .ZN(new_n607_));
  XNOR2_X1  g406(.A(KEYINPUT70), .B(G190gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n607_), .B(new_n608_), .Z(new_n609_));
  INV_X1    g408(.A(KEYINPUT36), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n607_), .B(new_n608_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n612_), .A2(KEYINPUT36), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n611_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n614_), .A2(KEYINPUT73), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT73), .ZN(new_n616_));
  NAND3_X1  g415(.A1(new_n611_), .A2(new_n613_), .A3(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n615_), .A2(new_n617_), .ZN(new_n618_));
  OAI21_X1  g417(.A(KEYINPUT74), .B1(new_n605_), .B2(new_n618_), .ZN(new_n619_));
  INV_X1    g418(.A(new_n617_), .ZN(new_n620_));
  AOI21_X1  g419(.A(new_n616_), .B1(new_n611_), .B2(new_n613_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n620_), .A2(new_n621_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n591_), .A2(new_n601_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n623_), .A2(KEYINPUT71), .ZN(new_n624_));
  INV_X1    g423(.A(new_n604_), .ZN(new_n625_));
  NAND3_X1  g424(.A1(new_n591_), .A2(new_n588_), .A3(new_n601_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n624_), .A2(new_n625_), .A3(new_n626_), .ZN(new_n627_));
  INV_X1    g426(.A(KEYINPUT74), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n622_), .A2(new_n627_), .A3(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n611_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n605_), .A2(KEYINPUT72), .A3(new_n630_), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n624_), .A2(new_n625_), .A3(new_n630_), .A4(new_n626_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT72), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n632_), .A2(new_n633_), .ZN(new_n634_));
  NAND4_X1  g433(.A1(new_n619_), .A2(new_n629_), .A3(new_n631_), .A4(new_n634_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n635_), .A2(KEYINPUT37), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT75), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n605_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n627_), .A2(KEYINPUT75), .ZN(new_n639_));
  NAND4_X1  g438(.A1(new_n638_), .A2(new_n639_), .A3(new_n611_), .A4(new_n613_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT37), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n641_), .A3(new_n632_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n636_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n643_), .A2(KEYINPUT76), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT76), .ZN(new_n645_));
  NAND3_X1  g444(.A1(new_n636_), .A2(new_n642_), .A3(new_n645_), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n587_), .B1(new_n644_), .B2(new_n646_), .ZN(new_n647_));
  AND2_X1   g446(.A1(new_n574_), .A2(new_n647_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n515_), .A2(new_n516_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n648_), .A2(new_n527_), .A3(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(KEYINPUT38), .ZN(new_n652_));
  OR2_X1    g451(.A1(new_n651_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n640_), .A2(new_n632_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n587_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n283_), .A2(new_n566_), .ZN(new_n657_));
  NAND3_X1  g456(.A1(new_n571_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n658_));
  OAI21_X1  g457(.A(G1gat), .B1(new_n658_), .B2(new_n649_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n651_), .A2(new_n652_), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n653_), .A2(new_n659_), .A3(new_n660_), .ZN(G1324gat));
  INV_X1    g460(.A(KEYINPUT39), .ZN(new_n662_));
  AND3_X1   g461(.A1(new_n571_), .A2(new_n656_), .A3(new_n657_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n457_), .A2(new_n485_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  AOI21_X1  g464(.A(new_n528_), .B1(new_n663_), .B2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n662_), .B1(new_n666_), .B2(KEYINPUT98), .ZN(new_n667_));
  OAI21_X1  g466(.A(new_n667_), .B1(KEYINPUT98), .B2(new_n666_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n648_), .A2(new_n528_), .A3(new_n665_), .ZN(new_n669_));
  OR3_X1    g468(.A1(new_n666_), .A2(KEYINPUT98), .A3(KEYINPUT39), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n668_), .A2(new_n669_), .A3(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT40), .ZN(new_n672_));
  XNOR2_X1  g471(.A(new_n671_), .B(new_n672_), .ZN(G1325gat));
  INV_X1    g472(.A(new_n422_), .ZN(new_n674_));
  OAI21_X1  g473(.A(G15gat), .B1(new_n658_), .B2(new_n674_), .ZN(new_n675_));
  XOR2_X1   g474(.A(KEYINPUT99), .B(KEYINPUT41), .Z(new_n676_));
  XNOR2_X1  g475(.A(new_n675_), .B(new_n676_), .ZN(new_n677_));
  INV_X1    g476(.A(new_n648_), .ZN(new_n678_));
  OR2_X1    g477(.A1(new_n674_), .A2(G15gat), .ZN(new_n679_));
  OAI21_X1  g478(.A(new_n677_), .B1(new_n678_), .B2(new_n679_), .ZN(G1326gat));
  OAI21_X1  g479(.A(G22gat), .B1(new_n658_), .B2(new_n371_), .ZN(new_n681_));
  XNOR2_X1  g480(.A(new_n681_), .B(KEYINPUT100), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n682_), .B(KEYINPUT42), .ZN(new_n683_));
  OR2_X1    g482(.A1(new_n678_), .A2(G22gat), .ZN(new_n684_));
  OAI21_X1  g483(.A(new_n683_), .B1(new_n371_), .B2(new_n684_), .ZN(G1327gat));
  NAND2_X1  g484(.A1(new_n657_), .A2(new_n587_), .ZN(new_n686_));
  AND3_X1   g485(.A1(new_n636_), .A2(new_n642_), .A3(new_n645_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n645_), .B1(new_n636_), .B2(new_n642_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  INV_X1    g488(.A(new_n689_), .ZN(new_n690_));
  OAI21_X1  g489(.A(KEYINPUT43), .B1(new_n523_), .B2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT43), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n571_), .A2(new_n692_), .A3(new_n689_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n686_), .B1(new_n691_), .B2(new_n693_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(KEYINPUT44), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n650_), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n694_), .A2(KEYINPUT44), .ZN(new_n697_));
  OAI21_X1  g496(.A(G29gat), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n654_), .A2(new_n586_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n574_), .A2(new_n699_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n650_), .A2(new_n533_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT101), .ZN(new_n702_));
  OAI21_X1  g501(.A(new_n698_), .B1(new_n700_), .B2(new_n702_), .ZN(G1328gat));
  INV_X1    g502(.A(new_n697_), .ZN(new_n704_));
  AOI21_X1  g503(.A(new_n664_), .B1(new_n694_), .B2(KEYINPUT44), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n706_), .A2(G36gat), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n708_));
  NOR2_X1   g507(.A1(new_n664_), .A2(G36gat), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n708_), .B1(new_n700_), .B2(new_n710_), .ZN(new_n711_));
  NAND4_X1  g510(.A1(new_n574_), .A2(KEYINPUT45), .A3(new_n699_), .A4(new_n709_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(KEYINPUT102), .B(KEYINPUT46), .ZN(new_n713_));
  NAND4_X1  g512(.A1(new_n707_), .A2(new_n711_), .A3(new_n712_), .A4(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(new_n713_), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n711_), .A2(new_n712_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n534_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n715_), .B1(new_n716_), .B2(new_n717_), .ZN(new_n718_));
  AND2_X1   g517(.A1(new_n714_), .A2(new_n718_), .ZN(G1329gat));
  OAI21_X1  g518(.A(new_n538_), .B1(new_n700_), .B2(new_n674_), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n704_), .A2(G43gat), .A3(new_n422_), .ZN(new_n721_));
  INV_X1    g520(.A(new_n695_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n720_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT47), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n725_), .B(new_n720_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1330gat));
  NAND4_X1  g526(.A1(new_n704_), .A2(G50gat), .A3(new_n489_), .A4(new_n695_), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n325_), .B1(new_n700_), .B2(new_n371_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT103), .ZN(G1331gat));
  NAND4_X1  g530(.A1(new_n571_), .A2(new_n656_), .A3(new_n566_), .A4(new_n283_), .ZN(new_n732_));
  NOR3_X1   g531(.A1(new_n732_), .A2(new_n233_), .A3(new_n649_), .ZN(new_n733_));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n734_), .B1(new_n523_), .B2(new_n572_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n571_), .A2(KEYINPUT104), .A3(new_n566_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n735_), .A2(new_n283_), .A3(new_n736_), .ZN(new_n737_));
  INV_X1    g536(.A(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n647_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT105), .B1(new_n738_), .B2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT105), .ZN(new_n741_));
  NAND3_X1  g540(.A1(new_n737_), .A2(new_n741_), .A3(new_n647_), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n740_), .A2(new_n650_), .A3(new_n742_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n733_), .B1(new_n743_), .B2(new_n233_), .ZN(G1332gat));
  OAI21_X1  g543(.A(G64gat), .B1(new_n732_), .B2(new_n664_), .ZN(new_n745_));
  XOR2_X1   g544(.A(KEYINPUT106), .B(KEYINPUT48), .Z(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n740_), .A2(new_n742_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n665_), .A2(new_n234_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n747_), .B1(new_n748_), .B2(new_n749_), .ZN(G1333gat));
  OAI21_X1  g549(.A(G71gat), .B1(new_n732_), .B2(new_n674_), .ZN(new_n751_));
  XNOR2_X1  g550(.A(new_n751_), .B(KEYINPUT49), .ZN(new_n752_));
  OR2_X1    g551(.A1(new_n674_), .A2(G71gat), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n752_), .B1(new_n748_), .B2(new_n753_), .ZN(G1334gat));
  OAI21_X1  g553(.A(G78gat), .B1(new_n732_), .B2(new_n371_), .ZN(new_n755_));
  XNOR2_X1  g554(.A(new_n755_), .B(KEYINPUT50), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n371_), .A2(G78gat), .ZN(new_n757_));
  OAI21_X1  g556(.A(new_n756_), .B1(new_n748_), .B2(new_n757_), .ZN(G1335gat));
  AND4_X1   g557(.A1(new_n283_), .A2(new_n735_), .A3(new_n699_), .A4(new_n736_), .ZN(new_n759_));
  AOI21_X1  g558(.A(G85gat), .B1(new_n759_), .B2(new_n650_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n691_), .A2(new_n693_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n572_), .B1(new_n281_), .B2(new_n282_), .ZN(new_n762_));
  AND3_X1   g561(.A1(new_n762_), .A2(KEYINPUT107), .A3(new_n587_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT107), .B1(new_n762_), .B2(new_n587_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n763_), .A2(new_n764_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n761_), .A2(new_n766_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n767_), .A2(new_n212_), .A3(new_n649_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n760_), .A2(new_n768_), .ZN(G1336gat));
  AOI21_X1  g568(.A(G92gat), .B1(new_n759_), .B2(new_n665_), .ZN(new_n770_));
  NOR3_X1   g569(.A1(new_n767_), .A2(new_n213_), .A3(new_n664_), .ZN(new_n771_));
  NOR2_X1   g570(.A1(new_n770_), .A2(new_n771_), .ZN(G1337gat));
  OAI21_X1  g571(.A(G99gat), .B1(new_n767_), .B2(new_n674_), .ZN(new_n773_));
  INV_X1    g572(.A(new_n759_), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n422_), .B1(new_n220_), .B2(new_n221_), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n773_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  XNOR2_X1  g575(.A(new_n776_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND4_X1  g576(.A1(new_n737_), .A2(new_n204_), .A3(new_n489_), .A4(new_n699_), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n759_), .A2(KEYINPUT108), .A3(new_n204_), .A4(new_n489_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n780_), .A2(new_n781_), .ZN(new_n782_));
  AOI211_X1 g581(.A(new_n371_), .B(new_n765_), .C1(new_n691_), .C2(new_n693_), .ZN(new_n783_));
  OAI21_X1  g582(.A(KEYINPUT109), .B1(new_n783_), .B2(new_n204_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n761_), .A2(new_n489_), .A3(new_n766_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n786_));
  NAND3_X1  g585(.A1(new_n785_), .A2(new_n786_), .A3(G106gat), .ZN(new_n787_));
  NAND3_X1  g586(.A1(new_n784_), .A2(KEYINPUT52), .A3(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789_));
  OAI211_X1 g588(.A(KEYINPUT109), .B(new_n789_), .C1(new_n783_), .C2(new_n204_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n782_), .A2(new_n788_), .A3(new_n790_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n791_), .A2(KEYINPUT53), .ZN(new_n792_));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793_));
  NAND4_X1  g592(.A1(new_n782_), .A2(new_n788_), .A3(new_n793_), .A4(new_n790_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(G1339gat));
  INV_X1    g594(.A(new_n423_), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n665_), .A2(new_n649_), .ZN(new_n797_));
  INV_X1    g596(.A(KEYINPUT57), .ZN(new_n798_));
  NAND4_X1  g597(.A1(new_n546_), .A2(new_n550_), .A3(new_n556_), .A4(new_n554_), .ZN(new_n799_));
  OAI21_X1  g598(.A(new_n551_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n800_));
  AND3_X1   g599(.A1(new_n799_), .A2(new_n562_), .A3(new_n800_), .ZN(new_n801_));
  NOR2_X1   g600(.A1(new_n564_), .A2(new_n801_), .ZN(new_n802_));
  AND3_X1   g601(.A1(new_n259_), .A2(new_n270_), .A3(new_n277_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n277_), .B1(new_n259_), .B2(new_n270_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n802_), .B1(new_n803_), .B2(new_n804_), .ZN(new_n805_));
  NAND2_X1  g604(.A1(new_n805_), .A2(KEYINPUT111), .ZN(new_n806_));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n279_), .A2(new_n807_), .A3(new_n802_), .ZN(new_n808_));
  AND2_X1   g607(.A1(new_n806_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT55), .B1(new_n252_), .B2(new_n258_), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n255_), .A2(new_n256_), .ZN(new_n811_));
  XNOR2_X1  g610(.A(new_n249_), .B(new_n264_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n260_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT55), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n813_), .B1(new_n814_), .B2(new_n257_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n275_), .B1(new_n810_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(KEYINPUT56), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT110), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT56), .B(new_n275_), .C1(new_n810_), .C2(new_n815_), .ZN(new_n820_));
  NAND3_X1  g619(.A1(new_n818_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n816_), .A2(KEYINPUT110), .A3(new_n817_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n803_), .A2(new_n566_), .ZN(new_n823_));
  NAND3_X1  g622(.A1(new_n821_), .A2(new_n822_), .A3(new_n823_), .ZN(new_n824_));
  AOI211_X1 g623(.A(new_n798_), .B(new_n655_), .C1(new_n809_), .C2(new_n824_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n818_), .A2(new_n819_), .A3(new_n820_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n822_), .A2(new_n823_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n806_), .B(new_n808_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n828_));
  AOI21_X1  g627(.A(KEYINPUT57), .B1(new_n828_), .B2(new_n654_), .ZN(new_n829_));
  NOR2_X1   g628(.A1(new_n825_), .A2(new_n829_), .ZN(new_n830_));
  INV_X1    g629(.A(new_n820_), .ZN(new_n831_));
  INV_X1    g630(.A(KEYINPUT112), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n803_), .B1(new_n831_), .B2(new_n832_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n818_), .A2(KEYINPUT112), .A3(new_n820_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n833_), .A2(new_n802_), .A3(new_n834_), .ZN(new_n835_));
  INV_X1    g634(.A(KEYINPUT58), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n835_), .A2(new_n836_), .ZN(new_n837_));
  NAND4_X1  g636(.A1(new_n833_), .A2(new_n834_), .A3(KEYINPUT58), .A4(new_n802_), .ZN(new_n838_));
  NAND3_X1  g637(.A1(new_n689_), .A2(new_n837_), .A3(new_n838_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n586_), .B1(new_n830_), .B2(new_n839_), .ZN(new_n840_));
  OAI211_X1 g639(.A(new_n586_), .B(new_n566_), .C1(new_n687_), .C2(new_n688_), .ZN(new_n841_));
  OAI21_X1  g640(.A(KEYINPUT54), .B1(new_n841_), .B2(new_n283_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843_));
  INV_X1    g642(.A(new_n283_), .ZN(new_n844_));
  NAND4_X1  g643(.A1(new_n647_), .A2(new_n843_), .A3(new_n566_), .A4(new_n844_), .ZN(new_n845_));
  AND2_X1   g644(.A1(new_n842_), .A2(new_n845_), .ZN(new_n846_));
  OAI211_X1 g645(.A(new_n796_), .B(new_n797_), .C1(new_n840_), .C2(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(G113gat), .B1(new_n848_), .B2(new_n572_), .ZN(new_n849_));
  OAI21_X1  g648(.A(KEYINPUT59), .B1(new_n847_), .B2(KEYINPUT113), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n828_), .A2(new_n654_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n851_), .A2(new_n798_), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n828_), .A2(KEYINPUT57), .A3(new_n654_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n852_), .A2(new_n839_), .A3(new_n853_), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n854_), .A2(new_n587_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n842_), .A2(new_n845_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n423_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  INV_X1    g656(.A(KEYINPUT113), .ZN(new_n858_));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859_));
  NAND4_X1  g658(.A1(new_n857_), .A2(new_n858_), .A3(new_n859_), .A4(new_n797_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n850_), .A2(KEYINPUT114), .A3(new_n860_), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT114), .B1(new_n850_), .B2(new_n860_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n862_), .ZN(new_n863_));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n572_), .A2(new_n864_), .A3(G113gat), .ZN(new_n865_));
  OAI21_X1  g664(.A(new_n865_), .B1(new_n864_), .B2(G113gat), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n849_), .B1(new_n863_), .B2(new_n866_), .ZN(G1340gat));
  NOR2_X1   g666(.A1(new_n844_), .A2(G120gat), .ZN(new_n868_));
  OAI211_X1 g667(.A(new_n857_), .B(new_n797_), .C1(KEYINPUT60), .C2(new_n868_), .ZN(new_n869_));
  NAND4_X1  g668(.A1(new_n850_), .A2(new_n869_), .A3(new_n283_), .A4(new_n860_), .ZN(new_n870_));
  NAND2_X1  g669(.A1(new_n870_), .A2(G120gat), .ZN(new_n871_));
  OAI21_X1  g670(.A(new_n871_), .B1(KEYINPUT60), .B2(new_n869_), .ZN(G1341gat));
  AOI21_X1  g671(.A(G127gat), .B1(new_n848_), .B2(new_n586_), .ZN(new_n873_));
  AND2_X1   g672(.A1(new_n586_), .A2(G127gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n873_), .B1(new_n863_), .B2(new_n874_), .ZN(G1342gat));
  AOI21_X1  g674(.A(G134gat), .B1(new_n848_), .B2(new_n655_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(KEYINPUT116), .B(G134gat), .ZN(new_n877_));
  NOR2_X1   g676(.A1(new_n690_), .A2(new_n877_), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n876_), .B1(new_n863_), .B2(new_n878_), .ZN(G1343gat));
  AOI22_X1  g678(.A1(new_n854_), .A2(new_n587_), .B1(new_n842_), .B2(new_n845_), .ZN(new_n880_));
  INV_X1    g679(.A(new_n880_), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n371_), .A2(new_n422_), .ZN(new_n882_));
  NAND3_X1  g681(.A1(new_n881_), .A2(new_n797_), .A3(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n572_), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n885_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g685(.A1(new_n884_), .A2(new_n283_), .ZN(new_n887_));
  XNOR2_X1  g686(.A(new_n887_), .B(G148gat), .ZN(G1345gat));
  OAI21_X1  g687(.A(G155gat), .B1(new_n883_), .B2(new_n587_), .ZN(new_n889_));
  NOR3_X1   g688(.A1(new_n880_), .A2(new_n371_), .A3(new_n422_), .ZN(new_n890_));
  NAND4_X1  g689(.A1(new_n890_), .A2(new_n303_), .A3(new_n586_), .A4(new_n797_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n889_), .A2(new_n891_), .ZN(new_n892_));
  XNOR2_X1  g691(.A(KEYINPUT117), .B(KEYINPUT61), .ZN(new_n893_));
  XNOR2_X1  g692(.A(new_n892_), .B(new_n893_), .ZN(G1346gat));
  NOR3_X1   g693(.A1(new_n883_), .A2(new_n304_), .A3(new_n690_), .ZN(new_n895_));
  NAND2_X1  g694(.A1(new_n884_), .A2(new_n655_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n895_), .B1(new_n896_), .B2(new_n304_), .ZN(G1347gat));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n898_));
  NOR2_X1   g697(.A1(new_n650_), .A2(new_n664_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n899_), .A2(new_n422_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n880_), .A2(new_n489_), .A3(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n901_), .A2(new_n572_), .ZN(new_n902_));
  AOI21_X1  g701(.A(new_n898_), .B1(new_n902_), .B2(G169gat), .ZN(new_n903_));
  AOI211_X1 g702(.A(KEYINPUT62), .B(new_n383_), .C1(new_n901_), .C2(new_n572_), .ZN(new_n904_));
  INV_X1    g703(.A(new_n901_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n566_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n906_));
  XOR2_X1   g705(.A(new_n906_), .B(KEYINPUT118), .Z(new_n907_));
  OAI22_X1  g706(.A1(new_n903_), .A2(new_n904_), .B1(new_n905_), .B2(new_n907_), .ZN(G1348gat));
  AOI21_X1  g707(.A(G176gat), .B1(new_n901_), .B2(new_n283_), .ZN(new_n909_));
  OAI21_X1  g708(.A(KEYINPUT119), .B1(new_n880_), .B2(new_n489_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n900_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT119), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n912_), .B(new_n371_), .C1(new_n840_), .C2(new_n846_), .ZN(new_n913_));
  AND3_X1   g712(.A1(new_n910_), .A2(new_n911_), .A3(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(new_n844_), .A2(new_n384_), .ZN(new_n915_));
  AOI21_X1  g714(.A(new_n909_), .B1(new_n914_), .B2(new_n915_), .ZN(G1349gat));
  NOR3_X1   g715(.A1(new_n905_), .A2(new_n587_), .A3(new_n392_), .ZN(new_n917_));
  NAND4_X1  g716(.A1(new_n910_), .A2(new_n913_), .A3(new_n586_), .A4(new_n911_), .ZN(new_n918_));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n919_));
  XNOR2_X1  g718(.A(new_n918_), .B(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(new_n917_), .B1(new_n920_), .B2(new_n376_), .ZN(G1350gat));
  NOR2_X1   g720(.A1(new_n905_), .A2(new_n690_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n655_), .A2(new_n389_), .ZN(new_n923_));
  XOR2_X1   g722(.A(new_n923_), .B(KEYINPUT121), .Z(new_n924_));
  OAI22_X1  g723(.A1(new_n922_), .A2(new_n377_), .B1(new_n905_), .B2(new_n924_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n925_), .A2(KEYINPUT122), .ZN(new_n926_));
  INV_X1    g725(.A(KEYINPUT122), .ZN(new_n927_));
  OAI221_X1 g726(.A(new_n927_), .B1(new_n905_), .B2(new_n924_), .C1(new_n922_), .C2(new_n377_), .ZN(new_n928_));
  NAND2_X1  g727(.A1(new_n926_), .A2(new_n928_), .ZN(G1351gat));
  NAND3_X1  g728(.A1(new_n890_), .A2(new_n572_), .A3(new_n899_), .ZN(new_n930_));
  AND3_X1   g729(.A1(new_n930_), .A2(KEYINPUT123), .A3(new_n341_), .ZN(new_n931_));
  AOI21_X1  g730(.A(KEYINPUT123), .B1(new_n930_), .B2(new_n341_), .ZN(new_n932_));
  NOR2_X1   g731(.A1(new_n930_), .A2(new_n341_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n931_), .A2(new_n932_), .A3(new_n933_), .ZN(G1352gat));
  NAND2_X1  g733(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n935_));
  NAND4_X1  g734(.A1(new_n890_), .A2(new_n283_), .A3(new_n899_), .A4(new_n935_), .ZN(new_n936_));
  NOR2_X1   g735(.A1(KEYINPUT124), .A2(G204gat), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(KEYINPUT125), .ZN(new_n938_));
  XNOR2_X1  g737(.A(new_n936_), .B(new_n938_), .ZN(G1353gat));
  NAND3_X1  g738(.A1(new_n881_), .A2(new_n882_), .A3(new_n899_), .ZN(new_n940_));
  NOR2_X1   g739(.A1(new_n940_), .A2(new_n587_), .ZN(new_n941_));
  OR2_X1    g740(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n941_), .A2(new_n942_), .ZN(new_n943_));
  XOR2_X1   g742(.A(KEYINPUT63), .B(G211gat), .Z(new_n944_));
  AOI21_X1  g743(.A(new_n943_), .B1(new_n941_), .B2(new_n944_), .ZN(G1354gat));
  XNOR2_X1  g744(.A(KEYINPUT126), .B(G218gat), .ZN(new_n946_));
  OR3_X1    g745(.A1(new_n940_), .A2(new_n654_), .A3(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948_));
  OAI21_X1  g747(.A(new_n946_), .B1(new_n940_), .B2(new_n690_), .ZN(new_n949_));
  AND3_X1   g748(.A1(new_n947_), .A2(new_n948_), .A3(new_n949_), .ZN(new_n950_));
  AOI21_X1  g749(.A(new_n948_), .B1(new_n947_), .B2(new_n949_), .ZN(new_n951_));
  NOR2_X1   g750(.A1(new_n950_), .A2(new_n951_), .ZN(G1355gat));
endmodule


