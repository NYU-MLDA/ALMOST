//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 0 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n643_, new_n644_, new_n645_, new_n647_, new_n648_,
    new_n649_, new_n650_, new_n651_, new_n652_, new_n653_, new_n654_,
    new_n655_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n864_, new_n865_, new_n866_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n877_, new_n878_, new_n879_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n918_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n929_, new_n930_, new_n931_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n941_, new_n942_, new_n943_;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT95), .B(G85gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  XNOR2_X1  g003(.A(KEYINPUT0), .B(G57gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT86), .ZN(new_n209_));
  AND2_X1   g008(.A1(new_n209_), .A2(KEYINPUT3), .ZN(new_n210_));
  NOR2_X1   g009(.A1(new_n209_), .A2(KEYINPUT3), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n208_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  AND2_X1   g011(.A1(G141gat), .A2(G148gat), .ZN(new_n213_));
  INV_X1    g012(.A(KEYINPUT2), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n214_), .A2(KEYINPUT87), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n209_), .A2(KEYINPUT3), .ZN(new_n216_));
  AOI22_X1  g015(.A1(new_n213_), .A2(new_n215_), .B1(new_n216_), .B2(new_n207_), .ZN(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT87), .B(KEYINPUT2), .ZN(new_n218_));
  OAI211_X1 g017(.A(new_n212_), .B(new_n217_), .C1(new_n213_), .C2(new_n218_), .ZN(new_n219_));
  XOR2_X1   g018(.A(G155gat), .B(G162gat), .Z(new_n220_));
  NAND2_X1  g019(.A1(new_n219_), .A2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n213_), .A2(new_n207_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223_));
  NAND2_X1  g022(.A1(new_n223_), .A2(KEYINPUT1), .ZN(new_n224_));
  OAI21_X1  g023(.A(new_n224_), .B1(G155gat), .B2(G162gat), .ZN(new_n225_));
  NOR2_X1   g024(.A1(new_n223_), .A2(KEYINPUT1), .ZN(new_n226_));
  OAI21_X1  g025(.A(new_n222_), .B1(new_n225_), .B2(new_n226_), .ZN(new_n227_));
  AND2_X1   g026(.A1(new_n221_), .A2(new_n227_), .ZN(new_n228_));
  INV_X1    g027(.A(KEYINPUT88), .ZN(new_n229_));
  NAND2_X1  g028(.A1(new_n228_), .A2(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n221_), .A2(new_n227_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT88), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  XNOR2_X1  g032(.A(G127gat), .B(G134gat), .ZN(new_n234_));
  XNOR2_X1  g033(.A(G113gat), .B(G120gat), .ZN(new_n235_));
  XNOR2_X1  g034(.A(new_n234_), .B(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n233_), .A2(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n228_), .A2(new_n236_), .ZN(new_n239_));
  AND2_X1   g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(G225gat), .A2(G233gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n240_), .A2(new_n241_), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT96), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n238_), .A2(new_n245_), .ZN(new_n246_));
  OAI21_X1  g045(.A(new_n246_), .B1(new_n240_), .B2(new_n245_), .ZN(new_n247_));
  XOR2_X1   g046(.A(new_n241_), .B(KEYINPUT94), .Z(new_n248_));
  NAND2_X1  g047(.A1(new_n247_), .A2(new_n248_), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n206_), .B1(new_n244_), .B2(new_n250_), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n242_), .B(KEYINPUT96), .ZN(new_n252_));
  INV_X1    g051(.A(new_n206_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(new_n249_), .ZN(new_n254_));
  AOI21_X1  g053(.A(KEYINPUT101), .B1(new_n251_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n251_), .A2(KEYINPUT101), .A3(new_n254_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n256_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G169gat), .A2(G176gat), .ZN(new_n260_));
  INV_X1    g059(.A(new_n260_), .ZN(new_n261_));
  XNOR2_X1  g060(.A(KEYINPUT22), .B(G169gat), .ZN(new_n262_));
  INV_X1    g061(.A(G176gat), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n261_), .B1(new_n262_), .B2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265_));
  XOR2_X1   g064(.A(new_n265_), .B(KEYINPUT23), .Z(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT83), .B(G190gat), .ZN(new_n267_));
  NOR2_X1   g066(.A1(new_n267_), .A2(G183gat), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n264_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  INV_X1    g068(.A(G169gat), .ZN(new_n270_));
  NAND2_X1  g069(.A1(new_n270_), .A2(new_n263_), .ZN(new_n271_));
  NOR2_X1   g070(.A1(new_n271_), .A2(KEYINPUT24), .ZN(new_n272_));
  NAND3_X1  g071(.A1(new_n271_), .A2(KEYINPUT24), .A3(new_n260_), .ZN(new_n273_));
  AOI211_X1 g072(.A(new_n272_), .B(new_n266_), .C1(KEYINPUT84), .C2(new_n273_), .ZN(new_n274_));
  OAI21_X1  g073(.A(new_n274_), .B1(KEYINPUT84), .B2(new_n273_), .ZN(new_n275_));
  XOR2_X1   g074(.A(KEYINPUT25), .B(G183gat), .Z(new_n276_));
  NAND2_X1  g075(.A1(new_n267_), .A2(KEYINPUT26), .ZN(new_n277_));
  OR2_X1    g076(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n276_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n269_), .B1(new_n275_), .B2(new_n279_), .ZN(new_n280_));
  XNOR2_X1  g079(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n281_));
  XNOR2_X1  g080(.A(new_n280_), .B(new_n281_), .ZN(new_n282_));
  XOR2_X1   g081(.A(G71gat), .B(G99gat), .Z(new_n283_));
  XNOR2_X1  g082(.A(KEYINPUT30), .B(G15gat), .ZN(new_n284_));
  XNOR2_X1  g083(.A(new_n283_), .B(new_n284_), .ZN(new_n285_));
  XNOR2_X1  g084(.A(new_n282_), .B(new_n285_), .ZN(new_n286_));
  NAND2_X1  g085(.A1(G227gat), .A2(G233gat), .ZN(new_n287_));
  INV_X1    g086(.A(G43gat), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n287_), .B(new_n288_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(new_n236_), .B(new_n289_), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n286_), .B(new_n290_), .ZN(new_n291_));
  INV_X1    g090(.A(new_n291_), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n233_), .A2(KEYINPUT29), .ZN(new_n293_));
  XNOR2_X1  g092(.A(KEYINPUT89), .B(KEYINPUT28), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G22gat), .B(G50gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT21), .ZN(new_n299_));
  XOR2_X1   g098(.A(G211gat), .B(G218gat), .Z(new_n300_));
  INV_X1    g099(.A(KEYINPUT90), .ZN(new_n301_));
  INV_X1    g100(.A(G197gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n302_), .A2(G204gat), .ZN(new_n303_));
  AOI211_X1 g102(.A(new_n299_), .B(new_n300_), .C1(new_n301_), .C2(new_n303_), .ZN(new_n304_));
  INV_X1    g103(.A(G204gat), .ZN(new_n305_));
  NAND2_X1  g104(.A1(new_n305_), .A2(G197gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n303_), .ZN(new_n307_));
  AND2_X1   g106(.A1(new_n304_), .A2(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n304_), .A2(new_n307_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n300_), .A2(new_n299_), .ZN(new_n310_));
  NOR3_X1   g109(.A1(new_n308_), .A2(new_n309_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n312_));
  OAI21_X1  g111(.A(new_n311_), .B1(new_n312_), .B2(new_n228_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(G228gat), .A3(G233gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n312_), .B1(new_n230_), .B2(new_n232_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(G228gat), .A2(G233gat), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n311_), .A2(new_n316_), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n314_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  XOR2_X1   g117(.A(G78gat), .B(G106gat), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n318_), .B(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(new_n319_), .ZN(new_n321_));
  NAND2_X1  g120(.A1(new_n318_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(KEYINPUT91), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n298_), .A2(new_n320_), .A3(new_n323_), .ZN(new_n324_));
  INV_X1    g123(.A(new_n320_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n323_), .ZN(new_n326_));
  OAI21_X1  g125(.A(new_n325_), .B1(new_n297_), .B2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n324_), .A2(new_n327_), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n266_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(new_n331_), .B(KEYINPUT92), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n332_), .A2(new_n264_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n266_), .A2(new_n272_), .ZN(new_n334_));
  XOR2_X1   g133(.A(KEYINPUT26), .B(G190gat), .Z(new_n335_));
  OAI211_X1 g134(.A(new_n334_), .B(new_n273_), .C1(new_n276_), .C2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n333_), .A2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n311_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n338_), .B(KEYINPUT20), .C1(new_n311_), .C2(new_n280_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(KEYINPUT19), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n339_), .A2(new_n341_), .ZN(new_n342_));
  OR2_X1    g141(.A1(new_n337_), .A2(new_n311_), .ZN(new_n343_));
  INV_X1    g142(.A(new_n341_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n280_), .A2(new_n311_), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n343_), .A2(KEYINPUT20), .A3(new_n344_), .A4(new_n345_), .ZN(new_n346_));
  NAND2_X1  g145(.A1(new_n342_), .A2(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348_));
  INV_X1    g147(.A(G92gat), .ZN(new_n349_));
  XNOR2_X1  g148(.A(new_n348_), .B(new_n349_), .ZN(new_n350_));
  XNOR2_X1  g149(.A(KEYINPUT18), .B(G64gat), .ZN(new_n351_));
  XOR2_X1   g150(.A(new_n350_), .B(new_n351_), .Z(new_n352_));
  NAND2_X1  g151(.A1(new_n347_), .A2(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(new_n352_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n342_), .A2(new_n354_), .A3(new_n346_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT27), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  XNOR2_X1  g157(.A(KEYINPUT100), .B(KEYINPUT20), .ZN(new_n359_));
  NAND3_X1  g158(.A1(new_n343_), .A2(new_n345_), .A3(new_n359_), .ZN(new_n360_));
  NAND2_X1  g159(.A1(new_n360_), .A2(new_n341_), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(new_n341_), .B2(new_n339_), .ZN(new_n362_));
  XOR2_X1   g161(.A(new_n352_), .B(KEYINPUT102), .Z(new_n363_));
  NAND2_X1  g162(.A1(new_n362_), .A2(new_n363_), .ZN(new_n364_));
  NAND3_X1  g163(.A1(new_n364_), .A2(KEYINPUT27), .A3(new_n355_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n358_), .A2(new_n365_), .ZN(new_n366_));
  NOR2_X1   g165(.A1(new_n329_), .A2(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n259_), .A2(new_n292_), .A3(new_n367_), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n251_), .A2(new_n254_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n362_), .A2(KEYINPUT32), .A3(new_n354_), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n354_), .A2(KEYINPUT32), .ZN(new_n371_));
  INV_X1    g170(.A(new_n371_), .ZN(new_n372_));
  OAI211_X1 g171(.A(new_n369_), .B(new_n370_), .C1(new_n372_), .C2(new_n347_), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT33), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n254_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n375_), .A2(KEYINPUT97), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT97), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n254_), .A2(new_n377_), .A3(new_n374_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n376_), .A2(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(new_n247_), .A2(new_n241_), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT98), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n240_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n238_), .A2(new_n239_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n383_), .A2(KEYINPUT98), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n382_), .A2(new_n248_), .A3(new_n384_), .ZN(new_n385_));
  NAND3_X1  g184(.A1(new_n380_), .A2(new_n206_), .A3(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(KEYINPUT99), .ZN(new_n387_));
  INV_X1    g186(.A(KEYINPUT93), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n356_), .A2(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n353_), .A2(KEYINPUT93), .A3(new_n355_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n389_), .A2(new_n390_), .ZN(new_n391_));
  NAND4_X1  g190(.A1(new_n252_), .A2(KEYINPUT33), .A3(new_n253_), .A4(new_n249_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n387_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n373_), .B1(new_n379_), .B2(new_n393_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n257_), .ZN(new_n395_));
  NOR3_X1   g194(.A1(new_n395_), .A2(new_n328_), .A3(new_n255_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n366_), .ZN(new_n397_));
  AOI22_X1  g196(.A1(new_n394_), .A2(new_n328_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n368_), .B1(new_n398_), .B2(new_n292_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G15gat), .B(G22gat), .ZN(new_n400_));
  INV_X1    g199(.A(G1gat), .ZN(new_n401_));
  INV_X1    g200(.A(G8gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT14), .B1(new_n401_), .B2(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(new_n403_), .ZN(new_n404_));
  XNOR2_X1  g203(.A(G1gat), .B(G8gat), .ZN(new_n405_));
  XNOR2_X1  g204(.A(new_n404_), .B(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G29gat), .B(G36gat), .ZN(new_n407_));
  INV_X1    g206(.A(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G43gat), .B(G50gat), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n409_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n411_), .A2(new_n407_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n412_), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n406_), .B(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(G229gat), .A2(G233gat), .ZN(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n414_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT15), .ZN(new_n418_));
  XNOR2_X1  g217(.A(new_n413_), .B(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(new_n406_), .ZN(new_n420_));
  OR2_X1    g219(.A1(new_n406_), .A2(new_n413_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n417_), .B1(new_n422_), .B2(new_n416_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G113gat), .B(G141gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(G169gat), .B(G197gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(new_n424_), .B(new_n425_), .ZN(new_n426_));
  XNOR2_X1  g225(.A(new_n423_), .B(new_n426_), .ZN(new_n427_));
  AND2_X1   g226(.A1(new_n399_), .A2(new_n427_), .ZN(new_n428_));
  INV_X1    g227(.A(G57gat), .ZN(new_n429_));
  INV_X1    g228(.A(G64gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(G57gat), .A2(G64gat), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n431_), .A2(new_n432_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n433_), .A2(KEYINPUT11), .ZN(new_n434_));
  XNOR2_X1  g233(.A(G71gat), .B(G78gat), .ZN(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT11), .ZN(new_n437_));
  NAND3_X1  g236(.A1(new_n431_), .A2(new_n437_), .A3(new_n432_), .ZN(new_n438_));
  NAND3_X1  g237(.A1(new_n434_), .A2(new_n436_), .A3(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n433_), .A2(new_n435_), .A3(KEYINPUT11), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n439_), .A2(new_n440_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n441_), .A2(KEYINPUT68), .ZN(new_n442_));
  INV_X1    g241(.A(KEYINPUT68), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n439_), .A2(new_n443_), .A3(new_n440_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n442_), .A2(KEYINPUT12), .A3(new_n444_), .ZN(new_n445_));
  INV_X1    g244(.A(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n448_));
  NOR2_X1   g247(.A1(new_n447_), .A2(new_n448_), .ZN(new_n449_));
  OR2_X1    g248(.A1(G85gat), .A2(G92gat), .ZN(new_n450_));
  NAND2_X1  g249(.A1(G85gat), .A2(G92gat), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  XNOR2_X1  g251(.A(KEYINPUT64), .B(KEYINPUT9), .ZN(new_n453_));
  OAI21_X1  g252(.A(new_n449_), .B1(new_n452_), .B2(new_n453_), .ZN(new_n454_));
  INV_X1    g253(.A(KEYINPUT9), .ZN(new_n455_));
  NAND3_X1  g254(.A1(new_n455_), .A2(G85gat), .A3(G92gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(KEYINPUT10), .B(G99gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n456_), .B1(new_n457_), .B2(G106gat), .ZN(new_n458_));
  OAI21_X1  g257(.A(KEYINPUT65), .B1(new_n454_), .B2(new_n458_), .ZN(new_n459_));
  NOR2_X1   g258(.A1(new_n451_), .A2(KEYINPUT9), .ZN(new_n460_));
  INV_X1    g259(.A(G99gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(KEYINPUT10), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT10), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(G99gat), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n462_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(G106gat), .ZN(new_n466_));
  AOI21_X1  g265(.A(new_n460_), .B1(new_n465_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT65), .ZN(new_n468_));
  AND2_X1   g267(.A1(new_n455_), .A2(KEYINPUT64), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n455_), .A2(KEYINPUT64), .ZN(new_n470_));
  OAI211_X1 g269(.A(new_n451_), .B(new_n450_), .C1(new_n469_), .C2(new_n470_), .ZN(new_n471_));
  NAND4_X1  g270(.A1(new_n467_), .A2(new_n468_), .A3(new_n471_), .A4(new_n449_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(new_n459_), .A2(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(KEYINPUT67), .ZN(new_n474_));
  INV_X1    g273(.A(KEYINPUT8), .ZN(new_n475_));
  OAI21_X1  g274(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n476_));
  INV_X1    g275(.A(new_n476_), .ZN(new_n477_));
  NOR3_X1   g276(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n477_), .A2(new_n478_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT6), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT66), .ZN(new_n483_));
  NAND3_X1  g282(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n482_), .A2(new_n483_), .A3(new_n484_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT66), .B1(new_n447_), .B2(new_n448_), .ZN(new_n486_));
  NAND3_X1  g285(.A1(new_n479_), .A2(new_n485_), .A3(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n452_), .ZN(new_n488_));
  AOI21_X1  g287(.A(new_n475_), .B1(new_n487_), .B2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n450_), .A2(new_n475_), .A3(new_n451_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n490_), .B1(new_n479_), .B2(new_n449_), .ZN(new_n491_));
  OAI211_X1 g290(.A(new_n473_), .B(new_n474_), .C1(new_n489_), .C2(new_n491_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(new_n491_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n483_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n495_));
  INV_X1    g294(.A(KEYINPUT7), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n496_), .A2(new_n461_), .A3(new_n466_), .ZN(new_n497_));
  NAND2_X1  g296(.A1(new_n497_), .A2(new_n476_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n495_), .A2(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n452_), .B1(new_n499_), .B2(new_n485_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n494_), .B1(new_n500_), .B2(new_n475_), .ZN(new_n501_));
  AOI21_X1  g300(.A(new_n474_), .B1(new_n501_), .B2(new_n473_), .ZN(new_n502_));
  OAI21_X1  g301(.A(new_n446_), .B1(new_n493_), .B2(new_n502_), .ZN(new_n503_));
  AND2_X1   g302(.A1(new_n459_), .A2(new_n472_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n487_), .A2(new_n488_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n491_), .B1(new_n505_), .B2(KEYINPUT8), .ZN(new_n506_));
  OAI211_X1 g305(.A(new_n440_), .B(new_n439_), .C1(new_n504_), .C2(new_n506_), .ZN(new_n507_));
  OAI211_X1 g306(.A(new_n473_), .B(new_n441_), .C1(new_n489_), .C2(new_n491_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n508_), .A2(KEYINPUT12), .ZN(new_n509_));
  AOI22_X1  g308(.A1(new_n503_), .A2(KEYINPUT69), .B1(new_n507_), .B2(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(G230gat), .A2(G233gat), .ZN(new_n511_));
  OAI21_X1  g310(.A(KEYINPUT67), .B1(new_n504_), .B2(new_n506_), .ZN(new_n512_));
  AOI211_X1 g311(.A(KEYINPUT69), .B(new_n445_), .C1(new_n512_), .C2(new_n492_), .ZN(new_n513_));
  INV_X1    g312(.A(new_n513_), .ZN(new_n514_));
  NAND3_X1  g313(.A1(new_n510_), .A2(new_n511_), .A3(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(new_n507_), .A2(new_n508_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n511_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  XNOR2_X1  g318(.A(G120gat), .B(G148gat), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n520_), .B(new_n305_), .ZN(new_n521_));
  XNOR2_X1  g320(.A(KEYINPUT5), .B(G176gat), .ZN(new_n522_));
  XOR2_X1   g321(.A(new_n521_), .B(new_n522_), .Z(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n519_), .A2(new_n524_), .ZN(new_n525_));
  INV_X1    g324(.A(KEYINPUT70), .ZN(new_n526_));
  NAND3_X1  g325(.A1(new_n515_), .A2(new_n518_), .A3(new_n523_), .ZN(new_n527_));
  NAND3_X1  g326(.A1(new_n525_), .A2(new_n526_), .A3(new_n527_), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n519_), .A2(KEYINPUT70), .A3(new_n524_), .ZN(new_n529_));
  AND2_X1   g328(.A1(new_n528_), .A2(new_n529_), .ZN(new_n530_));
  OR2_X1    g329(.A1(new_n530_), .A2(KEYINPUT13), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n530_), .A2(KEYINPUT13), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G127gat), .B(G155gat), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n535_), .B(KEYINPUT79), .ZN(new_n536_));
  XNOR2_X1  g335(.A(new_n536_), .B(KEYINPUT78), .ZN(new_n537_));
  XNOR2_X1  g336(.A(G183gat), .B(G211gat), .ZN(new_n538_));
  XNOR2_X1  g337(.A(new_n538_), .B(KEYINPUT16), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n537_), .B(new_n539_), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT17), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n541_), .B(KEYINPUT80), .Z(new_n542_));
  XNOR2_X1  g341(.A(new_n406_), .B(new_n441_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n545_), .A2(KEYINPUT68), .ZN(new_n546_));
  OR2_X1    g345(.A1(new_n545_), .A2(KEYINPUT68), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n542_), .A2(new_n546_), .A3(new_n547_), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n540_), .A2(KEYINPUT17), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n549_), .A2(new_n545_), .A3(new_n541_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n550_), .A2(KEYINPUT81), .ZN(new_n551_));
  OR2_X1    g350(.A1(new_n550_), .A2(KEYINPUT81), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n548_), .A2(new_n551_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n419_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n554_), .B1(new_n512_), .B2(new_n492_), .ZN(new_n555_));
  XOR2_X1   g354(.A(KEYINPUT71), .B(KEYINPUT34), .Z(new_n556_));
  NAND2_X1  g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT35), .ZN(new_n559_));
  NOR2_X1   g358(.A1(new_n558_), .A2(new_n559_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n413_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n473_), .B(new_n561_), .C1(new_n489_), .C2(new_n491_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n558_), .A2(new_n559_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n562_), .A2(new_n563_), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n555_), .A2(new_n560_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT73), .ZN(new_n566_));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n562_), .A2(new_n567_), .A3(new_n563_), .ZN(new_n568_));
  AOI21_X1  g367(.A(new_n567_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n569_));
  NOR3_X1   g368(.A1(new_n555_), .A2(new_n568_), .A3(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n560_), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n566_), .B1(new_n570_), .B2(new_n571_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n419_), .B1(new_n493_), .B2(new_n502_), .ZN(new_n573_));
  NAND3_X1  g372(.A1(new_n562_), .A2(new_n567_), .A3(new_n563_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n564_), .A2(KEYINPUT72), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n573_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n576_), .A2(KEYINPUT73), .A3(new_n560_), .ZN(new_n577_));
  AOI21_X1  g376(.A(new_n565_), .B1(new_n572_), .B2(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(G190gat), .B(G218gat), .Z(new_n579_));
  XNOR2_X1  g378(.A(G134gat), .B(G162gat), .ZN(new_n580_));
  XNOR2_X1  g379(.A(new_n579_), .B(new_n580_), .ZN(new_n581_));
  XNOR2_X1  g380(.A(new_n581_), .B(KEYINPUT36), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(KEYINPUT77), .B1(new_n578_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n565_), .ZN(new_n585_));
  AND3_X1   g384(.A1(new_n576_), .A2(KEYINPUT73), .A3(new_n560_), .ZN(new_n586_));
  AOI21_X1  g385(.A(KEYINPUT73), .B1(new_n576_), .B2(new_n560_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n585_), .B1(new_n586_), .B2(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT77), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(new_n582_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n584_), .A2(new_n590_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT36), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n581_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(KEYINPUT74), .B(KEYINPUT75), .Z(new_n594_));
  XNOR2_X1  g393(.A(new_n593_), .B(new_n594_), .ZN(new_n595_));
  OAI211_X1 g394(.A(new_n585_), .B(new_n595_), .C1(new_n586_), .C2(new_n587_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT76), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n572_), .A2(new_n577_), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT76), .ZN(new_n599_));
  NAND4_X1  g398(.A1(new_n598_), .A2(new_n599_), .A3(new_n585_), .A4(new_n595_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n597_), .A2(new_n600_), .ZN(new_n601_));
  OAI21_X1  g400(.A(KEYINPUT37), .B1(new_n591_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n588_), .A2(new_n582_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(new_n603_), .A2(new_n596_), .ZN(new_n604_));
  INV_X1    g403(.A(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(KEYINPUT37), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n602_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR3_X1   g408(.A1(new_n534_), .A2(new_n553_), .A3(new_n609_), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n610_), .A2(KEYINPUT82), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(KEYINPUT82), .ZN(new_n612_));
  AND3_X1   g411(.A1(new_n428_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n613_), .A2(KEYINPUT103), .ZN(new_n614_));
  NAND3_X1  g413(.A1(new_n428_), .A2(new_n611_), .A3(new_n612_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT103), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n614_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n401_), .A3(new_n258_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT38), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n618_), .A2(KEYINPUT38), .A3(new_n401_), .A4(new_n258_), .ZN(new_n622_));
  INV_X1    g421(.A(new_n427_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(new_n534_), .A2(new_n623_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n605_), .A2(new_n553_), .ZN(new_n625_));
  AND3_X1   g424(.A1(new_n399_), .A2(new_n624_), .A3(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(G1gat), .B1(new_n627_), .B2(new_n259_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n621_), .A2(new_n622_), .A3(new_n628_), .ZN(G1324gat));
  NAND2_X1  g428(.A1(new_n366_), .A2(new_n402_), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n614_), .B2(new_n617_), .ZN(new_n631_));
  INV_X1    g430(.A(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n626_), .A2(new_n366_), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n633_), .B1(new_n634_), .B2(G8gat), .ZN(new_n635_));
  AOI211_X1 g434(.A(KEYINPUT39), .B(new_n402_), .C1(new_n626_), .C2(new_n366_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n635_), .A2(new_n636_), .ZN(new_n637_));
  INV_X1    g436(.A(new_n637_), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n632_), .A2(KEYINPUT40), .A3(new_n638_), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT40), .ZN(new_n640_));
  OAI21_X1  g439(.A(new_n640_), .B1(new_n631_), .B2(new_n637_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n639_), .A2(new_n641_), .ZN(G1325gat));
  OAI21_X1  g441(.A(G15gat), .B1(new_n627_), .B2(new_n291_), .ZN(new_n643_));
  XNOR2_X1  g442(.A(new_n643_), .B(KEYINPUT41), .ZN(new_n644_));
  NOR3_X1   g443(.A1(new_n615_), .A2(G15gat), .A3(new_n291_), .ZN(new_n645_));
  OR2_X1    g444(.A1(new_n644_), .A2(new_n645_), .ZN(G1326gat));
  NOR2_X1   g445(.A1(new_n328_), .A2(G22gat), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT104), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n613_), .A2(new_n648_), .ZN(new_n649_));
  NAND2_X1  g448(.A1(new_n626_), .A2(new_n329_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT42), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n650_), .A2(new_n651_), .A3(G22gat), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n651_), .B1(new_n650_), .B2(G22gat), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n649_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT105), .ZN(new_n655_));
  XNOR2_X1  g454(.A(new_n654_), .B(new_n655_), .ZN(G1327gat));
  INV_X1    g455(.A(G29gat), .ZN(new_n657_));
  INV_X1    g456(.A(new_n553_), .ZN(new_n658_));
  NOR3_X1   g457(.A1(new_n534_), .A2(new_n658_), .A3(new_n623_), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  AND3_X1   g459(.A1(new_n399_), .A2(new_n660_), .A3(new_n609_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n660_), .B1(new_n399_), .B2(new_n609_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n659_), .B1(new_n661_), .B2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n664_));
  AOI211_X1 g463(.A(new_n657_), .B(new_n259_), .C1(new_n663_), .C2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(new_n659_), .ZN(new_n666_));
  NAND2_X1  g465(.A1(new_n399_), .A2(new_n609_), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n667_), .A2(KEYINPUT43), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n399_), .A2(new_n660_), .A3(new_n609_), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n666_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n670_), .A2(KEYINPUT44), .ZN(new_n671_));
  NAND3_X1  g470(.A1(new_n399_), .A2(new_n605_), .A3(new_n659_), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n673_));
  NAND2_X1  g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NAND4_X1  g473(.A1(new_n399_), .A2(KEYINPUT106), .A3(new_n605_), .A4(new_n659_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n258_), .A3(new_n675_), .ZN(new_n676_));
  AOI22_X1  g475(.A1(new_n665_), .A2(new_n671_), .B1(new_n657_), .B2(new_n676_), .ZN(G1328gat));
  INV_X1    g476(.A(KEYINPUT46), .ZN(new_n678_));
  INV_X1    g477(.A(G36gat), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n397_), .B1(new_n663_), .B2(new_n664_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n679_), .B1(new_n680_), .B2(new_n671_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n397_), .A2(G36gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n674_), .A2(new_n675_), .A3(new_n682_), .ZN(new_n683_));
  XNOR2_X1  g482(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n684_));
  XOR2_X1   g483(.A(new_n684_), .B(KEYINPUT108), .Z(new_n685_));
  INV_X1    g484(.A(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(new_n683_), .B(new_n686_), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n678_), .B1(new_n681_), .B2(new_n687_), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n366_), .B1(new_n670_), .B2(KEYINPUT44), .ZN(new_n689_));
  NOR2_X1   g488(.A1(new_n663_), .A2(new_n664_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G36gat), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n683_), .B(new_n685_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(new_n692_), .A3(KEYINPUT46), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n688_), .A2(new_n693_), .ZN(G1329gat));
  NAND3_X1  g493(.A1(new_n674_), .A2(new_n292_), .A3(new_n675_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(new_n288_), .ZN(new_n696_));
  OAI211_X1 g495(.A(G43gat), .B(new_n292_), .C1(new_n670_), .C2(KEYINPUT44), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n697_), .B2(new_n690_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n698_), .A2(KEYINPUT47), .ZN(new_n699_));
  INV_X1    g498(.A(KEYINPUT47), .ZN(new_n700_));
  OAI211_X1 g499(.A(new_n700_), .B(new_n696_), .C1(new_n697_), .C2(new_n690_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(G1330gat));
  NAND3_X1  g501(.A1(new_n674_), .A2(new_n329_), .A3(new_n675_), .ZN(new_n703_));
  INV_X1    g502(.A(G50gat), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OAI211_X1 g504(.A(G50gat), .B(new_n329_), .C1(new_n670_), .C2(KEYINPUT44), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n705_), .B1(new_n706_), .B2(new_n690_), .ZN(new_n707_));
  INV_X1    g506(.A(KEYINPUT109), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  OAI211_X1 g508(.A(KEYINPUT109), .B(new_n705_), .C1(new_n706_), .C2(new_n690_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1331gat));
  NOR2_X1   g510(.A1(new_n533_), .A2(new_n427_), .ZN(new_n712_));
  AND2_X1   g511(.A1(new_n399_), .A2(new_n712_), .ZN(new_n713_));
  AND3_X1   g512(.A1(new_n713_), .A2(new_n658_), .A3(new_n608_), .ZN(new_n714_));
  AOI21_X1  g513(.A(G57gat), .B1(new_n714_), .B2(new_n258_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n713_), .A2(new_n625_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n259_), .A2(new_n429_), .ZN(new_n717_));
  AOI21_X1  g516(.A(new_n715_), .B1(new_n716_), .B2(new_n717_), .ZN(G1332gat));
  AOI21_X1  g517(.A(new_n430_), .B1(new_n716_), .B2(new_n366_), .ZN(new_n719_));
  XOR2_X1   g518(.A(new_n719_), .B(KEYINPUT48), .Z(new_n720_));
  NAND3_X1  g519(.A1(new_n714_), .A2(new_n430_), .A3(new_n366_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1333gat));
  INV_X1    g521(.A(G71gat), .ZN(new_n723_));
  AOI21_X1  g522(.A(new_n723_), .B1(new_n716_), .B2(new_n292_), .ZN(new_n724_));
  XOR2_X1   g523(.A(new_n724_), .B(KEYINPUT49), .Z(new_n725_));
  NAND3_X1  g524(.A1(new_n714_), .A2(new_n723_), .A3(new_n292_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1334gat));
  INV_X1    g526(.A(G78gat), .ZN(new_n728_));
  AOI21_X1  g527(.A(new_n728_), .B1(new_n716_), .B2(new_n329_), .ZN(new_n729_));
  XOR2_X1   g528(.A(new_n729_), .B(KEYINPUT50), .Z(new_n730_));
  NOR2_X1   g529(.A1(new_n328_), .A2(G78gat), .ZN(new_n731_));
  XNOR2_X1  g530(.A(new_n731_), .B(KEYINPUT110), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n714_), .A2(new_n732_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n730_), .A2(new_n733_), .ZN(G1335gat));
  NAND2_X1  g533(.A1(new_n712_), .A2(new_n553_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n399_), .A2(new_n605_), .A3(new_n736_), .ZN(new_n737_));
  AOI21_X1  g536(.A(G85gat), .B1(new_n737_), .B2(new_n258_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n735_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n258_), .A2(G85gat), .ZN(new_n740_));
  XNOR2_X1  g539(.A(new_n740_), .B(KEYINPUT111), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n738_), .B1(new_n739_), .B2(new_n741_), .ZN(G1336gat));
  AOI21_X1  g541(.A(G92gat), .B1(new_n737_), .B2(new_n366_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n397_), .A2(new_n349_), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n743_), .B1(new_n739_), .B2(new_n744_), .ZN(G1337gat));
  NAND3_X1  g544(.A1(new_n737_), .A2(new_n465_), .A3(new_n292_), .ZN(new_n746_));
  AND2_X1   g545(.A1(new_n746_), .A2(KEYINPUT112), .ZN(new_n747_));
  AND2_X1   g546(.A1(new_n739_), .A2(new_n292_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n747_), .B1(new_n748_), .B2(new_n461_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(KEYINPUT51), .ZN(new_n750_));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n751_));
  OAI211_X1 g550(.A(new_n751_), .B(new_n747_), .C1(new_n748_), .C2(new_n461_), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n750_), .A2(new_n752_), .ZN(G1338gat));
  NAND3_X1  g552(.A1(new_n737_), .A2(new_n466_), .A3(new_n329_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n329_), .B(new_n736_), .C1(new_n661_), .C2(new_n662_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n756_));
  AND3_X1   g555(.A1(new_n755_), .A2(new_n756_), .A3(G106gat), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n756_), .B1(new_n755_), .B2(G106gat), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n754_), .B1(new_n757_), .B2(new_n758_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n759_), .A2(KEYINPUT53), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n761_));
  OAI211_X1 g560(.A(new_n761_), .B(new_n754_), .C1(new_n757_), .C2(new_n758_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n760_), .A2(new_n762_), .ZN(G1339gat));
  NAND4_X1  g562(.A1(new_n533_), .A2(new_n658_), .A3(new_n608_), .A4(new_n623_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(KEYINPUT113), .B(KEYINPUT54), .ZN(new_n765_));
  INV_X1    g564(.A(new_n765_), .ZN(new_n766_));
  XNOR2_X1  g565(.A(new_n764_), .B(new_n766_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n527_), .A2(new_n427_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n509_), .A2(new_n507_), .ZN(new_n769_));
  AOI21_X1  g568(.A(new_n445_), .B1(new_n512_), .B2(new_n492_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT69), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n769_), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  NOR3_X1   g571(.A1(new_n772_), .A2(new_n517_), .A3(new_n513_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n517_), .B1(new_n772_), .B2(new_n513_), .ZN(new_n774_));
  AOI21_X1  g573(.A(new_n773_), .B1(KEYINPUT55), .B2(new_n774_), .ZN(new_n775_));
  AND4_X1   g574(.A1(KEYINPUT55), .A2(new_n510_), .A3(new_n511_), .A4(new_n514_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n524_), .B1(new_n775_), .B2(new_n776_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT56), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n777_), .A2(new_n778_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n774_), .A2(KEYINPUT55), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n780_), .A2(new_n515_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n773_), .A2(new_n774_), .A3(KEYINPUT55), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n524_), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n768_), .B1(new_n779_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT114), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n416_), .B1(new_n422_), .B2(new_n786_), .ZN(new_n787_));
  AOI21_X1  g586(.A(KEYINPUT114), .B1(new_n420_), .B2(new_n421_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n414_), .A2(new_n415_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n790_), .A2(new_n426_), .ZN(new_n791_));
  OAI22_X1  g590(.A1(new_n789_), .A2(new_n791_), .B1(new_n423_), .B2(new_n426_), .ZN(new_n792_));
  XNOR2_X1  g591(.A(new_n792_), .B(KEYINPUT115), .ZN(new_n793_));
  NAND3_X1  g592(.A1(new_n528_), .A2(new_n793_), .A3(new_n529_), .ZN(new_n794_));
  INV_X1    g593(.A(new_n794_), .ZN(new_n795_));
  OAI21_X1  g594(.A(new_n604_), .B1(new_n785_), .B2(new_n795_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT57), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n796_), .A2(new_n797_), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n779_), .A2(new_n784_), .ZN(new_n799_));
  AND2_X1   g598(.A1(new_n793_), .A2(new_n527_), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT58), .B1(new_n799_), .B2(new_n800_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n801_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n799_), .A2(KEYINPUT58), .A3(new_n800_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n802_), .A2(new_n609_), .A3(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n768_), .ZN(new_n805_));
  AOI21_X1  g604(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n524_), .ZN(new_n806_));
  AOI211_X1 g605(.A(new_n778_), .B(new_n523_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n807_));
  OAI21_X1  g606(.A(new_n805_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n605_), .B1(new_n808_), .B2(new_n794_), .ZN(new_n809_));
  AOI21_X1  g608(.A(KEYINPUT116), .B1(new_n809_), .B2(KEYINPUT57), .ZN(new_n810_));
  OAI211_X1 g609(.A(KEYINPUT57), .B(new_n604_), .C1(new_n785_), .C2(new_n795_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  OAI211_X1 g612(.A(new_n798_), .B(new_n804_), .C1(new_n810_), .C2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n658_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n801_), .A2(new_n608_), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n817_), .A2(new_n803_), .B1(new_n797_), .B2(new_n796_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n811_), .A2(new_n812_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n808_), .A2(new_n794_), .ZN(new_n820_));
  NAND4_X1  g619(.A1(new_n820_), .A2(KEYINPUT116), .A3(KEYINPUT57), .A4(new_n604_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n818_), .A2(KEYINPUT117), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n767_), .B1(new_n816_), .B2(new_n823_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n367_), .A2(new_n258_), .A3(new_n292_), .ZN(new_n825_));
  OAI21_X1  g624(.A(KEYINPUT118), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n827_));
  INV_X1    g626(.A(new_n825_), .ZN(new_n828_));
  AND3_X1   g627(.A1(new_n818_), .A2(KEYINPUT117), .A3(new_n822_), .ZN(new_n829_));
  AOI21_X1  g628(.A(KEYINPUT117), .B1(new_n818_), .B2(new_n822_), .ZN(new_n830_));
  NOR3_X1   g629(.A1(new_n829_), .A2(new_n830_), .A3(new_n658_), .ZN(new_n831_));
  OAI211_X1 g630(.A(new_n827_), .B(new_n828_), .C1(new_n831_), .C2(new_n767_), .ZN(new_n832_));
  NAND2_X1  g631(.A1(new_n826_), .A2(new_n832_), .ZN(new_n833_));
  AOI21_X1  g632(.A(G113gat), .B1(new_n833_), .B2(new_n427_), .ZN(new_n834_));
  NOR2_X1   g633(.A1(new_n810_), .A2(new_n813_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n804_), .A2(new_n798_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n815_), .B1(new_n835_), .B2(new_n836_), .ZN(new_n837_));
  NAND3_X1  g636(.A1(new_n837_), .A2(new_n553_), .A3(new_n823_), .ZN(new_n838_));
  INV_X1    g637(.A(new_n767_), .ZN(new_n839_));
  AOI21_X1  g638(.A(new_n825_), .B1(new_n838_), .B2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841_));
  NOR2_X1   g640(.A1(new_n840_), .A2(new_n841_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n814_), .A2(new_n553_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n839_), .A2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n825_), .A2(KEYINPUT59), .ZN(new_n845_));
  AOI21_X1  g644(.A(new_n842_), .B1(new_n844_), .B2(new_n845_), .ZN(new_n846_));
  AND2_X1   g645(.A1(new_n427_), .A2(G113gat), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n834_), .B1(new_n846_), .B2(new_n847_), .ZN(G1340gat));
  NAND2_X1  g647(.A1(new_n844_), .A2(new_n845_), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n534_), .B(new_n849_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n850_));
  XOR2_X1   g649(.A(KEYINPUT119), .B(G120gat), .Z(new_n851_));
  NAND2_X1  g650(.A1(new_n850_), .A2(new_n851_), .ZN(new_n852_));
  NOR2_X1   g651(.A1(new_n533_), .A2(KEYINPUT60), .ZN(new_n853_));
  MUX2_X1   g652(.A(new_n853_), .B(KEYINPUT60), .S(new_n851_), .Z(new_n854_));
  NAND2_X1  g653(.A1(new_n838_), .A2(new_n839_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n827_), .B1(new_n855_), .B2(new_n828_), .ZN(new_n856_));
  AOI211_X1 g655(.A(KEYINPUT118), .B(new_n825_), .C1(new_n838_), .C2(new_n839_), .ZN(new_n857_));
  OAI21_X1  g656(.A(new_n854_), .B1(new_n856_), .B2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n852_), .A2(new_n858_), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n859_), .A2(KEYINPUT120), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861_));
  NAND3_X1  g660(.A1(new_n852_), .A2(new_n858_), .A3(new_n861_), .ZN(new_n862_));
  NAND2_X1  g661(.A1(new_n860_), .A2(new_n862_), .ZN(G1341gat));
  AOI21_X1  g662(.A(G127gat), .B1(new_n833_), .B2(new_n658_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n658_), .A2(G127gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n865_), .B(KEYINPUT121), .ZN(new_n866_));
  AOI21_X1  g665(.A(new_n864_), .B1(new_n846_), .B2(new_n866_), .ZN(G1342gat));
  AOI21_X1  g666(.A(G134gat), .B1(new_n833_), .B2(new_n605_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n609_), .A2(G134gat), .ZN(new_n869_));
  OAI211_X1 g668(.A(new_n849_), .B(new_n869_), .C1(new_n840_), .C2(new_n841_), .ZN(new_n870_));
  INV_X1    g669(.A(new_n870_), .ZN(new_n871_));
  OAI21_X1  g670(.A(KEYINPUT122), .B1(new_n868_), .B2(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(KEYINPUT122), .ZN(new_n873_));
  AOI21_X1  g672(.A(new_n604_), .B1(new_n826_), .B2(new_n832_), .ZN(new_n874_));
  OAI211_X1 g673(.A(new_n873_), .B(new_n870_), .C1(new_n874_), .C2(G134gat), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n872_), .A2(new_n875_), .ZN(G1343gat));
  NOR3_X1   g675(.A1(new_n259_), .A2(new_n328_), .A3(new_n366_), .ZN(new_n877_));
  AND3_X1   g676(.A1(new_n855_), .A2(new_n291_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n427_), .ZN(new_n879_));
  XNOR2_X1  g678(.A(new_n879_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n534_), .ZN(new_n881_));
  XNOR2_X1  g680(.A(new_n881_), .B(G148gat), .ZN(G1345gat));
  NAND4_X1  g681(.A1(new_n855_), .A2(new_n658_), .A3(new_n291_), .A4(new_n877_), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n883_), .A2(KEYINPUT123), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(KEYINPUT123), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  XNOR2_X1  g685(.A(KEYINPUT61), .B(G155gat), .ZN(new_n887_));
  INV_X1    g686(.A(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n884_), .A2(new_n885_), .A3(new_n887_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n889_), .A2(new_n890_), .ZN(G1346gat));
  AOI21_X1  g690(.A(G162gat), .B1(new_n878_), .B2(new_n605_), .ZN(new_n892_));
  AND2_X1   g691(.A1(new_n609_), .A2(G162gat), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n878_), .B2(new_n893_), .ZN(G1347gat));
  INV_X1    g693(.A(KEYINPUT62), .ZN(new_n895_));
  NOR4_X1   g694(.A1(new_n258_), .A2(new_n329_), .A3(new_n397_), .A4(new_n291_), .ZN(new_n896_));
  AND2_X1   g695(.A1(new_n844_), .A2(new_n896_), .ZN(new_n897_));
  NAND2_X1  g696(.A1(new_n897_), .A2(new_n427_), .ZN(new_n898_));
  INV_X1    g697(.A(new_n898_), .ZN(new_n899_));
  OAI21_X1  g698(.A(new_n895_), .B1(new_n899_), .B2(new_n270_), .ZN(new_n900_));
  NAND3_X1  g699(.A1(new_n898_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n899_), .A2(new_n262_), .ZN(new_n902_));
  NAND3_X1  g701(.A1(new_n900_), .A2(new_n901_), .A3(new_n902_), .ZN(G1348gat));
  AOI21_X1  g702(.A(G176gat), .B1(new_n897_), .B2(new_n534_), .ZN(new_n904_));
  AND3_X1   g703(.A1(new_n896_), .A2(G176gat), .A3(new_n534_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n904_), .B1(new_n855_), .B2(new_n905_), .ZN(G1349gat));
  NAND2_X1  g705(.A1(new_n897_), .A2(new_n658_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n907_), .A2(G183gat), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n276_), .B2(new_n907_), .ZN(G1350gat));
  NAND2_X1  g708(.A1(new_n897_), .A2(new_n609_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(G190gat), .ZN(new_n911_));
  OR2_X1    g710(.A1(new_n604_), .A2(new_n335_), .ZN(new_n912_));
  XNOR2_X1  g711(.A(new_n912_), .B(KEYINPUT124), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n897_), .A2(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n911_), .A2(new_n914_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT125), .ZN(new_n916_));
  INV_X1    g715(.A(KEYINPUT125), .ZN(new_n917_));
  NAND3_X1  g716(.A1(new_n911_), .A2(new_n917_), .A3(new_n914_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n916_), .A2(new_n918_), .ZN(G1351gat));
  NOR3_X1   g718(.A1(new_n258_), .A2(new_n328_), .A3(new_n397_), .ZN(new_n920_));
  NAND3_X1  g719(.A1(new_n855_), .A2(new_n291_), .A3(new_n920_), .ZN(new_n921_));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(new_n923_));
  NAND4_X1  g722(.A1(new_n855_), .A2(KEYINPUT126), .A3(new_n291_), .A4(new_n920_), .ZN(new_n924_));
  NAND2_X1  g723(.A1(new_n923_), .A2(new_n924_), .ZN(new_n925_));
  AOI21_X1  g724(.A(G197gat), .B1(new_n925_), .B2(new_n427_), .ZN(new_n926_));
  AOI211_X1 g725(.A(new_n302_), .B(new_n623_), .C1(new_n923_), .C2(new_n924_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(new_n926_), .A2(new_n927_), .ZN(G1352gat));
  NAND2_X1  g727(.A1(new_n925_), .A2(new_n534_), .ZN(new_n929_));
  NAND2_X1  g728(.A1(new_n929_), .A2(G204gat), .ZN(new_n930_));
  NAND3_X1  g729(.A1(new_n925_), .A2(new_n305_), .A3(new_n534_), .ZN(new_n931_));
  NAND2_X1  g730(.A1(new_n930_), .A2(new_n931_), .ZN(G1353gat));
  AOI21_X1  g731(.A(new_n553_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n933_));
  NAND2_X1  g732(.A1(new_n925_), .A2(new_n933_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(KEYINPUT127), .ZN(new_n936_));
  INV_X1    g735(.A(new_n936_), .ZN(new_n937_));
  NAND2_X1  g736(.A1(new_n934_), .A2(new_n937_), .ZN(new_n938_));
  NAND3_X1  g737(.A1(new_n925_), .A2(new_n936_), .A3(new_n933_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n938_), .A2(new_n939_), .ZN(G1354gat));
  NAND2_X1  g739(.A1(new_n925_), .A2(new_n605_), .ZN(new_n941_));
  INV_X1    g740(.A(G218gat), .ZN(new_n942_));
  NOR2_X1   g741(.A1(new_n608_), .A2(new_n942_), .ZN(new_n943_));
  AOI22_X1  g742(.A1(new_n941_), .A2(new_n942_), .B1(new_n925_), .B2(new_n943_), .ZN(G1355gat));
endmodule


