//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 0 1 0 1 1 1 1 1 0 1 0 1 0 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n709_, new_n710_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n822_, new_n823_, new_n824_, new_n825_, new_n826_, new_n828_,
    new_n829_, new_n831_, new_n832_, new_n834_, new_n835_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n849_, new_n850_,
    new_n851_, new_n853_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n861_, new_n862_, new_n864_,
    new_n865_, new_n866_, new_n867_, new_n868_, new_n869_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n883_, new_n884_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n893_, new_n894_;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202_));
  NAND2_X1  g001(.A1(G232gat), .A2(G233gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT34), .ZN(new_n204_));
  AND2_X1   g003(.A1(new_n204_), .A2(KEYINPUT35), .ZN(new_n205_));
  NOR2_X1   g004(.A1(new_n204_), .A2(KEYINPUT35), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n205_), .A2(new_n206_), .ZN(new_n207_));
  INV_X1    g006(.A(KEYINPUT68), .ZN(new_n208_));
  XNOR2_X1  g007(.A(G85gat), .B(G92gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT6), .ZN(new_n211_));
  XNOR2_X1  g010(.A(new_n210_), .B(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT66), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n213_), .A2(KEYINPUT7), .ZN(new_n214_));
  NOR2_X1   g013(.A1(G99gat), .A2(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(KEYINPUT7), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n216_), .B1(new_n217_), .B2(new_n215_), .ZN(new_n218_));
  AOI21_X1  g017(.A(new_n212_), .B1(new_n218_), .B2(KEYINPUT67), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n220_));
  OAI211_X1 g019(.A(new_n220_), .B(new_n216_), .C1(new_n217_), .C2(new_n215_), .ZN(new_n221_));
  AOI21_X1  g020(.A(new_n209_), .B1(new_n219_), .B2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n208_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT66), .ZN(new_n226_));
  AOI21_X1  g025(.A(new_n215_), .B1(new_n214_), .B2(new_n226_), .ZN(new_n227_));
  AOI211_X1 g026(.A(G99gat), .B(G106gat), .C1(new_n213_), .C2(KEYINPUT7), .ZN(new_n228_));
  OAI21_X1  g027(.A(KEYINPUT67), .B1(new_n227_), .B2(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(new_n212_), .ZN(new_n230_));
  NAND3_X1  g029(.A1(new_n229_), .A2(new_n230_), .A3(new_n221_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n209_), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(KEYINPUT68), .A3(KEYINPUT8), .ZN(new_n234_));
  OAI211_X1 g033(.A(new_n223_), .B(new_n232_), .C1(new_n218_), .C2(new_n212_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n224_), .A2(new_n234_), .A3(new_n235_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(KEYINPUT9), .ZN(new_n237_));
  XOR2_X1   g036(.A(KEYINPUT10), .B(G99gat), .Z(new_n238_));
  INV_X1    g037(.A(G106gat), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(G85gat), .ZN(new_n241_));
  INV_X1    g040(.A(G92gat), .ZN(new_n242_));
  OR3_X1    g041(.A1(new_n241_), .A2(new_n242_), .A3(KEYINPUT9), .ZN(new_n243_));
  NAND4_X1  g042(.A1(new_n237_), .A2(new_n230_), .A3(new_n240_), .A4(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(G29gat), .B(G36gat), .ZN(new_n245_));
  XNOR2_X1  g044(.A(new_n245_), .B(KEYINPUT70), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G43gat), .B(G50gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(new_n246_), .B(new_n247_), .ZN(new_n248_));
  INV_X1    g047(.A(new_n248_), .ZN(new_n249_));
  XOR2_X1   g048(.A(KEYINPUT71), .B(KEYINPUT15), .Z(new_n250_));
  NAND2_X1  g049(.A1(new_n249_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(new_n250_), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n248_), .A2(new_n252_), .ZN(new_n253_));
  AOI22_X1  g052(.A1(new_n236_), .A2(new_n244_), .B1(new_n251_), .B2(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n223_), .B1(new_n231_), .B2(new_n232_), .ZN(new_n255_));
  OAI21_X1  g054(.A(new_n235_), .B1(new_n255_), .B2(KEYINPUT68), .ZN(new_n256_));
  AOI211_X1 g055(.A(new_n208_), .B(new_n223_), .C1(new_n231_), .C2(new_n232_), .ZN(new_n257_));
  OAI211_X1 g056(.A(new_n244_), .B(new_n248_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(new_n258_), .ZN(new_n259_));
  OAI21_X1  g058(.A(new_n207_), .B1(new_n254_), .B2(new_n259_), .ZN(new_n260_));
  INV_X1    g059(.A(KEYINPUT73), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  OAI211_X1 g061(.A(KEYINPUT73), .B(new_n207_), .C1(new_n254_), .C2(new_n259_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n251_), .A2(new_n253_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n244_), .B1(new_n256_), .B2(new_n257_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n265_), .A2(new_n266_), .ZN(new_n267_));
  NAND3_X1  g066(.A1(new_n267_), .A2(new_n258_), .A3(new_n205_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n268_), .A2(KEYINPUT72), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n270_));
  NAND4_X1  g069(.A1(new_n267_), .A2(new_n270_), .A3(new_n258_), .A4(new_n205_), .ZN(new_n271_));
  NAND2_X1  g070(.A1(new_n269_), .A2(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(G190gat), .B(G218gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(G134gat), .B(G162gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  NOR2_X1   g074(.A1(new_n275_), .A2(KEYINPUT36), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n264_), .A2(new_n272_), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT37), .ZN(new_n278_));
  AOI22_X1  g077(.A1(new_n262_), .A2(new_n263_), .B1(new_n269_), .B2(new_n271_), .ZN(new_n279_));
  XOR2_X1   g078(.A(new_n275_), .B(KEYINPUT36), .Z(new_n280_));
  INV_X1    g079(.A(new_n280_), .ZN(new_n281_));
  OAI211_X1 g080(.A(new_n277_), .B(new_n278_), .C1(new_n279_), .C2(new_n281_), .ZN(new_n282_));
  NAND2_X1  g081(.A1(new_n282_), .A2(KEYINPUT75), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n264_), .A2(new_n272_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n284_), .A2(new_n280_), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT75), .ZN(new_n286_));
  NAND4_X1  g085(.A1(new_n285_), .A2(new_n286_), .A3(new_n278_), .A4(new_n277_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(new_n277_), .A2(KEYINPUT74), .ZN(new_n288_));
  NOR2_X1   g087(.A1(new_n288_), .A2(new_n278_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n285_), .A2(KEYINPUT74), .A3(new_n277_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n283_), .A2(new_n287_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  XNOR2_X1  g090(.A(G57gat), .B(G64gat), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n292_), .A2(KEYINPUT11), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(KEYINPUT11), .ZN(new_n294_));
  XOR2_X1   g093(.A(G71gat), .B(G78gat), .Z(new_n295_));
  NAND3_X1  g094(.A1(new_n293_), .A2(new_n294_), .A3(new_n295_), .ZN(new_n296_));
  OR2_X1    g095(.A1(new_n294_), .A2(new_n295_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n296_), .A2(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G231gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  XNOR2_X1  g099(.A(G15gat), .B(G22gat), .ZN(new_n301_));
  XNOR2_X1  g100(.A(KEYINPUT76), .B(G8gat), .ZN(new_n302_));
  AND2_X1   g101(.A1(new_n302_), .A2(G1gat), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT14), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n301_), .B1(new_n303_), .B2(new_n304_), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G1gat), .B(G8gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XNOR2_X1  g106(.A(new_n300_), .B(new_n307_), .ZN(new_n308_));
  NOR2_X1   g107(.A1(new_n308_), .A2(KEYINPUT79), .ZN(new_n309_));
  XNOR2_X1  g108(.A(G183gat), .B(G211gat), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n310_), .B(KEYINPUT78), .ZN(new_n311_));
  XOR2_X1   g110(.A(G127gat), .B(G155gat), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(KEYINPUT77), .B(KEYINPUT16), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n313_), .B(new_n314_), .ZN(new_n315_));
  NAND2_X1  g114(.A1(new_n315_), .A2(KEYINPUT17), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n309_), .B(new_n316_), .Z(new_n317_));
  NOR2_X1   g116(.A1(new_n315_), .A2(KEYINPUT17), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n308_), .A2(new_n318_), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n317_), .A2(new_n319_), .ZN(new_n320_));
  XNOR2_X1  g119(.A(new_n320_), .B(KEYINPUT80), .ZN(new_n321_));
  INV_X1    g120(.A(new_n321_), .ZN(new_n322_));
  NOR2_X1   g121(.A1(new_n291_), .A2(new_n322_), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT81), .ZN(new_n324_));
  OAI211_X1 g123(.A(new_n244_), .B(new_n298_), .C1(new_n256_), .C2(new_n257_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT64), .B(KEYINPUT65), .ZN(new_n326_));
  NAND2_X1  g125(.A1(G230gat), .A2(G233gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n326_), .B(new_n327_), .ZN(new_n328_));
  NAND2_X1  g127(.A1(new_n325_), .A2(new_n328_), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n329_), .A2(KEYINPUT69), .ZN(new_n330_));
  INV_X1    g129(.A(KEYINPUT69), .ZN(new_n331_));
  NAND3_X1  g130(.A1(new_n325_), .A2(new_n331_), .A3(new_n328_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT12), .ZN(new_n333_));
  INV_X1    g132(.A(new_n298_), .ZN(new_n334_));
  AOI21_X1  g133(.A(new_n333_), .B1(new_n266_), .B2(new_n334_), .ZN(new_n335_));
  AOI211_X1 g134(.A(KEYINPUT12), .B(new_n298_), .C1(new_n236_), .C2(new_n244_), .ZN(new_n336_));
  OAI211_X1 g135(.A(new_n330_), .B(new_n332_), .C1(new_n335_), .C2(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n266_), .A2(new_n334_), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n338_), .A2(new_n325_), .ZN(new_n339_));
  INV_X1    g138(.A(new_n328_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n337_), .A2(new_n341_), .ZN(new_n342_));
  XNOR2_X1  g141(.A(G120gat), .B(G148gat), .ZN(new_n343_));
  XNOR2_X1  g142(.A(new_n343_), .B(KEYINPUT5), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G176gat), .B(G204gat), .ZN(new_n345_));
  XOR2_X1   g144(.A(new_n344_), .B(new_n345_), .Z(new_n346_));
  INV_X1    g145(.A(new_n346_), .ZN(new_n347_));
  XNOR2_X1  g146(.A(new_n342_), .B(new_n347_), .ZN(new_n348_));
  OR2_X1    g147(.A1(new_n348_), .A2(KEYINPUT13), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(KEYINPUT13), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n323_), .A2(new_n324_), .A3(new_n352_), .ZN(new_n353_));
  NOR2_X1   g152(.A1(G155gat), .A2(G162gat), .ZN(new_n354_));
  XNOR2_X1  g153(.A(new_n354_), .B(KEYINPUT89), .ZN(new_n355_));
  INV_X1    g154(.A(G155gat), .ZN(new_n356_));
  INV_X1    g155(.A(G162gat), .ZN(new_n357_));
  NOR2_X1   g156(.A1(new_n356_), .A2(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  NOR2_X1   g159(.A1(G141gat), .A2(G148gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(new_n361_), .B(KEYINPUT3), .ZN(new_n362_));
  NAND2_X1  g161(.A1(G141gat), .A2(G148gat), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT2), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n360_), .A2(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n359_), .A2(KEYINPUT1), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT1), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n358_), .A2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n355_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT88), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n361_), .A2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(KEYINPUT88), .B1(G141gat), .B2(G148gat), .ZN(new_n373_));
  AOI22_X1  g172(.A1(new_n372_), .A2(new_n373_), .B1(G141gat), .B2(G148gat), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n370_), .A2(new_n374_), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n366_), .A2(new_n375_), .ZN(new_n376_));
  XOR2_X1   g175(.A(G127gat), .B(G134gat), .Z(new_n377_));
  XOR2_X1   g176(.A(G113gat), .B(G120gat), .Z(new_n378_));
  XOR2_X1   g177(.A(new_n377_), .B(new_n378_), .Z(new_n379_));
  NAND2_X1  g178(.A1(new_n376_), .A2(new_n379_), .ZN(new_n380_));
  AOI22_X1  g179(.A1(new_n365_), .A2(new_n360_), .B1(new_n370_), .B2(new_n374_), .ZN(new_n381_));
  INV_X1    g180(.A(new_n379_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(G225gat), .A2(G233gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n387_), .B(G85gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(KEYINPUT0), .B(G57gat), .ZN(new_n389_));
  XOR2_X1   g188(.A(new_n388_), .B(new_n389_), .Z(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n380_), .A2(new_n383_), .A3(KEYINPUT4), .ZN(new_n392_));
  OR3_X1    g191(.A1(new_n381_), .A2(new_n382_), .A3(KEYINPUT4), .ZN(new_n393_));
  AND2_X1   g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  OAI211_X1 g193(.A(new_n386_), .B(new_n391_), .C1(new_n394_), .C2(new_n385_), .ZN(new_n395_));
  AOI21_X1  g194(.A(new_n385_), .B1(new_n392_), .B2(new_n393_), .ZN(new_n396_));
  INV_X1    g195(.A(new_n386_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n390_), .B1(new_n396_), .B2(new_n397_), .ZN(new_n398_));
  INV_X1    g197(.A(KEYINPUT98), .ZN(new_n399_));
  NAND3_X1  g198(.A1(new_n395_), .A2(new_n398_), .A3(new_n399_), .ZN(new_n400_));
  OAI211_X1 g199(.A(KEYINPUT98), .B(new_n390_), .C1(new_n396_), .C2(new_n397_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n400_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(new_n402_), .ZN(new_n403_));
  AND3_X1   g202(.A1(KEYINPUT23), .A2(G183gat), .A3(G190gat), .ZN(new_n404_));
  AOI21_X1  g203(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n405_));
  NOR2_X1   g204(.A1(G183gat), .A2(G190gat), .ZN(new_n406_));
  OR3_X1    g205(.A1(new_n404_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  NAND2_X1  g206(.A1(G169gat), .A2(G176gat), .ZN(new_n408_));
  NAND2_X1  g207(.A1(new_n407_), .A2(new_n408_), .ZN(new_n409_));
  INV_X1    g208(.A(KEYINPUT22), .ZN(new_n410_));
  NAND2_X1  g209(.A1(new_n410_), .A2(G169gat), .ZN(new_n411_));
  AOI21_X1  g210(.A(G176gat), .B1(new_n411_), .B2(KEYINPUT85), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT22), .B(G169gat), .ZN(new_n413_));
  OAI21_X1  g212(.A(new_n412_), .B1(KEYINPUT85), .B2(new_n413_), .ZN(new_n414_));
  OR2_X1    g213(.A1(new_n414_), .A2(KEYINPUT86), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(KEYINPUT86), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n409_), .B1(new_n415_), .B2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(new_n417_), .ZN(new_n418_));
  NOR2_X1   g217(.A1(G169gat), .A2(G176gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT84), .ZN(new_n420_));
  AND2_X1   g219(.A1(new_n408_), .A2(KEYINPUT24), .ZN(new_n421_));
  OR2_X1    g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(KEYINPUT24), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n422_), .A2(new_n423_), .ZN(new_n424_));
  XNOR2_X1  g223(.A(KEYINPUT25), .B(G183gat), .ZN(new_n425_));
  XNOR2_X1  g224(.A(KEYINPUT26), .B(G190gat), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  NOR2_X1   g226(.A1(new_n404_), .A2(new_n405_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n427_), .A2(new_n428_), .ZN(new_n429_));
  INV_X1    g228(.A(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n424_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n418_), .A2(new_n431_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(G227gat), .A2(G233gat), .ZN(new_n433_));
  INV_X1    g232(.A(G71gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(G99gat), .ZN(new_n436_));
  XNOR2_X1  g235(.A(new_n435_), .B(new_n436_), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n432_), .B(new_n437_), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n438_), .B(new_n379_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(G15gat), .B(G43gat), .ZN(new_n440_));
  XNOR2_X1  g239(.A(new_n440_), .B(KEYINPUT87), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n441_), .B(KEYINPUT30), .ZN(new_n442_));
  XNOR2_X1  g241(.A(new_n442_), .B(KEYINPUT31), .ZN(new_n443_));
  INV_X1    g242(.A(new_n443_), .ZN(new_n444_));
  OR2_X1    g243(.A1(new_n439_), .A2(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n439_), .A2(new_n444_), .ZN(new_n446_));
  AOI21_X1  g245(.A(new_n403_), .B1(new_n445_), .B2(new_n446_), .ZN(new_n447_));
  INV_X1    g246(.A(KEYINPUT29), .ZN(new_n448_));
  INV_X1    g247(.A(G228gat), .ZN(new_n449_));
  INV_X1    g248(.A(G233gat), .ZN(new_n450_));
  NOR2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  INV_X1    g250(.A(new_n451_), .ZN(new_n452_));
  OAI22_X1  g251(.A1(new_n381_), .A2(new_n448_), .B1(KEYINPUT91), .B2(new_n452_), .ZN(new_n453_));
  INV_X1    g252(.A(KEYINPUT90), .ZN(new_n454_));
  XOR2_X1   g253(.A(G197gat), .B(G204gat), .Z(new_n455_));
  NAND2_X1  g254(.A1(new_n455_), .A2(KEYINPUT21), .ZN(new_n456_));
  XNOR2_X1  g255(.A(G211gat), .B(G218gat), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n454_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  INV_X1    g257(.A(new_n457_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n459_), .A2(new_n455_), .A3(KEYINPUT90), .A4(KEYINPUT21), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n459_), .B1(KEYINPUT21), .B2(new_n455_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n455_), .A2(KEYINPUT21), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n461_), .A2(new_n464_), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  OAI21_X1  g265(.A(G78gat), .B1(new_n453_), .B2(new_n466_), .ZN(new_n467_));
  INV_X1    g266(.A(KEYINPUT91), .ZN(new_n468_));
  AOI22_X1  g267(.A1(new_n376_), .A2(KEYINPUT29), .B1(new_n468_), .B2(new_n451_), .ZN(new_n469_));
  INV_X1    g268(.A(G78gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n469_), .A2(new_n470_), .A3(new_n465_), .ZN(new_n471_));
  AOI21_X1  g270(.A(G106gat), .B1(new_n467_), .B2(new_n471_), .ZN(new_n472_));
  INV_X1    g271(.A(new_n472_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n467_), .A2(new_n471_), .A3(G106gat), .ZN(new_n474_));
  XNOR2_X1  g273(.A(G22gat), .B(G50gat), .ZN(new_n475_));
  INV_X1    g274(.A(new_n475_), .ZN(new_n476_));
  NAND3_X1  g275(.A1(new_n473_), .A2(new_n474_), .A3(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(new_n474_), .ZN(new_n478_));
  OAI21_X1  g277(.A(new_n475_), .B1(new_n478_), .B2(new_n472_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n477_), .A2(new_n479_), .ZN(new_n480_));
  OAI21_X1  g279(.A(KEYINPUT28), .B1(new_n376_), .B2(KEYINPUT29), .ZN(new_n481_));
  OR3_X1    g280(.A1(new_n376_), .A2(KEYINPUT28), .A3(KEYINPUT29), .ZN(new_n482_));
  NOR2_X1   g281(.A1(new_n451_), .A2(new_n468_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  AND3_X1   g283(.A1(new_n481_), .A2(new_n482_), .A3(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n484_), .B1(new_n482_), .B2(new_n481_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  INV_X1    g286(.A(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n480_), .A2(new_n488_), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n477_), .A2(new_n479_), .A3(new_n487_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n489_), .A2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(G226gat), .A2(G233gat), .ZN(new_n492_));
  XNOR2_X1  g291(.A(new_n492_), .B(KEYINPUT19), .ZN(new_n493_));
  INV_X1    g292(.A(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT20), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n408_), .B(KEYINPUT92), .ZN(new_n496_));
  INV_X1    g295(.A(G176gat), .ZN(new_n497_));
  AOI21_X1  g296(.A(new_n496_), .B1(new_n497_), .B2(new_n413_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n498_), .A2(new_n407_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n431_), .A2(new_n499_), .ZN(new_n500_));
  AOI21_X1  g299(.A(new_n495_), .B1(new_n500_), .B2(new_n465_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n418_), .A2(new_n466_), .A3(new_n431_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n494_), .B1(new_n501_), .B2(new_n502_), .ZN(new_n503_));
  AOI21_X1  g302(.A(new_n429_), .B1(new_n422_), .B2(new_n423_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n504_), .B1(new_n407_), .B2(new_n498_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n505_), .A2(KEYINPUT93), .A3(new_n466_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT93), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n507_), .B1(new_n500_), .B2(new_n465_), .ZN(new_n508_));
  NAND2_X1  g307(.A1(new_n506_), .A2(new_n508_), .ZN(new_n509_));
  OAI21_X1  g308(.A(new_n465_), .B1(new_n417_), .B2(new_n504_), .ZN(new_n510_));
  AND3_X1   g309(.A1(new_n510_), .A2(KEYINPUT20), .A3(new_n494_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n503_), .B1(new_n509_), .B2(new_n511_), .ZN(new_n512_));
  XNOR2_X1  g311(.A(G8gat), .B(G36gat), .ZN(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT18), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G64gat), .B(G92gat), .ZN(new_n515_));
  XOR2_X1   g314(.A(new_n514_), .B(new_n515_), .Z(new_n516_));
  NAND2_X1  g315(.A1(new_n512_), .A2(new_n516_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n516_), .ZN(new_n518_));
  AND2_X1   g317(.A1(new_n509_), .A2(new_n511_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n518_), .B1(new_n519_), .B2(new_n503_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT27), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n522_), .B1(new_n512_), .B2(new_n516_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT96), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n465_), .B1(new_n500_), .B2(new_n524_), .ZN(new_n525_));
  NAND2_X1  g324(.A1(new_n505_), .A2(KEYINPUT96), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  XNOR2_X1  g326(.A(KEYINPUT95), .B(KEYINPUT20), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n510_), .A2(new_n528_), .ZN(new_n529_));
  AOI21_X1  g328(.A(new_n494_), .B1(new_n527_), .B2(new_n529_), .ZN(new_n530_));
  AND3_X1   g329(.A1(new_n501_), .A2(new_n502_), .A3(new_n494_), .ZN(new_n531_));
  OAI21_X1  g330(.A(new_n518_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n532_));
  AOI22_X1  g331(.A1(new_n521_), .A2(new_n522_), .B1(new_n523_), .B2(new_n532_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n491_), .A2(new_n533_), .A3(KEYINPUT99), .ZN(new_n534_));
  AOI21_X1  g333(.A(KEYINPUT99), .B1(new_n491_), .B2(new_n533_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n447_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND2_X1  g335(.A1(new_n516_), .A2(KEYINPUT32), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n538_), .B1(new_n530_), .B2(new_n531_), .ZN(new_n539_));
  INV_X1    g338(.A(KEYINPUT97), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n539_), .A2(new_n540_), .ZN(new_n541_));
  OAI211_X1 g340(.A(KEYINPUT97), .B(new_n538_), .C1(new_n530_), .C2(new_n531_), .ZN(new_n542_));
  NAND2_X1  g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n512_), .A2(new_n537_), .ZN(new_n544_));
  NAND3_X1  g343(.A1(new_n403_), .A2(new_n543_), .A3(new_n544_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n394_), .A2(new_n385_), .ZN(new_n546_));
  OAI211_X1 g345(.A(new_n546_), .B(new_n391_), .C1(new_n385_), .C2(new_n384_), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n517_), .A2(new_n520_), .A3(new_n547_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT33), .ZN(new_n549_));
  XNOR2_X1  g348(.A(new_n398_), .B(new_n549_), .ZN(new_n550_));
  OAI21_X1  g349(.A(KEYINPUT94), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  NOR3_X1   g350(.A1(new_n519_), .A2(new_n518_), .A3(new_n503_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n503_), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n509_), .A2(new_n511_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n516_), .B1(new_n553_), .B2(new_n554_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n552_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(new_n398_), .B(KEYINPUT33), .ZN(new_n557_));
  INV_X1    g356(.A(KEYINPUT94), .ZN(new_n558_));
  NAND4_X1  g357(.A1(new_n556_), .A2(new_n557_), .A3(new_n558_), .A4(new_n547_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n545_), .A2(new_n551_), .A3(new_n559_), .ZN(new_n560_));
  NAND3_X1  g359(.A1(new_n489_), .A2(new_n402_), .A3(new_n490_), .ZN(new_n561_));
  INV_X1    g360(.A(new_n561_), .ZN(new_n562_));
  AOI22_X1  g361(.A1(new_n560_), .A2(new_n491_), .B1(new_n562_), .B2(new_n533_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n445_), .A2(new_n446_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n536_), .B1(new_n563_), .B2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n251_), .A2(new_n253_), .A3(new_n307_), .ZN(new_n566_));
  XNOR2_X1  g365(.A(new_n566_), .B(KEYINPUT83), .ZN(new_n567_));
  OR2_X1    g366(.A1(new_n307_), .A2(new_n248_), .ZN(new_n568_));
  XNOR2_X1  g367(.A(new_n568_), .B(KEYINPUT82), .ZN(new_n569_));
  NAND2_X1  g368(.A1(G229gat), .A2(G233gat), .ZN(new_n570_));
  AND2_X1   g369(.A1(new_n569_), .A2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(new_n307_), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n569_), .B1(new_n572_), .B2(new_n249_), .ZN(new_n573_));
  INV_X1    g372(.A(new_n570_), .ZN(new_n574_));
  AOI22_X1  g373(.A1(new_n567_), .A2(new_n571_), .B1(new_n573_), .B2(new_n574_), .ZN(new_n575_));
  XNOR2_X1  g374(.A(G113gat), .B(G141gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(G169gat), .B(G197gat), .ZN(new_n577_));
  XOR2_X1   g376(.A(new_n576_), .B(new_n577_), .Z(new_n578_));
  XNOR2_X1  g377(.A(new_n575_), .B(new_n578_), .ZN(new_n579_));
  AND2_X1   g378(.A1(new_n565_), .A2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n353_), .A2(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n324_), .B1(new_n323_), .B2(new_n352_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n202_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n582_), .ZN(new_n584_));
  NAND4_X1  g383(.A1(new_n584_), .A2(KEYINPUT100), .A3(new_n353_), .A4(new_n580_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n583_), .A2(new_n585_), .ZN(new_n586_));
  NOR3_X1   g385(.A1(new_n586_), .A2(G1gat), .A3(new_n402_), .ZN(new_n587_));
  XOR2_X1   g386(.A(KEYINPUT101), .B(KEYINPUT38), .Z(new_n588_));
  OR2_X1    g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n579_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n351_), .A2(new_n590_), .ZN(new_n591_));
  NAND2_X1  g390(.A1(new_n591_), .A2(new_n320_), .ZN(new_n592_));
  INV_X1    g391(.A(KEYINPUT102), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n592_), .A2(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n285_), .A2(new_n277_), .ZN(new_n595_));
  AND2_X1   g394(.A1(new_n565_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n591_), .A2(KEYINPUT102), .A3(new_n320_), .ZN(new_n597_));
  AND3_X1   g396(.A1(new_n594_), .A2(new_n596_), .A3(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  OAI21_X1  g398(.A(G1gat), .B1(new_n599_), .B2(new_n402_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n587_), .A2(new_n588_), .ZN(new_n601_));
  NAND3_X1  g400(.A1(new_n589_), .A2(new_n600_), .A3(new_n601_), .ZN(G1324gat));
  NOR2_X1   g401(.A1(new_n533_), .A2(new_n302_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n583_), .A2(new_n585_), .A3(new_n603_), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n604_), .B(KEYINPUT103), .ZN(new_n605_));
  INV_X1    g404(.A(new_n533_), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n598_), .A2(new_n606_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n607_), .A2(G8gat), .ZN(new_n608_));
  NAND2_X1  g407(.A1(new_n608_), .A2(KEYINPUT39), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT39), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n607_), .A2(new_n610_), .A3(G8gat), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n609_), .A2(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n605_), .A2(new_n612_), .ZN(new_n613_));
  INV_X1    g412(.A(KEYINPUT40), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n605_), .A2(new_n612_), .A3(KEYINPUT40), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(G1325gat));
  INV_X1    g416(.A(G15gat), .ZN(new_n618_));
  AOI21_X1  g417(.A(new_n618_), .B1(new_n598_), .B2(new_n564_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT41), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  NAND4_X1  g420(.A1(new_n583_), .A2(new_n585_), .A3(new_n618_), .A4(new_n564_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n619_), .A2(new_n620_), .ZN(new_n623_));
  NAND3_X1  g422(.A1(new_n621_), .A2(new_n622_), .A3(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT104), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(G1326gat));
  OAI21_X1  g425(.A(G22gat), .B1(new_n599_), .B2(new_n491_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT42), .ZN(new_n628_));
  OR2_X1    g427(.A1(new_n491_), .A2(G22gat), .ZN(new_n629_));
  OAI21_X1  g428(.A(new_n628_), .B1(new_n586_), .B2(new_n629_), .ZN(G1327gat));
  NOR2_X1   g429(.A1(new_n321_), .A2(new_n595_), .ZN(new_n631_));
  NAND3_X1  g430(.A1(new_n591_), .A2(new_n565_), .A3(new_n631_), .ZN(new_n632_));
  XOR2_X1   g431(.A(new_n632_), .B(KEYINPUT107), .Z(new_n633_));
  AOI21_X1  g432(.A(G29gat), .B1(new_n633_), .B2(new_n403_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n565_), .A2(new_n291_), .ZN(new_n635_));
  NAND2_X1  g434(.A1(new_n283_), .A2(new_n287_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n289_), .A2(new_n290_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OAI21_X1  g437(.A(KEYINPUT43), .B1(new_n638_), .B2(KEYINPUT105), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n321_), .B1(new_n635_), .B2(new_n639_), .ZN(new_n640_));
  NAND4_X1  g439(.A1(new_n565_), .A2(new_n291_), .A3(KEYINPUT105), .A4(KEYINPUT43), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n640_), .A2(new_n591_), .A3(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT44), .ZN(new_n643_));
  AND2_X1   g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  AND2_X1   g443(.A1(new_n640_), .A2(new_n641_), .ZN(new_n645_));
  INV_X1    g444(.A(KEYINPUT106), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n645_), .A2(new_n646_), .A3(KEYINPUT44), .A4(new_n591_), .ZN(new_n647_));
  OAI21_X1  g446(.A(KEYINPUT106), .B1(new_n642_), .B2(new_n643_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n644_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n403_), .A2(G29gat), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n634_), .B1(new_n649_), .B2(new_n650_), .ZN(G1328gat));
  INV_X1    g450(.A(KEYINPUT46), .ZN(new_n652_));
  INV_X1    g451(.A(G36gat), .ZN(new_n653_));
  AOI21_X1  g452(.A(new_n653_), .B1(new_n649_), .B2(new_n606_), .ZN(new_n654_));
  NAND3_X1  g453(.A1(new_n633_), .A2(new_n653_), .A3(new_n606_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT45), .ZN(new_n656_));
  XNOR2_X1  g455(.A(new_n655_), .B(new_n656_), .ZN(new_n657_));
  OAI21_X1  g456(.A(new_n652_), .B1(new_n654_), .B2(new_n657_), .ZN(new_n658_));
  XNOR2_X1  g457(.A(new_n655_), .B(KEYINPUT45), .ZN(new_n659_));
  AOI211_X1 g458(.A(new_n533_), .B(new_n644_), .C1(new_n647_), .C2(new_n648_), .ZN(new_n660_));
  OAI211_X1 g459(.A(new_n659_), .B(KEYINPUT46), .C1(new_n660_), .C2(new_n653_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n658_), .A2(new_n661_), .ZN(G1329gat));
  AOI21_X1  g461(.A(G43gat), .B1(new_n633_), .B2(new_n564_), .ZN(new_n663_));
  AND2_X1   g462(.A1(new_n564_), .A2(G43gat), .ZN(new_n664_));
  AOI21_X1  g463(.A(new_n663_), .B1(new_n649_), .B2(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT47), .ZN(new_n666_));
  XNOR2_X1  g465(.A(new_n665_), .B(new_n666_), .ZN(G1330gat));
  INV_X1    g466(.A(G50gat), .ZN(new_n668_));
  INV_X1    g467(.A(new_n491_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n633_), .A2(new_n668_), .A3(new_n669_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT108), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n649_), .A2(new_n669_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n671_), .B1(new_n672_), .B2(G50gat), .ZN(new_n673_));
  AOI211_X1 g472(.A(KEYINPUT108), .B(new_n668_), .C1(new_n649_), .C2(new_n669_), .ZN(new_n674_));
  OAI21_X1  g473(.A(new_n670_), .B1(new_n673_), .B2(new_n674_), .ZN(G1331gat));
  NOR2_X1   g474(.A1(new_n352_), .A2(new_n579_), .ZN(new_n676_));
  AND2_X1   g475(.A1(new_n676_), .A2(new_n565_), .ZN(new_n677_));
  AND2_X1   g476(.A1(new_n677_), .A2(new_n323_), .ZN(new_n678_));
  INV_X1    g477(.A(G57gat), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n678_), .A2(new_n679_), .A3(new_n403_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n596_), .A2(new_n676_), .A3(new_n321_), .ZN(new_n681_));
  OAI21_X1  g480(.A(G57gat), .B1(new_n681_), .B2(new_n402_), .ZN(new_n682_));
  NAND2_X1  g481(.A1(new_n680_), .A2(new_n682_), .ZN(G1332gat));
  OAI21_X1  g482(.A(G64gat), .B1(new_n681_), .B2(new_n533_), .ZN(new_n684_));
  XOR2_X1   g483(.A(KEYINPUT109), .B(KEYINPUT48), .Z(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(new_n686_));
  INV_X1    g485(.A(G64gat), .ZN(new_n687_));
  NAND3_X1  g486(.A1(new_n678_), .A2(new_n687_), .A3(new_n606_), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n686_), .A2(new_n688_), .ZN(G1333gat));
  INV_X1    g488(.A(new_n564_), .ZN(new_n690_));
  OAI21_X1  g489(.A(G71gat), .B1(new_n681_), .B2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(new_n691_), .B(KEYINPUT49), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n678_), .A2(new_n434_), .A3(new_n564_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n692_), .A2(new_n693_), .ZN(G1334gat));
  OAI21_X1  g493(.A(G78gat), .B1(new_n681_), .B2(new_n491_), .ZN(new_n695_));
  XNOR2_X1  g494(.A(new_n695_), .B(KEYINPUT50), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n678_), .A2(new_n470_), .A3(new_n669_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1335gat));
  NAND2_X1  g497(.A1(new_n635_), .A2(new_n639_), .ZN(new_n699_));
  NAND4_X1  g498(.A1(new_n699_), .A2(new_n322_), .A3(new_n641_), .A4(new_n676_), .ZN(new_n700_));
  NAND2_X1  g499(.A1(new_n700_), .A2(KEYINPUT110), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT110), .ZN(new_n702_));
  NAND4_X1  g501(.A1(new_n640_), .A2(new_n702_), .A3(new_n641_), .A4(new_n676_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n701_), .A2(new_n703_), .ZN(new_n704_));
  OAI21_X1  g503(.A(G85gat), .B1(new_n704_), .B2(new_n402_), .ZN(new_n705_));
  AND2_X1   g504(.A1(new_n677_), .A2(new_n631_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(new_n241_), .A3(new_n403_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(G1336gat));
  OAI21_X1  g507(.A(G92gat), .B1(new_n704_), .B2(new_n533_), .ZN(new_n709_));
  NAND3_X1  g508(.A1(new_n706_), .A2(new_n242_), .A3(new_n606_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n709_), .A2(new_n710_), .ZN(G1337gat));
  INV_X1    g510(.A(KEYINPUT51), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n706_), .A2(new_n238_), .A3(new_n564_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n690_), .B1(new_n701_), .B2(new_n703_), .ZN(new_n714_));
  OAI211_X1 g513(.A(new_n712_), .B(new_n713_), .C1(new_n714_), .C2(new_n436_), .ZN(new_n715_));
  AND2_X1   g514(.A1(new_n715_), .A2(KEYINPUT112), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n715_), .A2(KEYINPUT112), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n713_), .B1(new_n714_), .B2(new_n436_), .ZN(new_n718_));
  AND3_X1   g517(.A1(new_n718_), .A2(KEYINPUT111), .A3(KEYINPUT51), .ZN(new_n719_));
  AOI21_X1  g518(.A(KEYINPUT111), .B1(new_n718_), .B2(KEYINPUT51), .ZN(new_n720_));
  OAI22_X1  g519(.A1(new_n716_), .A2(new_n717_), .B1(new_n719_), .B2(new_n720_), .ZN(G1338gat));
  NAND3_X1  g520(.A1(new_n706_), .A2(new_n239_), .A3(new_n669_), .ZN(new_n722_));
  OR2_X1    g521(.A1(new_n700_), .A2(new_n491_), .ZN(new_n723_));
  INV_X1    g522(.A(KEYINPUT52), .ZN(new_n724_));
  AND3_X1   g523(.A1(new_n723_), .A2(new_n724_), .A3(G106gat), .ZN(new_n725_));
  AOI21_X1  g524(.A(new_n724_), .B1(new_n723_), .B2(G106gat), .ZN(new_n726_));
  OAI21_X1  g525(.A(new_n722_), .B1(new_n725_), .B2(new_n726_), .ZN(new_n727_));
  XNOR2_X1  g526(.A(new_n727_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g527(.A1(new_n323_), .A2(new_n352_), .A3(new_n590_), .ZN(new_n729_));
  XNOR2_X1  g528(.A(new_n729_), .B(KEYINPUT54), .ZN(new_n730_));
  INV_X1    g529(.A(KEYINPUT113), .ZN(new_n731_));
  INV_X1    g530(.A(KEYINPUT55), .ZN(new_n732_));
  OAI21_X1  g531(.A(new_n325_), .B1(new_n336_), .B2(new_n335_), .ZN(new_n733_));
  AOI22_X1  g532(.A1(new_n337_), .A2(new_n732_), .B1(new_n340_), .B2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n338_), .A2(KEYINPUT12), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n266_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n735_), .A2(new_n736_), .ZN(new_n737_));
  NAND4_X1  g536(.A1(new_n737_), .A2(KEYINPUT55), .A3(new_n330_), .A4(new_n332_), .ZN(new_n738_));
  AOI21_X1  g537(.A(new_n347_), .B1(new_n734_), .B2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(new_n731_), .B1(new_n739_), .B2(KEYINPUT56), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n332_), .B1(new_n336_), .B2(new_n335_), .ZN(new_n741_));
  AOI21_X1  g540(.A(new_n331_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n742_));
  OAI21_X1  g541(.A(new_n732_), .B1(new_n741_), .B2(new_n742_), .ZN(new_n743_));
  NAND2_X1  g542(.A1(new_n733_), .A2(new_n340_), .ZN(new_n744_));
  NAND3_X1  g543(.A1(new_n743_), .A2(new_n738_), .A3(new_n744_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n745_), .A2(new_n346_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT56), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n746_), .A2(KEYINPUT113), .A3(new_n747_), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n745_), .A2(KEYINPUT56), .A3(new_n346_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT114), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND4_X1  g550(.A1(new_n745_), .A2(KEYINPUT114), .A3(KEYINPUT56), .A4(new_n346_), .ZN(new_n752_));
  NAND4_X1  g551(.A1(new_n740_), .A2(new_n748_), .A3(new_n751_), .A4(new_n752_), .ZN(new_n753_));
  NAND3_X1  g552(.A1(new_n337_), .A2(new_n341_), .A3(new_n347_), .ZN(new_n754_));
  AND2_X1   g553(.A1(new_n579_), .A2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n753_), .A2(new_n755_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n575_), .A2(new_n578_), .ZN(new_n757_));
  AOI21_X1  g556(.A(new_n578_), .B1(new_n573_), .B2(new_n570_), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n567_), .A2(new_n569_), .A3(new_n574_), .ZN(new_n759_));
  NAND2_X1  g558(.A1(new_n758_), .A2(new_n759_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n757_), .A2(new_n760_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n348_), .A2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n756_), .A2(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(KEYINPUT57), .B1(new_n764_), .B2(new_n595_), .ZN(new_n765_));
  AND3_X1   g564(.A1(new_n757_), .A2(new_n754_), .A3(new_n760_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n749_), .ZN(new_n767_));
  AOI21_X1  g566(.A(KEYINPUT56), .B1(new_n745_), .B2(new_n346_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n766_), .B1(new_n767_), .B2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT58), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n769_), .A2(new_n770_), .ZN(new_n771_));
  OAI211_X1 g570(.A(new_n766_), .B(KEYINPUT58), .C1(new_n767_), .C2(new_n768_), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n771_), .A2(new_n291_), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n762_), .B1(new_n753_), .B2(new_n755_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n595_), .A2(KEYINPUT57), .ZN(new_n775_));
  OAI21_X1  g574(.A(new_n773_), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(new_n322_), .B1(new_n765_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n730_), .A2(new_n777_), .ZN(new_n778_));
  OAI211_X1 g577(.A(new_n403_), .B(new_n564_), .C1(new_n534_), .C2(new_n535_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n779_), .A2(KEYINPUT59), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n778_), .A2(new_n780_), .ZN(new_n781_));
  OAI21_X1  g580(.A(KEYINPUT115), .B1(new_n765_), .B2(new_n776_), .ZN(new_n782_));
  INV_X1    g581(.A(new_n320_), .ZN(new_n783_));
  OR2_X1    g582(.A1(new_n774_), .A2(new_n775_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT57), .ZN(new_n785_));
  INV_X1    g584(.A(new_n595_), .ZN(new_n786_));
  OAI21_X1  g585(.A(new_n785_), .B1(new_n774_), .B2(new_n786_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788_));
  NAND4_X1  g587(.A1(new_n784_), .A2(new_n787_), .A3(new_n788_), .A4(new_n773_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n782_), .A2(new_n783_), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n779_), .B1(new_n790_), .B2(new_n730_), .ZN(new_n791_));
  INV_X1    g590(.A(KEYINPUT59), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n781_), .B1(new_n791_), .B2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(G113gat), .B1(new_n793_), .B2(new_n590_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n790_), .A2(new_n730_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n779_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  OR2_X1    g596(.A1(new_n590_), .A2(G113gat), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n794_), .B1(new_n797_), .B2(new_n798_), .ZN(G1340gat));
  XNOR2_X1  g598(.A(KEYINPUT116), .B(G120gat), .ZN(new_n800_));
  AOI21_X1  g599(.A(KEYINPUT60), .B1(new_n351_), .B2(new_n800_), .ZN(new_n801_));
  OR3_X1    g600(.A1(new_n797_), .A2(KEYINPUT60), .A3(new_n801_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n351_), .B1(new_n797_), .B2(new_n801_), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n803_), .A2(new_n793_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n802_), .B1(new_n804_), .B2(new_n800_), .ZN(G1341gat));
  AOI21_X1  g604(.A(G127gat), .B1(new_n791_), .B2(new_n321_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n793_), .ZN(new_n807_));
  XNOR2_X1  g606(.A(KEYINPUT117), .B(G127gat), .ZN(new_n808_));
  NOR2_X1   g607(.A1(new_n783_), .A2(new_n808_), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n806_), .B1(new_n807_), .B2(new_n809_), .ZN(G1342gat));
  NAND3_X1  g609(.A1(new_n795_), .A2(new_n786_), .A3(new_n796_), .ZN(new_n811_));
  INV_X1    g610(.A(G134gat), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n811_), .A2(new_n812_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n291_), .A2(G134gat), .ZN(new_n814_));
  XNOR2_X1  g613(.A(new_n814_), .B(KEYINPUT118), .ZN(new_n815_));
  OAI211_X1 g614(.A(new_n781_), .B(new_n815_), .C1(new_n791_), .C2(new_n792_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n813_), .A2(new_n816_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n817_), .A2(KEYINPUT119), .ZN(new_n818_));
  INV_X1    g617(.A(KEYINPUT119), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n813_), .A2(new_n816_), .A3(new_n819_), .ZN(new_n820_));
  NAND2_X1  g619(.A1(new_n818_), .A2(new_n820_), .ZN(G1343gat));
  NOR4_X1   g620(.A1(new_n606_), .A2(new_n564_), .A3(new_n491_), .A4(new_n402_), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n822_), .B(KEYINPUT120), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n795_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n825_), .A2(new_n579_), .ZN(new_n826_));
  XNOR2_X1  g625(.A(new_n826_), .B(G141gat), .ZN(G1344gat));
  NOR2_X1   g626(.A1(new_n824_), .A2(new_n352_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(KEYINPUT121), .B(G148gat), .ZN(new_n829_));
  XNOR2_X1  g628(.A(new_n828_), .B(new_n829_), .ZN(G1345gat));
  NOR2_X1   g629(.A1(new_n824_), .A2(new_n322_), .ZN(new_n831_));
  XOR2_X1   g630(.A(KEYINPUT61), .B(G155gat), .Z(new_n832_));
  XNOR2_X1  g631(.A(new_n831_), .B(new_n832_), .ZN(G1346gat));
  OAI21_X1  g632(.A(G162gat), .B1(new_n824_), .B2(new_n638_), .ZN(new_n834_));
  NAND2_X1  g633(.A1(new_n786_), .A2(new_n357_), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n834_), .B1(new_n824_), .B2(new_n835_), .ZN(G1347gat));
  INV_X1    g635(.A(KEYINPUT62), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n447_), .A2(new_n606_), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n838_), .A2(new_n669_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(new_n840_), .B1(new_n730_), .B2(new_n777_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n841_), .ZN(new_n842_));
  NOR2_X1   g641(.A1(new_n842_), .A2(new_n590_), .ZN(new_n843_));
  INV_X1    g642(.A(G169gat), .ZN(new_n844_));
  OAI21_X1  g643(.A(new_n837_), .B1(new_n843_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n843_), .A2(new_n413_), .ZN(new_n846_));
  OAI211_X1 g645(.A(KEYINPUT62), .B(G169gat), .C1(new_n842_), .C2(new_n590_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n845_), .A2(new_n846_), .A3(new_n847_), .ZN(G1348gat));
  AOI21_X1  g647(.A(G176gat), .B1(new_n841_), .B2(new_n351_), .ZN(new_n849_));
  AOI21_X1  g648(.A(new_n669_), .B1(new_n790_), .B2(new_n730_), .ZN(new_n850_));
  NOR3_X1   g649(.A1(new_n352_), .A2(new_n497_), .A3(new_n838_), .ZN(new_n851_));
  AOI21_X1  g650(.A(new_n849_), .B1(new_n850_), .B2(new_n851_), .ZN(G1349gat));
  NOR2_X1   g651(.A1(new_n783_), .A2(new_n425_), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n841_), .A2(new_n853_), .ZN(new_n854_));
  INV_X1    g653(.A(KEYINPUT122), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n322_), .A2(new_n838_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n850_), .A2(new_n857_), .ZN(new_n858_));
  INV_X1    g657(.A(new_n858_), .ZN(new_n859_));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860_));
  AOI21_X1  g659(.A(G183gat), .B1(new_n859_), .B2(new_n860_), .ZN(new_n861_));
  NAND2_X1  g660(.A1(new_n858_), .A2(KEYINPUT123), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n856_), .B1(new_n861_), .B2(new_n862_), .ZN(G1350gat));
  AND3_X1   g662(.A1(new_n841_), .A2(new_n786_), .A3(new_n426_), .ZN(new_n864_));
  INV_X1    g663(.A(G190gat), .ZN(new_n865_));
  AOI21_X1  g664(.A(new_n865_), .B1(new_n841_), .B2(new_n291_), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT124), .ZN(new_n867_));
  OR3_X1    g666(.A1(new_n864_), .A2(new_n866_), .A3(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(G1351gat));
  INV_X1    g669(.A(G197gat), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n561_), .A2(new_n564_), .A3(new_n533_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n795_), .A2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n871_), .B1(new_n873_), .B2(new_n590_), .ZN(new_n874_));
  INV_X1    g673(.A(KEYINPUT126), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  OAI211_X1 g675(.A(KEYINPUT126), .B(new_n871_), .C1(new_n873_), .C2(new_n590_), .ZN(new_n877_));
  NAND4_X1  g676(.A1(new_n795_), .A2(G197gat), .A3(new_n579_), .A4(new_n872_), .ZN(new_n878_));
  INV_X1    g677(.A(KEYINPUT125), .ZN(new_n879_));
  OR2_X1    g678(.A1(new_n878_), .A2(new_n879_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n878_), .A2(new_n879_), .ZN(new_n881_));
  AOI22_X1  g680(.A1(new_n876_), .A2(new_n877_), .B1(new_n880_), .B2(new_n881_), .ZN(G1352gat));
  INV_X1    g681(.A(new_n873_), .ZN(new_n883_));
  NAND2_X1  g682(.A1(new_n883_), .A2(new_n351_), .ZN(new_n884_));
  XNOR2_X1  g683(.A(new_n884_), .B(G204gat), .ZN(G1353gat));
  INV_X1    g684(.A(KEYINPUT63), .ZN(new_n886_));
  INV_X1    g685(.A(G211gat), .ZN(new_n887_));
  OAI21_X1  g686(.A(new_n320_), .B1(new_n886_), .B2(new_n887_), .ZN(new_n888_));
  XOR2_X1   g687(.A(new_n888_), .B(KEYINPUT127), .Z(new_n889_));
  NAND2_X1  g688(.A1(new_n883_), .A2(new_n889_), .ZN(new_n890_));
  NAND2_X1  g689(.A1(new_n886_), .A2(new_n887_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n890_), .B(new_n891_), .ZN(G1354gat));
  OR3_X1    g691(.A1(new_n873_), .A2(G218gat), .A3(new_n595_), .ZN(new_n893_));
  OAI21_X1  g692(.A(G218gat), .B1(new_n873_), .B2(new_n638_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n893_), .A2(new_n894_), .ZN(G1355gat));
endmodule


