//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n760_, new_n761_,
    new_n762_, new_n763_, new_n764_, new_n765_, new_n766_, new_n767_,
    new_n768_, new_n769_, new_n770_, new_n771_, new_n772_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n812_, new_n813_, new_n815_,
    new_n816_, new_n817_, new_n818_, new_n819_, new_n820_, new_n821_,
    new_n823_, new_n824_, new_n825_, new_n826_, new_n827_, new_n828_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n929_, new_n930_, new_n932_, new_n933_, new_n934_, new_n935_,
    new_n937_, new_n939_, new_n940_, new_n941_, new_n943_, new_n944_,
    new_n945_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n966_, new_n967_, new_n968_, new_n970_, new_n971_, new_n973_,
    new_n974_, new_n976_, new_n977_, new_n979_, new_n980_, new_n981_,
    new_n983_, new_n984_, new_n985_;
  INV_X1    g000(.A(KEYINPUT76), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203_));
  INV_X1    g002(.A(G1gat), .ZN(new_n204_));
  INV_X1    g003(.A(G8gat), .ZN(new_n205_));
  OAI21_X1  g004(.A(KEYINPUT14), .B1(new_n204_), .B2(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(new_n203_), .A2(new_n206_), .ZN(new_n207_));
  XNOR2_X1  g006(.A(G1gat), .B(G8gat), .ZN(new_n208_));
  OR2_X1    g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n207_), .A2(new_n208_), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  XNOR2_X1  g010(.A(G29gat), .B(G36gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G43gat), .B(G50gat), .ZN(new_n213_));
  OR2_X1    g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n213_), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n211_), .A2(new_n217_), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n216_), .A2(new_n209_), .A3(new_n210_), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n218_), .A2(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(G229gat), .A2(G233gat), .ZN(new_n221_));
  INV_X1    g020(.A(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(new_n220_), .A2(new_n222_), .ZN(new_n223_));
  INV_X1    g022(.A(KEYINPUT15), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n216_), .A2(new_n224_), .ZN(new_n225_));
  NAND3_X1  g024(.A1(new_n214_), .A2(KEYINPUT15), .A3(new_n215_), .ZN(new_n226_));
  NAND3_X1  g025(.A1(new_n225_), .A2(new_n211_), .A3(new_n226_), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n227_), .A2(new_n219_), .A3(new_n221_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G113gat), .B(G141gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G169gat), .ZN(new_n230_));
  XOR2_X1   g029(.A(new_n230_), .B(G197gat), .Z(new_n231_));
  AND3_X1   g030(.A1(new_n223_), .A2(new_n228_), .A3(new_n231_), .ZN(new_n232_));
  AOI21_X1  g031(.A(new_n231_), .B1(new_n223_), .B2(new_n228_), .ZN(new_n233_));
  OAI21_X1  g032(.A(new_n202_), .B1(new_n232_), .B2(new_n233_), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n223_), .A2(new_n228_), .ZN(new_n235_));
  INV_X1    g034(.A(new_n231_), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n235_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n223_), .A2(new_n228_), .A3(new_n231_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n237_), .A2(KEYINPUT76), .A3(new_n238_), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n234_), .A2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n241_));
  OR2_X1    g040(.A1(KEYINPUT72), .A2(KEYINPUT13), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G71gat), .B(G78gat), .ZN(new_n243_));
  XOR2_X1   g042(.A(G57gat), .B(G64gat), .Z(new_n244_));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n245_));
  AOI21_X1  g044(.A(new_n243_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  XOR2_X1   g047(.A(G71gat), .B(G78gat), .Z(new_n249_));
  XNOR2_X1  g048(.A(G57gat), .B(G64gat), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n249_), .B1(KEYINPUT11), .B2(new_n250_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT69), .ZN(new_n252_));
  NOR2_X1   g051(.A1(new_n244_), .A2(new_n245_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n248_), .A2(new_n252_), .A3(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  AOI21_X1  g054(.A(new_n253_), .B1(new_n248_), .B2(new_n252_), .ZN(new_n256_));
  NOR2_X1   g055(.A1(new_n255_), .A2(new_n256_), .ZN(new_n257_));
  INV_X1    g056(.A(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT68), .ZN(new_n259_));
  INV_X1    g058(.A(KEYINPUT7), .ZN(new_n260_));
  INV_X1    g059(.A(G99gat), .ZN(new_n261_));
  INV_X1    g060(.A(G106gat), .ZN(new_n262_));
  NAND4_X1  g061(.A1(new_n260_), .A2(new_n261_), .A3(new_n262_), .A4(KEYINPUT67), .ZN(new_n263_));
  OAI211_X1 g062(.A(new_n261_), .B(new_n262_), .C1(new_n260_), .C2(KEYINPUT67), .ZN(new_n264_));
  NAND2_X1  g063(.A1(new_n260_), .A2(KEYINPUT67), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT6), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(KEYINPUT66), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(KEYINPUT6), .ZN(new_n270_));
  NAND2_X1  g069(.A1(G99gat), .A2(G106gat), .ZN(new_n271_));
  AND3_X1   g070(.A1(new_n268_), .A2(new_n270_), .A3(new_n271_), .ZN(new_n272_));
  AOI21_X1  g071(.A(new_n271_), .B1(new_n268_), .B2(new_n270_), .ZN(new_n273_));
  OAI211_X1 g072(.A(new_n263_), .B(new_n266_), .C1(new_n272_), .C2(new_n273_), .ZN(new_n274_));
  XOR2_X1   g073(.A(G85gat), .B(G92gat), .Z(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n276_), .A2(KEYINPUT8), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT8), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n274_), .A2(new_n278_), .A3(new_n275_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  XOR2_X1   g079(.A(KEYINPUT65), .B(KEYINPUT9), .Z(new_n281_));
  INV_X1    g080(.A(G85gat), .ZN(new_n282_));
  INV_X1    g081(.A(G92gat), .ZN(new_n283_));
  NOR2_X1   g082(.A1(new_n282_), .A2(new_n283_), .ZN(new_n284_));
  NOR2_X1   g083(.A1(KEYINPUT65), .A2(KEYINPUT9), .ZN(new_n285_));
  AOI22_X1  g084(.A1(new_n275_), .A2(new_n281_), .B1(new_n284_), .B2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT10), .B(G99gat), .ZN(new_n287_));
  OAI221_X1 g086(.A(new_n286_), .B1(G106gat), .B2(new_n287_), .C1(new_n273_), .C2(new_n272_), .ZN(new_n288_));
  AOI21_X1  g087(.A(new_n259_), .B1(new_n280_), .B2(new_n288_), .ZN(new_n289_));
  AND3_X1   g088(.A1(new_n274_), .A2(new_n278_), .A3(new_n275_), .ZN(new_n290_));
  AOI21_X1  g089(.A(new_n278_), .B1(new_n274_), .B2(new_n275_), .ZN(new_n291_));
  OAI211_X1 g090(.A(new_n259_), .B(new_n288_), .C1(new_n290_), .C2(new_n291_), .ZN(new_n292_));
  INV_X1    g091(.A(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n258_), .B1(new_n289_), .B2(new_n293_), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n295_));
  OAI21_X1  g094(.A(new_n288_), .B1(new_n290_), .B2(new_n291_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT68), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n297_), .A2(new_n292_), .A3(new_n257_), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n294_), .A2(new_n295_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G230gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT64), .ZN(new_n301_));
  OAI211_X1 g100(.A(new_n299_), .B(new_n301_), .C1(new_n295_), .C2(new_n294_), .ZN(new_n302_));
  XOR2_X1   g101(.A(G120gat), .B(G148gat), .Z(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(G204gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(KEYINPUT5), .B(G176gat), .ZN(new_n305_));
  XOR2_X1   g104(.A(new_n304_), .B(new_n305_), .Z(new_n306_));
  INV_X1    g105(.A(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n307_), .A2(KEYINPUT71), .ZN(new_n308_));
  INV_X1    g107(.A(new_n301_), .ZN(new_n309_));
  AND2_X1   g108(.A1(new_n298_), .A2(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT12), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n294_), .A2(new_n311_), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n258_), .A2(KEYINPUT12), .A3(new_n296_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n302_), .A2(new_n308_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  AOI21_X1  g115(.A(new_n308_), .B1(new_n302_), .B2(new_n314_), .ZN(new_n317_));
  OAI211_X1 g116(.A(new_n241_), .B(new_n242_), .C1(new_n316_), .C2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n319_), .A2(KEYINPUT72), .A3(KEYINPUT13), .A4(new_n315_), .ZN(new_n320_));
  INV_X1    g119(.A(G211gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G127gat), .B(G155gat), .ZN(new_n322_));
  INV_X1    g121(.A(KEYINPUT16), .ZN(new_n323_));
  OR2_X1    g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n322_), .A2(new_n323_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n326_), .A2(G183gat), .ZN(new_n327_));
  XNOR2_X1  g126(.A(new_n322_), .B(KEYINPUT16), .ZN(new_n328_));
  INV_X1    g127(.A(G183gat), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n328_), .A2(new_n329_), .ZN(new_n330_));
  OAI21_X1  g129(.A(new_n321_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT17), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n326_), .A2(G183gat), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n328_), .A2(new_n329_), .ZN(new_n334_));
  NAND3_X1  g133(.A1(new_n333_), .A2(new_n334_), .A3(G211gat), .ZN(new_n335_));
  AND3_X1   g134(.A1(new_n331_), .A2(new_n332_), .A3(new_n335_), .ZN(new_n336_));
  AOI21_X1  g135(.A(new_n332_), .B1(new_n331_), .B2(new_n335_), .ZN(new_n337_));
  NOR2_X1   g136(.A1(new_n336_), .A2(new_n337_), .ZN(new_n338_));
  INV_X1    g137(.A(new_n211_), .ZN(new_n339_));
  OAI21_X1  g138(.A(new_n339_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n248_), .A2(new_n252_), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n250_), .A2(KEYINPUT11), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n343_), .A2(new_n211_), .A3(new_n254_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(G231gat), .A2(G233gat), .ZN(new_n345_));
  AND3_X1   g144(.A1(new_n340_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n346_));
  AOI21_X1  g145(.A(new_n345_), .B1(new_n340_), .B2(new_n344_), .ZN(new_n347_));
  NOR3_X1   g146(.A1(new_n338_), .A2(new_n346_), .A3(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n340_), .A2(new_n344_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n345_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n349_), .A2(new_n350_), .ZN(new_n351_));
  NAND3_X1  g150(.A1(new_n340_), .A2(new_n344_), .A3(new_n345_), .ZN(new_n352_));
  AOI21_X1  g151(.A(new_n337_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n353_));
  OAI21_X1  g152(.A(KEYINPUT74), .B1(new_n348_), .B2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(new_n337_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n355_), .B1(new_n346_), .B2(new_n347_), .ZN(new_n356_));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n351_), .A2(new_n352_), .ZN(new_n358_));
  OAI211_X1 g157(.A(new_n356_), .B(new_n357_), .C1(new_n358_), .C2(new_n338_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n354_), .A2(new_n359_), .ZN(new_n360_));
  XNOR2_X1  g159(.A(G190gat), .B(G218gat), .ZN(new_n361_));
  XNOR2_X1  g160(.A(G134gat), .B(G162gat), .ZN(new_n362_));
  XNOR2_X1  g161(.A(new_n361_), .B(new_n362_), .ZN(new_n363_));
  XOR2_X1   g162(.A(new_n363_), .B(KEYINPUT36), .Z(new_n364_));
  NAND3_X1  g163(.A1(new_n297_), .A2(new_n216_), .A3(new_n292_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(G232gat), .A2(G233gat), .ZN(new_n366_));
  XNOR2_X1  g165(.A(new_n366_), .B(KEYINPUT73), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT34), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT35), .ZN(new_n369_));
  OR2_X1    g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  AND2_X1   g169(.A1(new_n225_), .A2(new_n226_), .ZN(new_n371_));
  AOI22_X1  g170(.A1(new_n296_), .A2(new_n371_), .B1(new_n369_), .B2(new_n368_), .ZN(new_n372_));
  NAND3_X1  g171(.A1(new_n365_), .A2(new_n370_), .A3(new_n372_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(new_n370_), .B1(new_n365_), .B2(new_n372_), .ZN(new_n375_));
  OAI21_X1  g174(.A(new_n364_), .B1(new_n374_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n375_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n363_), .A2(KEYINPUT36), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n377_), .A2(new_n378_), .A3(new_n373_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n376_), .A2(new_n379_), .A3(KEYINPUT37), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT37), .B1(new_n376_), .B2(new_n379_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND4_X1  g181(.A1(new_n318_), .A2(new_n320_), .A3(new_n360_), .A4(new_n382_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n240_), .B1(new_n383_), .B2(KEYINPUT75), .ZN(new_n384_));
  INV_X1    g183(.A(G176gat), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n385_), .A2(KEYINPUT78), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT78), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n387_), .A2(G176gat), .ZN(new_n388_));
  INV_X1    g187(.A(G169gat), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT22), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT22), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(G169gat), .ZN(new_n392_));
  NAND4_X1  g191(.A1(new_n386_), .A2(new_n388_), .A3(new_n390_), .A4(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G169gat), .A2(G176gat), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n393_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(G190gat), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n329_), .A2(new_n396_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT23), .ZN(new_n398_));
  AOI21_X1  g197(.A(new_n398_), .B1(G183gat), .B2(G190gat), .ZN(new_n399_));
  NAND2_X1  g198(.A1(G183gat), .A2(G190gat), .ZN(new_n400_));
  NOR2_X1   g199(.A1(new_n400_), .A2(KEYINPUT23), .ZN(new_n401_));
  OAI21_X1  g200(.A(new_n397_), .B1(new_n399_), .B2(new_n401_), .ZN(new_n402_));
  NAND2_X1  g201(.A1(new_n402_), .A2(KEYINPUT89), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n400_), .A2(KEYINPUT23), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n398_), .A2(G183gat), .A3(G190gat), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(KEYINPUT89), .ZN(new_n407_));
  NAND3_X1  g206(.A1(new_n406_), .A2(new_n407_), .A3(new_n397_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n395_), .B1(new_n403_), .B2(new_n408_), .ZN(new_n409_));
  XOR2_X1   g208(.A(G211gat), .B(G218gat), .Z(new_n410_));
  INV_X1    g209(.A(KEYINPUT21), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n410_), .A2(new_n411_), .ZN(new_n412_));
  XOR2_X1   g211(.A(G197gat), .B(G204gat), .Z(new_n413_));
  XNOR2_X1  g212(.A(G211gat), .B(G218gat), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n414_), .A2(KEYINPUT21), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n412_), .A2(new_n413_), .A3(new_n415_), .ZN(new_n416_));
  INV_X1    g215(.A(new_n413_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n417_), .A2(KEYINPUT21), .A3(new_n414_), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n416_), .A2(new_n418_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n399_), .A2(KEYINPUT79), .ZN(new_n420_));
  NOR3_X1   g219(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n421_));
  INV_X1    g220(.A(KEYINPUT24), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n422_), .B1(G169gat), .B2(G176gat), .ZN(new_n423_));
  NAND2_X1  g222(.A1(new_n389_), .A2(new_n385_), .ZN(new_n424_));
  AOI21_X1  g223(.A(new_n421_), .B1(new_n423_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(KEYINPUT79), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n404_), .A2(new_n405_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n329_), .A2(KEYINPUT25), .ZN(new_n428_));
  INV_X1    g227(.A(KEYINPUT25), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n429_), .A2(G183gat), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n396_), .A2(KEYINPUT26), .ZN(new_n431_));
  INV_X1    g230(.A(KEYINPUT26), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n432_), .A2(G190gat), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n428_), .A2(new_n430_), .A3(new_n431_), .A4(new_n433_), .ZN(new_n434_));
  AND4_X1   g233(.A1(new_n420_), .A2(new_n425_), .A3(new_n427_), .A4(new_n434_), .ZN(new_n435_));
  OR3_X1    g234(.A1(new_n409_), .A2(new_n419_), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(G226gat), .A2(G233gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT19), .ZN(new_n438_));
  INV_X1    g237(.A(new_n438_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n420_), .A2(new_n427_), .A3(new_n397_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n440_), .A2(new_n394_), .A3(new_n393_), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n434_), .A2(KEYINPUT77), .ZN(new_n442_));
  XNOR2_X1  g241(.A(KEYINPUT25), .B(G183gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(KEYINPUT26), .B(G190gat), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT77), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n443_), .A2(new_n444_), .A3(new_n445_), .ZN(new_n446_));
  NAND4_X1  g245(.A1(new_n442_), .A2(new_n406_), .A3(new_n425_), .A4(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n441_), .A2(new_n447_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n448_), .A2(new_n419_), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n436_), .A2(KEYINPUT20), .A3(new_n439_), .A4(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(G8gat), .B(G36gat), .ZN(new_n451_));
  XNOR2_X1  g250(.A(new_n451_), .B(KEYINPUT18), .ZN(new_n452_));
  XNOR2_X1  g251(.A(new_n452_), .B(G64gat), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n453_), .B(new_n283_), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n419_), .B1(new_n409_), .B2(new_n435_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n441_), .A2(new_n447_), .A3(new_n418_), .A4(new_n416_), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n455_), .A2(KEYINPUT20), .A3(new_n456_), .ZN(new_n457_));
  INV_X1    g256(.A(KEYINPUT90), .ZN(new_n458_));
  AND3_X1   g257(.A1(new_n457_), .A2(new_n458_), .A3(new_n438_), .ZN(new_n459_));
  AOI21_X1  g258(.A(new_n458_), .B1(new_n457_), .B2(new_n438_), .ZN(new_n460_));
  OAI211_X1 g259(.A(new_n450_), .B(new_n454_), .C1(new_n459_), .C2(new_n460_), .ZN(new_n461_));
  XOR2_X1   g260(.A(KEYINPUT94), .B(KEYINPUT20), .Z(new_n462_));
  NAND3_X1  g261(.A1(new_n436_), .A2(new_n449_), .A3(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT95), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n463_), .A2(new_n464_), .A3(new_n438_), .ZN(new_n465_));
  AOI21_X1  g264(.A(new_n464_), .B1(new_n463_), .B2(new_n438_), .ZN(new_n466_));
  NOR2_X1   g265(.A1(new_n457_), .A2(new_n438_), .ZN(new_n467_));
  NOR3_X1   g266(.A1(new_n465_), .A2(new_n466_), .A3(new_n467_), .ZN(new_n468_));
  OAI211_X1 g267(.A(KEYINPUT27), .B(new_n461_), .C1(new_n468_), .C2(new_n454_), .ZN(new_n469_));
  INV_X1    g268(.A(KEYINPUT27), .ZN(new_n470_));
  NAND2_X1  g269(.A1(new_n457_), .A2(new_n438_), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT90), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n457_), .A2(new_n458_), .A3(new_n438_), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n472_), .A2(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n454_), .B1(new_n474_), .B2(new_n450_), .ZN(new_n475_));
  INV_X1    g274(.A(new_n461_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n470_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  AND2_X1   g276(.A1(new_n469_), .A2(new_n477_), .ZN(new_n478_));
  OAI21_X1  g277(.A(KEYINPUT81), .B1(G155gat), .B2(G162gat), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  NOR3_X1   g279(.A1(KEYINPUT81), .A2(G155gat), .A3(G162gat), .ZN(new_n481_));
  OR2_X1    g280(.A1(new_n480_), .A2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G155gat), .A2(G162gat), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n484_));
  INV_X1    g283(.A(KEYINPUT82), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n484_), .B(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT3), .ZN(new_n487_));
  INV_X1    g286(.A(G141gat), .ZN(new_n488_));
  INV_X1    g287(.A(G148gat), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n487_), .A2(new_n488_), .A3(new_n489_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n491_));
  OAI21_X1  g290(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n492_));
  NAND3_X1  g291(.A1(new_n490_), .A2(new_n491_), .A3(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n482_), .B(new_n483_), .C1(new_n486_), .C2(new_n493_), .ZN(new_n494_));
  NAND2_X1  g293(.A1(G141gat), .A2(G148gat), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n488_), .A2(new_n489_), .ZN(new_n496_));
  NOR2_X1   g295(.A1(new_n480_), .A2(new_n481_), .ZN(new_n497_));
  XNOR2_X1  g296(.A(new_n483_), .B(KEYINPUT1), .ZN(new_n498_));
  OAI211_X1 g297(.A(new_n495_), .B(new_n496_), .C1(new_n497_), .C2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n494_), .A2(new_n499_), .ZN(new_n500_));
  INV_X1    g299(.A(G120gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n501_), .A2(G113gat), .ZN(new_n502_));
  INV_X1    g301(.A(G113gat), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n503_), .A2(G120gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT80), .ZN(new_n505_));
  AND3_X1   g304(.A1(new_n502_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n505_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n507_));
  OAI21_X1  g306(.A(G127gat), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n503_), .A2(G120gat), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n501_), .A2(G113gat), .ZN(new_n510_));
  OAI21_X1  g309(.A(KEYINPUT80), .B1(new_n509_), .B2(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(G127gat), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n502_), .A2(new_n504_), .A3(new_n505_), .ZN(new_n513_));
  NAND3_X1  g312(.A1(new_n511_), .A2(new_n512_), .A3(new_n513_), .ZN(new_n514_));
  AND3_X1   g313(.A1(new_n508_), .A2(new_n514_), .A3(G134gat), .ZN(new_n515_));
  AOI21_X1  g314(.A(G134gat), .B1(new_n508_), .B2(new_n514_), .ZN(new_n516_));
  OAI21_X1  g315(.A(new_n500_), .B1(new_n515_), .B2(new_n516_), .ZN(new_n517_));
  OAI21_X1  g316(.A(new_n483_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n484_), .B(KEYINPUT82), .ZN(new_n519_));
  INV_X1    g318(.A(new_n493_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n518_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n496_), .A2(new_n495_), .ZN(new_n522_));
  INV_X1    g321(.A(KEYINPUT1), .ZN(new_n523_));
  XNOR2_X1  g322(.A(new_n483_), .B(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n522_), .B1(new_n482_), .B2(new_n524_), .ZN(new_n525_));
  NOR2_X1   g324(.A1(new_n521_), .A2(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(G134gat), .ZN(new_n527_));
  NOR3_X1   g326(.A1(new_n506_), .A2(new_n507_), .A3(G127gat), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n512_), .B1(new_n511_), .B2(new_n513_), .ZN(new_n529_));
  OAI21_X1  g328(.A(new_n527_), .B1(new_n528_), .B2(new_n529_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n508_), .A2(new_n514_), .A3(G134gat), .ZN(new_n531_));
  NAND3_X1  g330(.A1(new_n526_), .A2(new_n530_), .A3(new_n531_), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n517_), .A2(new_n532_), .A3(KEYINPUT4), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G225gat), .A2(G233gat), .ZN(new_n534_));
  INV_X1    g333(.A(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(KEYINPUT4), .ZN(new_n536_));
  OAI211_X1 g335(.A(new_n500_), .B(new_n536_), .C1(new_n515_), .C2(new_n516_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n533_), .A2(new_n535_), .A3(new_n537_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n517_), .A2(new_n532_), .A3(new_n534_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n538_), .A2(new_n539_), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G1gat), .B(G29gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(new_n541_), .B(KEYINPUT0), .ZN(new_n542_));
  INV_X1    g341(.A(G57gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(new_n542_), .B(new_n543_), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n544_), .B(new_n282_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n540_), .A2(new_n545_), .ZN(new_n546_));
  XNOR2_X1  g345(.A(new_n544_), .B(G85gat), .ZN(new_n547_));
  NAND3_X1  g346(.A1(new_n538_), .A2(new_n539_), .A3(new_n547_), .ZN(new_n548_));
  NAND2_X1  g347(.A1(new_n546_), .A2(new_n548_), .ZN(new_n549_));
  XNOR2_X1  g348(.A(G71gat), .B(G99gat), .ZN(new_n550_));
  INV_X1    g349(.A(new_n550_), .ZN(new_n551_));
  XNOR2_X1  g350(.A(new_n448_), .B(KEYINPUT30), .ZN(new_n552_));
  XNOR2_X1  g351(.A(G15gat), .B(G43gat), .ZN(new_n553_));
  NOR2_X1   g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n554_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n552_), .A2(new_n553_), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n551_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NOR2_X1   g357(.A1(new_n515_), .A2(new_n516_), .ZN(new_n559_));
  AND2_X1   g358(.A1(new_n559_), .A2(KEYINPUT31), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n559_), .A2(KEYINPUT31), .ZN(new_n561_));
  AND2_X1   g360(.A1(G227gat), .A2(G233gat), .ZN(new_n562_));
  OR3_X1    g361(.A1(new_n560_), .A2(new_n561_), .A3(new_n562_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n562_), .B1(new_n560_), .B2(new_n561_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n555_), .A2(new_n551_), .A3(new_n556_), .ZN(new_n565_));
  NAND4_X1  g364(.A1(new_n558_), .A2(new_n563_), .A3(new_n564_), .A4(new_n565_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n564_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n565_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n567_), .B1(new_n568_), .B2(new_n557_), .ZN(new_n569_));
  AOI21_X1  g368(.A(new_n549_), .B1(new_n566_), .B2(new_n569_), .ZN(new_n570_));
  XNOR2_X1  g369(.A(G22gat), .B(G50gat), .ZN(new_n571_));
  XNOR2_X1  g370(.A(new_n571_), .B(KEYINPUT28), .ZN(new_n572_));
  OAI21_X1  g371(.A(new_n572_), .B1(new_n500_), .B2(KEYINPUT29), .ZN(new_n573_));
  INV_X1    g372(.A(KEYINPUT29), .ZN(new_n574_));
  INV_X1    g373(.A(new_n572_), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n526_), .A2(new_n574_), .A3(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n577_), .B(KEYINPUT83), .ZN(new_n578_));
  NAND2_X1  g377(.A1(G228gat), .A2(G233gat), .ZN(new_n579_));
  INV_X1    g378(.A(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT86), .ZN(new_n581_));
  XNOR2_X1  g380(.A(KEYINPUT85), .B(KEYINPUT29), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  OAI211_X1 g382(.A(new_n581_), .B(new_n583_), .C1(new_n521_), .C2(new_n525_), .ZN(new_n584_));
  NAND2_X1  g383(.A1(new_n584_), .A2(new_n419_), .ZN(new_n585_));
  AOI21_X1  g384(.A(new_n581_), .B1(new_n500_), .B2(new_n583_), .ZN(new_n586_));
  OAI21_X1  g385(.A(new_n580_), .B1(new_n585_), .B2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT84), .ZN(new_n588_));
  AOI21_X1  g387(.A(new_n574_), .B1(new_n494_), .B2(new_n499_), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n419_), .A2(new_n579_), .ZN(new_n590_));
  OAI21_X1  g389(.A(new_n588_), .B1(new_n589_), .B2(new_n590_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n580_), .B1(new_n416_), .B2(new_n418_), .ZN(new_n592_));
  OAI211_X1 g391(.A(new_n592_), .B(KEYINPUT84), .C1(new_n526_), .C2(new_n574_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n591_), .A2(new_n593_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G78gat), .B(G106gat), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  AND3_X1   g395(.A1(new_n587_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n597_));
  AOI21_X1  g396(.A(new_n596_), .B1(new_n587_), .B2(new_n594_), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n578_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  NAND2_X1  g398(.A1(new_n599_), .A2(KEYINPUT87), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT87), .ZN(new_n601_));
  OAI211_X1 g400(.A(new_n578_), .B(new_n601_), .C1(new_n597_), .C2(new_n598_), .ZN(new_n602_));
  INV_X1    g401(.A(KEYINPUT88), .ZN(new_n603_));
  AND2_X1   g402(.A1(new_n587_), .A2(new_n594_), .ZN(new_n604_));
  OAI21_X1  g403(.A(new_n603_), .B1(new_n604_), .B2(new_n596_), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n598_), .A2(KEYINPUT88), .ZN(new_n606_));
  NAND2_X1  g405(.A1(new_n605_), .A2(new_n606_), .ZN(new_n607_));
  NAND3_X1  g406(.A1(new_n587_), .A2(new_n594_), .A3(new_n596_), .ZN(new_n608_));
  AND2_X1   g407(.A1(new_n608_), .A2(new_n577_), .ZN(new_n609_));
  AOI22_X1  g408(.A1(new_n600_), .A2(new_n602_), .B1(new_n607_), .B2(new_n609_), .ZN(new_n610_));
  NAND3_X1  g409(.A1(new_n478_), .A2(new_n570_), .A3(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n612_));
  XNOR2_X1  g411(.A(new_n611_), .B(new_n612_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n469_), .A2(new_n477_), .ZN(new_n614_));
  NOR3_X1   g413(.A1(new_n614_), .A2(new_n610_), .A3(new_n549_), .ZN(new_n615_));
  INV_X1    g414(.A(KEYINPUT91), .ZN(new_n616_));
  OAI21_X1  g415(.A(new_n616_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n617_));
  OAI21_X1  g416(.A(new_n450_), .B1(new_n459_), .B2(new_n460_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n454_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n618_), .A2(new_n619_), .ZN(new_n620_));
  NAND3_X1  g419(.A1(new_n620_), .A2(KEYINPUT91), .A3(new_n461_), .ZN(new_n621_));
  AND2_X1   g420(.A1(KEYINPUT92), .A2(KEYINPUT33), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n548_), .B(new_n622_), .ZN(new_n623_));
  NOR2_X1   g422(.A1(KEYINPUT92), .A2(KEYINPUT33), .ZN(new_n624_));
  AND2_X1   g423(.A1(new_n537_), .A2(new_n534_), .ZN(new_n625_));
  AND2_X1   g424(.A1(new_n625_), .A2(new_n533_), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n517_), .A2(new_n532_), .A3(new_n535_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n545_), .A2(new_n627_), .ZN(new_n628_));
  OAI21_X1  g427(.A(KEYINPUT93), .B1(new_n626_), .B2(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n625_), .A2(new_n533_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT93), .ZN(new_n631_));
  NAND4_X1  g430(.A1(new_n630_), .A2(new_n631_), .A3(new_n545_), .A4(new_n627_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n624_), .B1(new_n629_), .B2(new_n632_), .ZN(new_n633_));
  NAND4_X1  g432(.A1(new_n617_), .A2(new_n621_), .A3(new_n623_), .A4(new_n633_), .ZN(new_n634_));
  NAND2_X1  g433(.A1(new_n454_), .A2(KEYINPUT32), .ZN(new_n635_));
  NAND3_X1  g434(.A1(new_n474_), .A2(new_n450_), .A3(new_n635_), .ZN(new_n636_));
  OAI211_X1 g435(.A(new_n549_), .B(new_n636_), .C1(new_n468_), .C2(new_n635_), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n634_), .A2(new_n637_), .ZN(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(new_n610_), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n615_), .B1(new_n639_), .B2(KEYINPUT96), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n600_), .A2(new_n602_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n607_), .A2(new_n609_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n643_), .B1(new_n634_), .B2(new_n637_), .ZN(new_n644_));
  INV_X1    g443(.A(KEYINPUT96), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n640_), .A2(new_n646_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n566_), .A2(new_n569_), .ZN(new_n648_));
  INV_X1    g447(.A(new_n648_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n613_), .B1(new_n647_), .B2(new_n649_), .ZN(new_n650_));
  AOI211_X1 g449(.A(new_n384_), .B(new_n650_), .C1(KEYINPUT75), .C2(new_n383_), .ZN(new_n651_));
  NAND3_X1  g450(.A1(new_n651_), .A2(new_n204_), .A3(new_n549_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT38), .ZN(new_n653_));
  INV_X1    g452(.A(new_n376_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n379_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n650_), .A2(new_n656_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n318_), .A2(new_n320_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n360_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n240_), .ZN(new_n660_));
  NOR3_X1   g459(.A1(new_n658_), .A2(new_n659_), .A3(new_n660_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n657_), .A2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(new_n549_), .ZN(new_n663_));
  OAI21_X1  g462(.A(G1gat), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n653_), .A2(new_n664_), .ZN(G1324gat));
  NAND3_X1  g464(.A1(new_n651_), .A2(new_n205_), .A3(new_n614_), .ZN(new_n666_));
  NAND3_X1  g465(.A1(new_n657_), .A2(new_n614_), .A3(new_n661_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT39), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G8gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G8gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n671_), .A2(KEYINPUT98), .ZN(new_n672_));
  INV_X1    g471(.A(KEYINPUT98), .ZN(new_n673_));
  OAI211_X1 g472(.A(new_n666_), .B(new_n673_), .C1(new_n669_), .C2(new_n670_), .ZN(new_n674_));
  AND3_X1   g473(.A1(new_n672_), .A2(KEYINPUT40), .A3(new_n674_), .ZN(new_n675_));
  AOI21_X1  g474(.A(KEYINPUT40), .B1(new_n672_), .B2(new_n674_), .ZN(new_n676_));
  NOR2_X1   g475(.A1(new_n675_), .A2(new_n676_), .ZN(G1325gat));
  INV_X1    g476(.A(G15gat), .ZN(new_n678_));
  NAND3_X1  g477(.A1(new_n651_), .A2(new_n678_), .A3(new_n648_), .ZN(new_n679_));
  NAND3_X1  g478(.A1(new_n657_), .A2(new_n648_), .A3(new_n661_), .ZN(new_n680_));
  AND3_X1   g479(.A1(new_n680_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n681_));
  AOI21_X1  g480(.A(KEYINPUT41), .B1(new_n680_), .B2(G15gat), .ZN(new_n682_));
  OAI21_X1  g481(.A(new_n679_), .B1(new_n681_), .B2(new_n682_), .ZN(new_n683_));
  XOR2_X1   g482(.A(new_n683_), .B(KEYINPUT99), .Z(G1326gat));
  XNOR2_X1  g483(.A(new_n610_), .B(KEYINPUT100), .ZN(new_n685_));
  OAI21_X1  g484(.A(G22gat), .B1(new_n662_), .B2(new_n685_), .ZN(new_n686_));
  XNOR2_X1  g485(.A(KEYINPUT101), .B(KEYINPUT42), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(new_n688_));
  INV_X1    g487(.A(G22gat), .ZN(new_n689_));
  INV_X1    g488(.A(new_n685_), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n651_), .A2(new_n689_), .A3(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n688_), .A2(new_n691_), .ZN(G1327gat));
  INV_X1    g491(.A(new_n646_), .ZN(new_n693_));
  NOR2_X1   g492(.A1(new_n610_), .A2(new_n549_), .ZN(new_n694_));
  NAND2_X1  g493(.A1(new_n694_), .A2(new_n478_), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n695_), .B1(new_n644_), .B2(new_n645_), .ZN(new_n696_));
  OAI21_X1  g495(.A(new_n649_), .B1(new_n693_), .B2(new_n696_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n611_), .B(KEYINPUT97), .ZN(new_n698_));
  AOI21_X1  g497(.A(new_n382_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  OAI21_X1  g498(.A(KEYINPUT43), .B1(new_n699_), .B2(KEYINPUT103), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT43), .ZN(new_n702_));
  OAI211_X1 g501(.A(new_n701_), .B(new_n702_), .C1(new_n650_), .C2(new_n382_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n658_), .A2(new_n360_), .A3(new_n660_), .ZN(new_n704_));
  XNOR2_X1  g503(.A(new_n704_), .B(KEYINPUT102), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n700_), .A2(new_n703_), .A3(KEYINPUT44), .A4(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n706_), .A2(G29gat), .A3(new_n549_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n700_), .A2(new_n703_), .A3(new_n705_), .ZN(new_n708_));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n710_), .A2(KEYINPUT104), .ZN(new_n711_));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n708_), .A2(new_n712_), .A3(new_n709_), .ZN(new_n713_));
  AOI21_X1  g512(.A(new_n707_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n714_));
  INV_X1    g513(.A(KEYINPUT105), .ZN(new_n715_));
  INV_X1    g514(.A(new_n656_), .ZN(new_n716_));
  NOR2_X1   g515(.A1(new_n650_), .A2(new_n716_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n717_), .A2(new_n704_), .ZN(new_n718_));
  AOI21_X1  g517(.A(G29gat), .B1(new_n718_), .B2(new_n549_), .ZN(new_n719_));
  OR3_X1    g518(.A1(new_n714_), .A2(new_n715_), .A3(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n715_), .B1(new_n714_), .B2(new_n719_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n720_), .A2(new_n721_), .ZN(G1328gat));
  OR2_X1    g521(.A1(new_n614_), .A2(KEYINPUT106), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n614_), .A2(KEYINPUT106), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(new_n725_), .ZN(new_n726_));
  NOR2_X1   g525(.A1(new_n726_), .A2(G36gat), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n717_), .A2(new_n704_), .A3(new_n727_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n728_), .A2(KEYINPUT107), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n730_));
  NAND4_X1  g529(.A1(new_n717_), .A2(new_n730_), .A3(new_n704_), .A4(new_n727_), .ZN(new_n731_));
  AND3_X1   g530(.A1(new_n729_), .A2(KEYINPUT45), .A3(new_n731_), .ZN(new_n732_));
  AOI21_X1  g531(.A(KEYINPUT45), .B1(new_n729_), .B2(new_n731_), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n706_), .A2(new_n614_), .ZN(new_n735_));
  AOI21_X1  g534(.A(new_n735_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n736_));
  INV_X1    g535(.A(G36gat), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n734_), .B1(new_n736_), .B2(new_n737_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n738_), .A2(new_n739_), .ZN(new_n740_));
  OAI211_X1 g539(.A(new_n734_), .B(KEYINPUT46), .C1(new_n736_), .C2(new_n737_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1329gat));
  NAND3_X1  g541(.A1(new_n706_), .A2(G43gat), .A3(new_n648_), .ZN(new_n743_));
  AOI21_X1  g542(.A(new_n743_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n744_));
  AOI21_X1  g543(.A(G43gat), .B1(new_n718_), .B2(new_n648_), .ZN(new_n745_));
  OR3_X1    g544(.A1(new_n744_), .A2(KEYINPUT47), .A3(new_n745_), .ZN(new_n746_));
  OAI21_X1  g545(.A(KEYINPUT47), .B1(new_n744_), .B2(new_n745_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n746_), .A2(new_n747_), .ZN(G1330gat));
  NOR2_X1   g547(.A1(new_n685_), .A2(G50gat), .ZN(new_n749_));
  XNOR2_X1  g548(.A(new_n749_), .B(KEYINPUT108), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n718_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n706_), .A2(new_n643_), .ZN(new_n752_));
  AOI21_X1  g551(.A(new_n752_), .B1(new_n711_), .B2(new_n713_), .ZN(new_n753_));
  INV_X1    g552(.A(G50gat), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n751_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND2_X1  g554(.A1(new_n755_), .A2(KEYINPUT109), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n757_));
  OAI211_X1 g556(.A(new_n757_), .B(new_n751_), .C1(new_n753_), .C2(new_n754_), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n756_), .A2(new_n758_), .ZN(G1331gat));
  NAND2_X1  g558(.A1(new_n697_), .A2(new_n698_), .ZN(new_n760_));
  NAND2_X1  g559(.A1(new_n658_), .A2(new_n660_), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n761_), .A2(new_n659_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n760_), .A2(new_n382_), .A3(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n543_), .B1(new_n763_), .B2(new_n663_), .ZN(new_n764_));
  XOR2_X1   g563(.A(new_n764_), .B(KEYINPUT110), .Z(new_n765_));
  AOI21_X1  g564(.A(new_n648_), .B1(new_n640_), .B2(new_n646_), .ZN(new_n766_));
  OAI211_X1 g565(.A(new_n716_), .B(new_n762_), .C1(new_n766_), .C2(new_n613_), .ZN(new_n767_));
  NAND2_X1  g566(.A1(new_n767_), .A2(KEYINPUT111), .ZN(new_n768_));
  INV_X1    g567(.A(KEYINPUT111), .ZN(new_n769_));
  NAND4_X1  g568(.A1(new_n760_), .A2(new_n769_), .A3(new_n716_), .A4(new_n762_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n768_), .A2(new_n770_), .ZN(new_n771_));
  NOR3_X1   g570(.A1(new_n771_), .A2(new_n543_), .A3(new_n663_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n765_), .A2(new_n772_), .ZN(G1332gat));
  OR3_X1    g572(.A1(new_n763_), .A2(G64gat), .A3(new_n726_), .ZN(new_n774_));
  NAND3_X1  g573(.A1(new_n768_), .A2(new_n725_), .A3(new_n770_), .ZN(new_n775_));
  INV_X1    g574(.A(KEYINPUT112), .ZN(new_n776_));
  NAND3_X1  g575(.A1(new_n775_), .A2(new_n776_), .A3(G64gat), .ZN(new_n777_));
  INV_X1    g576(.A(new_n777_), .ZN(new_n778_));
  AOI21_X1  g577(.A(new_n776_), .B1(new_n775_), .B2(G64gat), .ZN(new_n779_));
  INV_X1    g578(.A(KEYINPUT48), .ZN(new_n780_));
  NOR3_X1   g579(.A1(new_n778_), .A2(new_n779_), .A3(new_n780_), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n775_), .A2(G64gat), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(KEYINPUT112), .ZN(new_n783_));
  AOI21_X1  g582(.A(KEYINPUT48), .B1(new_n783_), .B2(new_n777_), .ZN(new_n784_));
  OAI21_X1  g583(.A(new_n774_), .B1(new_n781_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(new_n787_));
  OAI211_X1 g586(.A(KEYINPUT113), .B(new_n774_), .C1(new_n781_), .C2(new_n784_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(G1333gat));
  OR3_X1    g588(.A1(new_n763_), .A2(G71gat), .A3(new_n649_), .ZN(new_n790_));
  OAI21_X1  g589(.A(G71gat), .B1(new_n771_), .B2(new_n649_), .ZN(new_n791_));
  AND2_X1   g590(.A1(new_n791_), .A2(KEYINPUT49), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n791_), .A2(KEYINPUT49), .ZN(new_n793_));
  OAI21_X1  g592(.A(new_n790_), .B1(new_n792_), .B2(new_n793_), .ZN(G1334gat));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n795_));
  INV_X1    g594(.A(new_n771_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n690_), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n795_), .B1(new_n797_), .B2(G78gat), .ZN(new_n798_));
  INV_X1    g597(.A(G78gat), .ZN(new_n799_));
  AOI211_X1 g598(.A(KEYINPUT50), .B(new_n799_), .C1(new_n796_), .C2(new_n690_), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n690_), .A2(new_n799_), .ZN(new_n801_));
  OAI22_X1  g600(.A1(new_n798_), .A2(new_n800_), .B1(new_n763_), .B2(new_n801_), .ZN(G1335gat));
  NOR2_X1   g601(.A1(new_n761_), .A2(new_n360_), .ZN(new_n803_));
  NAND2_X1  g602(.A1(new_n717_), .A2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(new_n804_), .ZN(new_n805_));
  NAND3_X1  g604(.A1(new_n805_), .A2(new_n282_), .A3(new_n549_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n700_), .A2(new_n703_), .A3(new_n803_), .ZN(new_n807_));
  OR2_X1    g606(.A1(new_n807_), .A2(KEYINPUT114), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n807_), .A2(KEYINPUT114), .ZN(new_n809_));
  AOI21_X1  g608(.A(new_n663_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n810_));
  OAI21_X1  g609(.A(new_n806_), .B1(new_n810_), .B2(new_n282_), .ZN(G1336gat));
  NAND3_X1  g610(.A1(new_n805_), .A2(new_n283_), .A3(new_n614_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n726_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n812_), .B1(new_n813_), .B2(new_n283_), .ZN(G1337gat));
  NOR3_X1   g613(.A1(new_n804_), .A2(new_n287_), .A3(new_n649_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n649_), .B1(new_n808_), .B2(new_n809_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n816_), .B1(new_n817_), .B2(new_n261_), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n818_), .A2(KEYINPUT51), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT51), .ZN(new_n820_));
  OAI211_X1 g619(.A(new_n820_), .B(new_n816_), .C1(new_n817_), .C2(new_n261_), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n819_), .A2(new_n821_), .ZN(G1338gat));
  NAND3_X1  g621(.A1(new_n805_), .A2(new_n262_), .A3(new_n643_), .ZN(new_n823_));
  NAND4_X1  g622(.A1(new_n700_), .A2(new_n703_), .A3(new_n643_), .A4(new_n803_), .ZN(new_n824_));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n824_), .A2(new_n825_), .A3(G106gat), .ZN(new_n826_));
  AOI21_X1  g625(.A(new_n825_), .B1(new_n824_), .B2(G106gat), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n823_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  XNOR2_X1  g627(.A(new_n828_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g628(.A(KEYINPUT118), .ZN(new_n830_));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n220_), .A2(new_n221_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n227_), .A2(new_n219_), .A3(new_n222_), .ZN(new_n833_));
  NAND3_X1  g632(.A1(new_n832_), .A2(new_n236_), .A3(new_n833_), .ZN(new_n834_));
  AND2_X1   g633(.A1(new_n834_), .A2(new_n238_), .ZN(new_n835_));
  INV_X1    g634(.A(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n319_), .B2(new_n315_), .ZN(new_n837_));
  INV_X1    g636(.A(KEYINPUT55), .ZN(new_n838_));
  AOI21_X1  g637(.A(new_n257_), .B1(new_n297_), .B2(new_n292_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n313_), .B1(new_n839_), .B2(KEYINPUT12), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n298_), .A2(new_n309_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n838_), .B1(new_n840_), .B2(new_n841_), .ZN(new_n842_));
  NAND4_X1  g641(.A1(new_n310_), .A2(new_n312_), .A3(KEYINPUT55), .A4(new_n313_), .ZN(new_n843_));
  OAI211_X1 g642(.A(new_n313_), .B(new_n298_), .C1(new_n839_), .C2(KEYINPUT12), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n301_), .ZN(new_n845_));
  NAND3_X1  g644(.A1(new_n842_), .A2(new_n843_), .A3(new_n845_), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n846_), .A2(new_n307_), .ZN(new_n847_));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n848_));
  NAND2_X1  g647(.A1(new_n847_), .A2(new_n848_), .ZN(new_n849_));
  NOR2_X1   g648(.A1(new_n306_), .A2(new_n848_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n846_), .A2(new_n850_), .ZN(new_n851_));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n851_), .A2(new_n852_), .ZN(new_n853_));
  NAND3_X1  g652(.A1(new_n846_), .A2(KEYINPUT116), .A3(new_n850_), .ZN(new_n854_));
  NAND3_X1  g653(.A1(new_n849_), .A2(new_n853_), .A3(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n302_), .A2(new_n306_), .A3(new_n314_), .ZN(new_n856_));
  NAND2_X1  g655(.A1(new_n856_), .A2(new_n240_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  AOI21_X1  g657(.A(new_n837_), .B1(new_n855_), .B2(new_n858_), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n831_), .B1(new_n859_), .B2(new_n656_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT58), .ZN(new_n861_));
  AOI21_X1  g660(.A(KEYINPUT56), .B1(new_n846_), .B2(new_n307_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n862_), .B1(new_n846_), .B2(new_n850_), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n856_), .A2(new_n835_), .ZN(new_n864_));
  INV_X1    g663(.A(KEYINPUT117), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n864_), .A2(new_n865_), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n856_), .A2(KEYINPUT117), .A3(new_n835_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n861_), .B1(new_n863_), .B2(new_n868_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n849_), .A2(new_n851_), .ZN(new_n870_));
  NAND4_X1  g669(.A1(new_n870_), .A2(KEYINPUT58), .A3(new_n867_), .A4(new_n866_), .ZN(new_n871_));
  INV_X1    g670(.A(new_n382_), .ZN(new_n872_));
  NAND3_X1  g671(.A1(new_n869_), .A2(new_n871_), .A3(new_n872_), .ZN(new_n873_));
  AOI21_X1  g672(.A(KEYINPUT116), .B1(new_n846_), .B2(new_n850_), .ZN(new_n874_));
  NOR2_X1   g673(.A1(new_n862_), .A2(new_n874_), .ZN(new_n875_));
  AOI21_X1  g674(.A(new_n857_), .B1(new_n875_), .B2(new_n854_), .ZN(new_n876_));
  OAI211_X1 g675(.A(KEYINPUT57), .B(new_n716_), .C1(new_n876_), .C2(new_n837_), .ZN(new_n877_));
  NAND3_X1  g676(.A1(new_n860_), .A2(new_n873_), .A3(new_n877_), .ZN(new_n878_));
  NAND2_X1  g677(.A1(new_n878_), .A2(new_n659_), .ZN(new_n879_));
  AOI21_X1  g678(.A(KEYINPUT115), .B1(new_n360_), .B2(new_n660_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT115), .ZN(new_n881_));
  AOI211_X1 g680(.A(new_n881_), .B(new_n240_), .C1(new_n354_), .C2(new_n359_), .ZN(new_n882_));
  NOR2_X1   g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  NAND4_X1  g682(.A1(new_n883_), .A2(new_n318_), .A3(new_n320_), .A4(new_n382_), .ZN(new_n884_));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n885_));
  XNOR2_X1  g684(.A(new_n884_), .B(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  AOI21_X1  g686(.A(new_n830_), .B1(new_n879_), .B2(new_n887_), .ZN(new_n888_));
  AOI211_X1 g687(.A(KEYINPUT118), .B(new_n886_), .C1(new_n878_), .C2(new_n659_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n649_), .A2(new_n663_), .ZN(new_n890_));
  NOR2_X1   g689(.A1(new_n643_), .A2(new_n614_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NOR3_X1   g691(.A1(new_n888_), .A2(new_n889_), .A3(new_n892_), .ZN(new_n893_));
  AOI21_X1  g692(.A(G113gat), .B1(new_n893_), .B2(new_n240_), .ZN(new_n894_));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n895_));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n888_), .A2(new_n889_), .ZN(new_n897_));
  INV_X1    g696(.A(new_n892_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n896_), .B1(new_n897_), .B2(new_n898_), .ZN(new_n899_));
  NAND3_X1  g698(.A1(new_n860_), .A2(KEYINPUT119), .A3(new_n873_), .ZN(new_n900_));
  NAND2_X1  g699(.A1(new_n900_), .A2(new_n877_), .ZN(new_n901_));
  AOI21_X1  g700(.A(KEYINPUT119), .B1(new_n860_), .B2(new_n873_), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n659_), .B1(new_n901_), .B2(new_n902_), .ZN(new_n903_));
  AOI211_X1 g702(.A(KEYINPUT59), .B(new_n892_), .C1(new_n903_), .C2(new_n887_), .ZN(new_n904_));
  OAI21_X1  g703(.A(new_n895_), .B1(new_n899_), .B2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n887_), .ZN(new_n906_));
  NAND3_X1  g705(.A1(new_n906_), .A2(new_n896_), .A3(new_n898_), .ZN(new_n907_));
  OAI211_X1 g706(.A(new_n907_), .B(KEYINPUT120), .C1(new_n896_), .C2(new_n893_), .ZN(new_n908_));
  NAND2_X1  g707(.A1(new_n905_), .A2(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n240_), .A2(G113gat), .ZN(new_n910_));
  XNOR2_X1  g709(.A(new_n910_), .B(KEYINPUT121), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n894_), .B1(new_n909_), .B2(new_n911_), .ZN(G1340gat));
  OAI211_X1 g711(.A(new_n907_), .B(new_n658_), .C1(new_n896_), .C2(new_n893_), .ZN(new_n913_));
  INV_X1    g712(.A(new_n913_), .ZN(new_n914_));
  XNOR2_X1  g713(.A(KEYINPUT122), .B(G120gat), .ZN(new_n915_));
  INV_X1    g714(.A(new_n893_), .ZN(new_n916_));
  INV_X1    g715(.A(new_n658_), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n915_), .B1(new_n917_), .B2(KEYINPUT60), .ZN(new_n918_));
  OAI21_X1  g717(.A(new_n918_), .B1(KEYINPUT60), .B2(new_n915_), .ZN(new_n919_));
  OAI22_X1  g718(.A1(new_n914_), .A2(new_n915_), .B1(new_n916_), .B2(new_n919_), .ZN(G1341gat));
  NAND3_X1  g719(.A1(new_n897_), .A2(new_n360_), .A3(new_n898_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n921_), .A2(new_n512_), .ZN(new_n922_));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n923_));
  NAND2_X1  g722(.A1(new_n922_), .A2(new_n923_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n921_), .A2(KEYINPUT123), .A3(new_n512_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n924_), .A2(new_n925_), .ZN(new_n926_));
  NOR2_X1   g725(.A1(new_n659_), .A2(new_n512_), .ZN(new_n927_));
  AOI21_X1  g726(.A(new_n926_), .B1(new_n909_), .B2(new_n927_), .ZN(G1342gat));
  NAND3_X1  g727(.A1(new_n893_), .A2(new_n527_), .A3(new_n656_), .ZN(new_n929_));
  AOI21_X1  g728(.A(new_n382_), .B1(new_n905_), .B2(new_n908_), .ZN(new_n930_));
  OAI21_X1  g729(.A(new_n929_), .B1(new_n930_), .B2(new_n527_), .ZN(G1343gat));
  INV_X1    g730(.A(new_n897_), .ZN(new_n932_));
  NAND3_X1  g731(.A1(new_n649_), .A2(new_n549_), .A3(new_n643_), .ZN(new_n933_));
  NOR3_X1   g732(.A1(new_n932_), .A2(new_n725_), .A3(new_n933_), .ZN(new_n934_));
  NAND2_X1  g733(.A1(new_n934_), .A2(new_n240_), .ZN(new_n935_));
  XNOR2_X1  g734(.A(new_n935_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g735(.A1(new_n934_), .A2(new_n658_), .ZN(new_n937_));
  XNOR2_X1  g736(.A(new_n937_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g737(.A1(new_n934_), .A2(new_n360_), .ZN(new_n939_));
  XNOR2_X1  g738(.A(KEYINPUT61), .B(G155gat), .ZN(new_n940_));
  XNOR2_X1  g739(.A(new_n940_), .B(KEYINPUT124), .ZN(new_n941_));
  XNOR2_X1  g740(.A(new_n939_), .B(new_n941_), .ZN(G1346gat));
  INV_X1    g741(.A(G162gat), .ZN(new_n943_));
  NAND3_X1  g742(.A1(new_n934_), .A2(new_n943_), .A3(new_n656_), .ZN(new_n944_));
  AND2_X1   g743(.A1(new_n934_), .A2(new_n872_), .ZN(new_n945_));
  OAI21_X1  g744(.A(new_n944_), .B1(new_n945_), .B2(new_n943_), .ZN(G1347gat));
  AND2_X1   g745(.A1(new_n725_), .A2(new_n570_), .ZN(new_n947_));
  NAND2_X1  g746(.A1(new_n947_), .A2(new_n685_), .ZN(new_n948_));
  AOI21_X1  g747(.A(new_n948_), .B1(new_n903_), .B2(new_n887_), .ZN(new_n949_));
  AOI21_X1  g748(.A(new_n389_), .B1(new_n949_), .B2(new_n240_), .ZN(new_n950_));
  OR2_X1    g749(.A1(new_n950_), .A2(KEYINPUT62), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n950_), .A2(KEYINPUT62), .ZN(new_n952_));
  NAND4_X1  g751(.A1(new_n949_), .A2(new_n390_), .A3(new_n392_), .A4(new_n240_), .ZN(new_n953_));
  NAND4_X1  g752(.A1(new_n951_), .A2(KEYINPUT125), .A3(new_n952_), .A4(new_n953_), .ZN(new_n954_));
  INV_X1    g753(.A(KEYINPUT125), .ZN(new_n955_));
  OAI21_X1  g754(.A(new_n953_), .B1(new_n950_), .B2(KEYINPUT62), .ZN(new_n956_));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n957_));
  AOI211_X1 g756(.A(new_n957_), .B(new_n389_), .C1(new_n949_), .C2(new_n240_), .ZN(new_n958_));
  OAI21_X1  g757(.A(new_n955_), .B1(new_n956_), .B2(new_n958_), .ZN(new_n959_));
  NAND2_X1  g758(.A1(new_n954_), .A2(new_n959_), .ZN(G1348gat));
  NOR2_X1   g759(.A1(new_n932_), .A2(new_n643_), .ZN(new_n961_));
  AND3_X1   g760(.A1(new_n947_), .A2(G176gat), .A3(new_n658_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n949_), .A2(new_n658_), .ZN(new_n963_));
  AND2_X1   g762(.A1(new_n386_), .A2(new_n388_), .ZN(new_n964_));
  AOI22_X1  g763(.A1(new_n961_), .A2(new_n962_), .B1(new_n963_), .B2(new_n964_), .ZN(G1349gat));
  INV_X1    g764(.A(new_n949_), .ZN(new_n966_));
  NOR3_X1   g765(.A1(new_n966_), .A2(new_n443_), .A3(new_n659_), .ZN(new_n967_));
  NAND3_X1  g766(.A1(new_n961_), .A2(new_n360_), .A3(new_n947_), .ZN(new_n968_));
  AOI21_X1  g767(.A(new_n967_), .B1(new_n968_), .B2(new_n329_), .ZN(G1350gat));
  OAI21_X1  g768(.A(G190gat), .B1(new_n966_), .B2(new_n382_), .ZN(new_n970_));
  NAND3_X1  g769(.A1(new_n949_), .A2(new_n656_), .A3(new_n444_), .ZN(new_n971_));
  NAND2_X1  g770(.A1(new_n970_), .A2(new_n971_), .ZN(G1351gat));
  AND4_X1   g771(.A1(new_n649_), .A2(new_n897_), .A3(new_n694_), .A4(new_n725_), .ZN(new_n973_));
  NAND2_X1  g772(.A1(new_n973_), .A2(new_n240_), .ZN(new_n974_));
  XNOR2_X1  g773(.A(new_n974_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g774(.A1(new_n973_), .A2(new_n658_), .ZN(new_n976_));
  XOR2_X1   g775(.A(KEYINPUT126), .B(G204gat), .Z(new_n977_));
  XNOR2_X1  g776(.A(new_n976_), .B(new_n977_), .ZN(G1353gat));
  AOI21_X1  g777(.A(new_n659_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n979_));
  NAND2_X1  g778(.A1(new_n973_), .A2(new_n979_), .ZN(new_n980_));
  OR2_X1    g779(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n981_));
  XNOR2_X1  g780(.A(new_n980_), .B(new_n981_), .ZN(G1354gat));
  NAND2_X1  g781(.A1(new_n973_), .A2(new_n656_), .ZN(new_n983_));
  XOR2_X1   g782(.A(KEYINPUT127), .B(G218gat), .Z(new_n984_));
  NOR2_X1   g783(.A1(new_n382_), .A2(new_n984_), .ZN(new_n985_));
  AOI22_X1  g784(.A1(new_n983_), .A2(new_n984_), .B1(new_n973_), .B2(new_n985_), .ZN(G1355gat));
endmodule


