//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:32:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n671_, new_n672_, new_n673_, new_n675_, new_n676_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n725_, new_n726_, new_n728_, new_n729_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n852_, new_n853_, new_n854_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n863_, new_n865_,
    new_n866_, new_n868_, new_n869_, new_n870_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n886_,
    new_n887_, new_n888_, new_n890_, new_n891_, new_n892_, new_n894_,
    new_n895_, new_n897_, new_n898_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_;
  INV_X1    g000(.A(KEYINPUT105), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G113gat), .B(G141gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT82), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G169gat), .B(G197gat), .ZN(new_n205_));
  XOR2_X1   g004(.A(new_n204_), .B(new_n205_), .Z(new_n206_));
  XNOR2_X1  g005(.A(KEYINPUT77), .B(KEYINPUT78), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209_));
  XOR2_X1   g008(.A(KEYINPUT76), .B(G8gat), .Z(new_n210_));
  XNOR2_X1  g009(.A(KEYINPUT75), .B(G1gat), .ZN(new_n211_));
  AOI21_X1  g010(.A(new_n209_), .B1(new_n210_), .B2(new_n211_), .ZN(new_n212_));
  XNOR2_X1  g011(.A(G1gat), .B(G8gat), .ZN(new_n213_));
  XOR2_X1   g012(.A(G15gat), .B(G22gat), .Z(new_n214_));
  NOR3_X1   g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n213_), .ZN(new_n216_));
  XOR2_X1   g015(.A(KEYINPUT75), .B(G1gat), .Z(new_n217_));
  XNOR2_X1  g016(.A(KEYINPUT76), .B(G8gat), .ZN(new_n218_));
  OAI21_X1  g017(.A(KEYINPUT14), .B1(new_n217_), .B2(new_n218_), .ZN(new_n219_));
  INV_X1    g018(.A(new_n214_), .ZN(new_n220_));
  AOI21_X1  g019(.A(new_n216_), .B1(new_n219_), .B2(new_n220_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n208_), .B1(new_n215_), .B2(new_n221_), .ZN(new_n222_));
  OAI21_X1  g021(.A(new_n213_), .B1(new_n212_), .B2(new_n214_), .ZN(new_n223_));
  NAND3_X1  g022(.A1(new_n219_), .A2(new_n216_), .A3(new_n220_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n223_), .A2(new_n207_), .A3(new_n224_), .ZN(new_n225_));
  XOR2_X1   g024(.A(G29gat), .B(G36gat), .Z(new_n226_));
  XOR2_X1   g025(.A(G43gat), .B(G50gat), .Z(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  XNOR2_X1  g027(.A(G29gat), .B(G36gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G43gat), .B(G50gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n229_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n228_), .A2(new_n231_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n222_), .A2(new_n225_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234_));
  NAND2_X1  g033(.A1(new_n233_), .A2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(KEYINPUT15), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n232_), .A2(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n228_), .A2(KEYINPUT15), .A3(new_n231_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n237_), .A2(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(new_n239_), .ZN(new_n240_));
  AND3_X1   g039(.A1(new_n223_), .A2(new_n207_), .A3(new_n224_), .ZN(new_n241_));
  AOI21_X1  g040(.A(new_n207_), .B1(new_n223_), .B2(new_n224_), .ZN(new_n242_));
  OAI21_X1  g041(.A(new_n240_), .B1(new_n241_), .B2(new_n242_), .ZN(new_n243_));
  NAND2_X1  g042(.A1(new_n243_), .A2(KEYINPUT81), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n222_), .A2(new_n225_), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT81), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n245_), .A2(new_n246_), .A3(new_n240_), .ZN(new_n247_));
  AOI21_X1  g046(.A(new_n235_), .B1(new_n244_), .B2(new_n247_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n231_), .B(new_n228_), .C1(new_n241_), .C2(new_n242_), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n234_), .B1(new_n249_), .B2(new_n233_), .ZN(new_n250_));
  OAI21_X1  g049(.A(new_n206_), .B1(new_n248_), .B2(new_n250_), .ZN(new_n251_));
  AND2_X1   g050(.A1(new_n233_), .A2(new_n234_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n246_), .B1(new_n245_), .B2(new_n240_), .ZN(new_n253_));
  AOI211_X1 g052(.A(KEYINPUT81), .B(new_n239_), .C1(new_n222_), .C2(new_n225_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n252_), .B1(new_n253_), .B2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n250_), .ZN(new_n256_));
  INV_X1    g055(.A(new_n206_), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n255_), .A2(new_n256_), .A3(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT83), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n251_), .A2(new_n258_), .A3(new_n259_), .ZN(new_n260_));
  OAI211_X1 g059(.A(KEYINPUT83), .B(new_n206_), .C1(new_n248_), .C2(new_n250_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  NAND2_X1  g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263_));
  INV_X1    g062(.A(KEYINPUT23), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n263_), .B(new_n264_), .ZN(new_n265_));
  NOR2_X1   g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266_));
  INV_X1    g065(.A(KEYINPUT84), .ZN(new_n267_));
  XNOR2_X1  g066(.A(new_n266_), .B(new_n267_), .ZN(new_n268_));
  INV_X1    g067(.A(KEYINPUT24), .ZN(new_n269_));
  AOI21_X1  g068(.A(new_n265_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  XNOR2_X1  g069(.A(KEYINPUT25), .B(G183gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(KEYINPUT26), .B(G190gat), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n266_), .B(KEYINPUT84), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n269_), .B1(G169gat), .B2(G176gat), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n274_), .A2(new_n275_), .ZN(new_n276_));
  NAND3_X1  g075(.A1(new_n270_), .A2(new_n273_), .A3(new_n276_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n278_), .B1(new_n264_), .B2(new_n263_), .ZN(new_n279_));
  OAI21_X1  g078(.A(new_n279_), .B1(new_n264_), .B2(new_n263_), .ZN(new_n280_));
  OAI21_X1  g079(.A(G169gat), .B1(KEYINPUT22), .B2(G176gat), .ZN(new_n281_));
  OR3_X1    g080(.A1(KEYINPUT22), .A2(G169gat), .A3(G176gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n280_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n277_), .A2(new_n283_), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT85), .ZN(new_n285_));
  NAND2_X1  g084(.A1(new_n284_), .A2(new_n285_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n277_), .A2(KEYINPUT85), .A3(new_n283_), .ZN(new_n287_));
  AND2_X1   g086(.A1(new_n286_), .A2(new_n287_), .ZN(new_n288_));
  XNOR2_X1  g087(.A(new_n288_), .B(KEYINPUT30), .ZN(new_n289_));
  NAND2_X1  g088(.A1(new_n289_), .A2(KEYINPUT88), .ZN(new_n290_));
  XNOR2_X1  g089(.A(new_n289_), .B(KEYINPUT88), .ZN(new_n291_));
  XOR2_X1   g090(.A(G71gat), .B(G99gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(KEYINPUT86), .B(G43gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(new_n292_), .B(new_n293_), .ZN(new_n294_));
  XOR2_X1   g093(.A(KEYINPUT87), .B(G15gat), .Z(new_n295_));
  NAND2_X1  g094(.A1(G227gat), .A2(G233gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n294_), .B(new_n297_), .ZN(new_n298_));
  MUX2_X1   g097(.A(new_n290_), .B(new_n291_), .S(new_n298_), .Z(new_n299_));
  XNOR2_X1  g098(.A(G127gat), .B(G134gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n300_), .B(KEYINPUT89), .ZN(new_n301_));
  XNOR2_X1  g100(.A(G113gat), .B(G120gat), .ZN(new_n302_));
  XNOR2_X1  g101(.A(new_n301_), .B(new_n302_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n303_), .B(KEYINPUT31), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n299_), .B(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(new_n305_), .ZN(new_n306_));
  XOR2_X1   g105(.A(G155gat), .B(G162gat), .Z(new_n307_));
  NAND3_X1  g106(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n308_), .B(KEYINPUT90), .ZN(new_n309_));
  INV_X1    g108(.A(KEYINPUT3), .ZN(new_n310_));
  INV_X1    g109(.A(G141gat), .ZN(new_n311_));
  INV_X1    g110(.A(G148gat), .ZN(new_n312_));
  NAND3_X1  g111(.A1(new_n310_), .A2(new_n311_), .A3(new_n312_), .ZN(new_n313_));
  OAI21_X1  g112(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n314_));
  NOR2_X1   g113(.A1(new_n311_), .A2(new_n312_), .ZN(new_n315_));
  OAI211_X1 g114(.A(new_n313_), .B(new_n314_), .C1(new_n315_), .C2(KEYINPUT2), .ZN(new_n316_));
  OAI21_X1  g115(.A(new_n307_), .B1(new_n309_), .B2(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n317_), .A2(KEYINPUT91), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT1), .ZN(new_n319_));
  NAND2_X1  g118(.A1(new_n307_), .A2(new_n319_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n311_), .A2(new_n312_), .ZN(new_n321_));
  INV_X1    g120(.A(new_n315_), .ZN(new_n322_));
  NAND3_X1  g121(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n320_), .A2(new_n321_), .A3(new_n322_), .A4(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n318_), .A2(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n317_), .A2(KEYINPUT91), .ZN(new_n326_));
  OR2_X1    g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n327_), .A2(KEYINPUT29), .ZN(new_n328_));
  XOR2_X1   g127(.A(G197gat), .B(G204gat), .Z(new_n329_));
  OR2_X1    g128(.A1(new_n329_), .A2(KEYINPUT21), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(KEYINPUT21), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G211gat), .B(G218gat), .ZN(new_n332_));
  NAND3_X1  g131(.A1(new_n330_), .A2(new_n331_), .A3(new_n332_), .ZN(new_n333_));
  OR2_X1    g132(.A1(new_n331_), .A2(new_n332_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n333_), .A2(new_n334_), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n328_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(G228gat), .A2(G233gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n337_), .B1(new_n335_), .B2(KEYINPUT93), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  OAI211_X1 g138(.A(new_n328_), .B(new_n335_), .C1(KEYINPUT93), .C2(new_n337_), .ZN(new_n340_));
  XNOR2_X1  g139(.A(G78gat), .B(G106gat), .ZN(new_n341_));
  XOR2_X1   g140(.A(new_n341_), .B(KEYINPUT94), .Z(new_n342_));
  NAND3_X1  g141(.A1(new_n339_), .A2(new_n340_), .A3(new_n342_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(new_n325_), .A2(new_n326_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT29), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n344_), .A2(new_n345_), .ZN(new_n346_));
  XOR2_X1   g145(.A(KEYINPUT92), .B(KEYINPUT28), .Z(new_n347_));
  OR2_X1    g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n346_), .A2(new_n347_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  XOR2_X1   g149(.A(G22gat), .B(G50gat), .Z(new_n351_));
  INV_X1    g150(.A(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n350_), .A2(new_n352_), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n349_), .A2(new_n351_), .A3(new_n348_), .ZN(new_n354_));
  NAND3_X1  g153(.A1(new_n343_), .A2(new_n353_), .A3(new_n354_), .ZN(new_n355_));
  NAND3_X1  g154(.A1(new_n339_), .A2(KEYINPUT95), .A3(new_n340_), .ZN(new_n356_));
  INV_X1    g155(.A(new_n341_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n339_), .A2(new_n340_), .ZN(new_n358_));
  INV_X1    g157(.A(KEYINPUT95), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n357_), .B1(new_n358_), .B2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n355_), .B1(new_n356_), .B2(new_n360_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n342_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n358_), .A2(new_n362_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n363_), .A2(new_n343_), .B1(new_n354_), .B2(new_n353_), .ZN(new_n364_));
  NOR2_X1   g163(.A1(new_n361_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(new_n365_), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n367_), .B(KEYINPUT19), .ZN(new_n368_));
  INV_X1    g167(.A(new_n335_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n286_), .A2(new_n369_), .A3(new_n287_), .ZN(new_n370_));
  INV_X1    g169(.A(KEYINPUT96), .ZN(new_n371_));
  NAND3_X1  g170(.A1(new_n370_), .A2(new_n371_), .A3(KEYINPUT20), .ZN(new_n372_));
  NOR3_X1   g171(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n373_));
  OAI21_X1  g172(.A(KEYINPUT97), .B1(new_n265_), .B2(new_n373_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n374_), .A2(new_n276_), .A3(new_n273_), .ZN(new_n375_));
  NOR3_X1   g174(.A1(new_n265_), .A2(KEYINPUT97), .A3(new_n373_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n283_), .B1(new_n375_), .B2(new_n376_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n377_), .A2(new_n335_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(new_n372_), .A2(new_n378_), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n371_), .B1(new_n370_), .B2(KEYINPUT20), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n368_), .B1(new_n379_), .B2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n288_), .A2(new_n369_), .ZN(new_n382_));
  OAI21_X1  g181(.A(KEYINPUT20), .B1(new_n377_), .B2(new_n335_), .ZN(new_n383_));
  OR3_X1    g182(.A1(new_n382_), .A2(new_n368_), .A3(new_n383_), .ZN(new_n384_));
  XOR2_X1   g183(.A(G8gat), .B(G36gat), .Z(new_n385_));
  XNOR2_X1  g184(.A(KEYINPUT98), .B(KEYINPUT18), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n385_), .B(new_n386_), .ZN(new_n387_));
  XNOR2_X1  g186(.A(G64gat), .B(G92gat), .ZN(new_n388_));
  XNOR2_X1  g187(.A(new_n387_), .B(new_n388_), .ZN(new_n389_));
  NAND2_X1  g188(.A1(new_n389_), .A2(KEYINPUT32), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n381_), .A2(new_n384_), .A3(new_n390_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n391_), .A2(KEYINPUT100), .ZN(new_n392_));
  INV_X1    g191(.A(KEYINPUT100), .ZN(new_n393_));
  NAND4_X1  g192(.A1(new_n381_), .A2(new_n384_), .A3(new_n393_), .A4(new_n390_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n392_), .A2(new_n394_), .ZN(new_n395_));
  INV_X1    g194(.A(new_n303_), .ZN(new_n396_));
  NAND2_X1  g195(.A1(new_n327_), .A2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(new_n344_), .A2(new_n303_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n397_), .A2(KEYINPUT4), .A3(new_n398_), .ZN(new_n399_));
  INV_X1    g198(.A(KEYINPUT99), .ZN(new_n400_));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OR3_X1    g201(.A1(new_n344_), .A2(KEYINPUT4), .A3(new_n303_), .ZN(new_n403_));
  NAND4_X1  g202(.A1(new_n399_), .A2(new_n400_), .A3(new_n402_), .A4(new_n403_), .ZN(new_n404_));
  AND3_X1   g203(.A1(new_n399_), .A2(new_n402_), .A3(new_n403_), .ZN(new_n405_));
  NAND3_X1  g204(.A1(new_n397_), .A2(new_n401_), .A3(new_n398_), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n406_), .A2(KEYINPUT99), .ZN(new_n407_));
  OAI21_X1  g206(.A(new_n404_), .B1(new_n405_), .B2(new_n407_), .ZN(new_n408_));
  XNOR2_X1  g207(.A(G1gat), .B(G29gat), .ZN(new_n409_));
  XNOR2_X1  g208(.A(new_n409_), .B(G85gat), .ZN(new_n410_));
  XNOR2_X1  g209(.A(KEYINPUT0), .B(G57gat), .ZN(new_n411_));
  XOR2_X1   g210(.A(new_n410_), .B(new_n411_), .Z(new_n412_));
  NAND2_X1  g211(.A1(new_n408_), .A2(new_n412_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n412_), .ZN(new_n414_));
  OAI211_X1 g213(.A(new_n414_), .B(new_n404_), .C1(new_n405_), .C2(new_n407_), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n413_), .A2(new_n415_), .ZN(new_n416_));
  OAI21_X1  g215(.A(new_n368_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n417_));
  NAND2_X1  g216(.A1(new_n370_), .A2(KEYINPUT20), .ZN(new_n418_));
  NAND2_X1  g217(.A1(new_n418_), .A2(KEYINPUT96), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n419_), .A2(new_n378_), .A3(new_n372_), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n417_), .B1(new_n420_), .B2(new_n368_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n421_), .A2(KEYINPUT32), .A3(new_n389_), .ZN(new_n422_));
  NAND3_X1  g221(.A1(new_n395_), .A2(new_n416_), .A3(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT101), .ZN(new_n424_));
  AND3_X1   g223(.A1(new_n408_), .A2(KEYINPUT33), .A3(new_n412_), .ZN(new_n425_));
  AOI21_X1  g224(.A(KEYINPUT33), .B1(new_n408_), .B2(new_n412_), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  AND3_X1   g226(.A1(new_n381_), .A2(new_n384_), .A3(new_n389_), .ZN(new_n428_));
  AOI21_X1  g227(.A(new_n389_), .B1(new_n381_), .B2(new_n384_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n399_), .A2(new_n401_), .A3(new_n403_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n397_), .A2(new_n402_), .A3(new_n398_), .ZN(new_n431_));
  AND3_X1   g230(.A1(new_n430_), .A2(new_n414_), .A3(new_n431_), .ZN(new_n432_));
  NOR3_X1   g231(.A1(new_n428_), .A2(new_n429_), .A3(new_n432_), .ZN(new_n433_));
  AOI22_X1  g232(.A1(new_n423_), .A2(new_n424_), .B1(new_n427_), .B2(new_n433_), .ZN(new_n434_));
  NAND4_X1  g233(.A1(new_n395_), .A2(new_n416_), .A3(KEYINPUT101), .A4(new_n422_), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n366_), .B1(new_n434_), .B2(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(KEYINPUT27), .ZN(new_n437_));
  OAI21_X1  g236(.A(new_n437_), .B1(new_n428_), .B2(new_n429_), .ZN(new_n438_));
  NAND2_X1  g237(.A1(new_n438_), .A2(KEYINPUT103), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT103), .ZN(new_n440_));
  OAI211_X1 g239(.A(new_n440_), .B(new_n437_), .C1(new_n428_), .C2(new_n429_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n389_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n421_), .A2(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT102), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n443_), .A2(new_n444_), .ZN(new_n445_));
  NAND3_X1  g244(.A1(new_n421_), .A2(KEYINPUT102), .A3(new_n442_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n428_), .A2(new_n437_), .ZN(new_n448_));
  AOI22_X1  g247(.A1(new_n439_), .A2(new_n441_), .B1(new_n447_), .B2(new_n448_), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n365_), .A2(new_n416_), .ZN(new_n450_));
  AND2_X1   g249(.A1(new_n449_), .A2(new_n450_), .ZN(new_n451_));
  OAI21_X1  g250(.A(new_n306_), .B1(new_n436_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n416_), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n305_), .A2(new_n453_), .A3(new_n365_), .A4(new_n449_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n262_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT37), .ZN(new_n456_));
  INV_X1    g255(.A(G85gat), .ZN(new_n457_));
  INV_X1    g256(.A(G92gat), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n457_), .A2(new_n458_), .ZN(new_n459_));
  NAND2_X1  g258(.A1(G85gat), .A2(G92gat), .ZN(new_n460_));
  INV_X1    g259(.A(KEYINPUT9), .ZN(new_n461_));
  AOI22_X1  g260(.A1(new_n459_), .A2(new_n460_), .B1(new_n461_), .B2(G92gat), .ZN(new_n462_));
  INV_X1    g261(.A(new_n462_), .ZN(new_n463_));
  INV_X1    g262(.A(KEYINPUT64), .ZN(new_n464_));
  NAND3_X1  g263(.A1(new_n459_), .A2(new_n461_), .A3(new_n460_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n463_), .A2(new_n464_), .A3(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(new_n465_), .ZN(new_n467_));
  OAI21_X1  g266(.A(KEYINPUT64), .B1(new_n467_), .B2(new_n462_), .ZN(new_n468_));
  XOR2_X1   g267(.A(KEYINPUT10), .B(G99gat), .Z(new_n469_));
  INV_X1    g268(.A(G106gat), .ZN(new_n470_));
  NAND2_X1  g269(.A1(G99gat), .A2(G106gat), .ZN(new_n471_));
  NAND2_X1  g270(.A1(new_n471_), .A2(KEYINPUT6), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n473_), .A2(G99gat), .A3(G106gat), .ZN(new_n474_));
  AOI22_X1  g273(.A1(new_n469_), .A2(new_n470_), .B1(new_n472_), .B2(new_n474_), .ZN(new_n475_));
  NAND3_X1  g274(.A1(new_n466_), .A2(new_n468_), .A3(new_n475_), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT8), .ZN(new_n477_));
  AOI21_X1  g276(.A(new_n473_), .B1(G99gat), .B2(G106gat), .ZN(new_n478_));
  NOR2_X1   g277(.A1(new_n471_), .A2(KEYINPUT6), .ZN(new_n479_));
  OAI21_X1  g278(.A(KEYINPUT65), .B1(new_n478_), .B2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT65), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n472_), .A2(new_n474_), .A3(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(KEYINPUT7), .ZN(new_n483_));
  INV_X1    g282(.A(G99gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n483_), .A2(new_n484_), .A3(new_n470_), .ZN(new_n485_));
  OAI21_X1  g284(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n486_));
  AND2_X1   g285(.A1(new_n485_), .A2(new_n486_), .ZN(new_n487_));
  NAND3_X1  g286(.A1(new_n480_), .A2(new_n482_), .A3(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n459_), .A2(new_n460_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n489_), .ZN(new_n490_));
  AOI21_X1  g289(.A(new_n477_), .B1(new_n488_), .B2(new_n490_), .ZN(new_n491_));
  NAND2_X1  g290(.A1(new_n472_), .A2(new_n474_), .ZN(new_n492_));
  AOI211_X1 g291(.A(KEYINPUT8), .B(new_n489_), .C1(new_n487_), .C2(new_n492_), .ZN(new_n493_));
  OAI211_X1 g292(.A(new_n232_), .B(new_n476_), .C1(new_n491_), .C2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT70), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(G232gat), .A2(G233gat), .ZN(new_n497_));
  XOR2_X1   g296(.A(new_n497_), .B(KEYINPUT34), .Z(new_n498_));
  INV_X1    g297(.A(KEYINPUT35), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XOR2_X1   g299(.A(new_n500_), .B(KEYINPUT71), .Z(new_n501_));
  OAI21_X1  g300(.A(new_n476_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n501_), .B1(new_n502_), .B2(new_n240_), .ZN(new_n503_));
  NAND2_X1  g302(.A1(new_n496_), .A2(new_n503_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n504_), .A2(KEYINPUT69), .ZN(new_n505_));
  INV_X1    g304(.A(KEYINPUT69), .ZN(new_n506_));
  NAND3_X1  g305(.A1(new_n496_), .A2(new_n506_), .A3(new_n503_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n505_), .A2(new_n507_), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n498_), .A2(new_n499_), .ZN(new_n509_));
  INV_X1    g308(.A(new_n509_), .ZN(new_n510_));
  NAND2_X1  g309(.A1(new_n508_), .A2(new_n510_), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n505_), .A2(new_n509_), .A3(new_n507_), .ZN(new_n512_));
  XOR2_X1   g311(.A(G190gat), .B(G218gat), .Z(new_n513_));
  XNOR2_X1  g312(.A(new_n513_), .B(KEYINPUT72), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G134gat), .B(G162gat), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n514_), .B(new_n515_), .ZN(new_n516_));
  INV_X1    g315(.A(KEYINPUT36), .ZN(new_n517_));
  XNOR2_X1  g316(.A(new_n516_), .B(new_n517_), .ZN(new_n518_));
  XNOR2_X1  g317(.A(new_n518_), .B(KEYINPUT74), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n511_), .A2(new_n512_), .A3(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n516_), .A2(new_n517_), .ZN(new_n522_));
  XNOR2_X1  g321(.A(new_n522_), .B(KEYINPUT73), .ZN(new_n523_));
  INV_X1    g322(.A(new_n523_), .ZN(new_n524_));
  AOI21_X1  g323(.A(new_n524_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n525_));
  OAI21_X1  g324(.A(new_n456_), .B1(new_n521_), .B2(new_n525_), .ZN(new_n526_));
  AND2_X1   g325(.A1(new_n511_), .A2(new_n512_), .ZN(new_n527_));
  OAI211_X1 g326(.A(KEYINPUT37), .B(new_n520_), .C1(new_n527_), .C2(new_n524_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n526_), .A2(new_n528_), .ZN(new_n529_));
  XNOR2_X1  g328(.A(G120gat), .B(G148gat), .ZN(new_n530_));
  XNOR2_X1  g329(.A(new_n530_), .B(KEYINPUT5), .ZN(new_n531_));
  XNOR2_X1  g330(.A(G176gat), .B(G204gat), .ZN(new_n532_));
  XOR2_X1   g331(.A(new_n531_), .B(new_n532_), .Z(new_n533_));
  INV_X1    g332(.A(KEYINPUT66), .ZN(new_n534_));
  XNOR2_X1  g333(.A(G57gat), .B(G64gat), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n536_));
  XOR2_X1   g335(.A(G71gat), .B(G78gat), .Z(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  NOR2_X1   g337(.A1(new_n535_), .A2(KEYINPUT11), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n536_), .A2(new_n537_), .ZN(new_n540_));
  OAI21_X1  g339(.A(new_n538_), .B1(new_n539_), .B2(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n487_), .A2(new_n492_), .ZN(new_n542_));
  NAND3_X1  g341(.A1(new_n542_), .A2(new_n477_), .A3(new_n490_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n485_), .A2(new_n486_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n544_), .B1(KEYINPUT65), .B2(new_n492_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n489_), .B1(new_n545_), .B2(new_n482_), .ZN(new_n546_));
  OAI21_X1  g345(.A(new_n543_), .B1(new_n546_), .B2(new_n477_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n541_), .B1(new_n547_), .B2(new_n476_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n476_), .B(new_n541_), .C1(new_n491_), .C2(new_n493_), .ZN(new_n549_));
  INV_X1    g348(.A(new_n549_), .ZN(new_n550_));
  NOR2_X1   g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G230gat), .A2(G233gat), .ZN(new_n552_));
  OAI21_X1  g351(.A(new_n534_), .B1(new_n551_), .B2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n552_), .ZN(new_n554_));
  OAI211_X1 g353(.A(KEYINPUT66), .B(new_n554_), .C1(new_n548_), .C2(new_n550_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n553_), .A2(new_n555_), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT67), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT12), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  OAI21_X1  g358(.A(new_n559_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n560_));
  INV_X1    g359(.A(new_n541_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n502_), .A2(new_n561_), .ZN(new_n562_));
  NOR2_X1   g361(.A1(new_n557_), .A2(KEYINPUT12), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n558_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND3_X1  g363(.A1(new_n560_), .A2(new_n552_), .A3(new_n564_), .ZN(new_n565_));
  INV_X1    g364(.A(new_n565_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n533_), .B1(new_n556_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n533_), .ZN(new_n568_));
  NAND4_X1  g367(.A1(new_n565_), .A2(new_n553_), .A3(new_n555_), .A4(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n567_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT68), .ZN(new_n571_));
  OAI21_X1  g370(.A(new_n570_), .B1(new_n571_), .B2(KEYINPUT13), .ZN(new_n572_));
  XNOR2_X1  g371(.A(KEYINPUT68), .B(KEYINPUT13), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n572_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  INV_X1    g373(.A(new_n574_), .ZN(new_n575_));
  XOR2_X1   g374(.A(G127gat), .B(G155gat), .Z(new_n576_));
  XNOR2_X1  g375(.A(G183gat), .B(G211gat), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n576_), .B(new_n577_), .ZN(new_n578_));
  XOR2_X1   g377(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n579_));
  XNOR2_X1  g378(.A(new_n578_), .B(new_n579_), .ZN(new_n580_));
  INV_X1    g379(.A(KEYINPUT17), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n580_), .A2(new_n581_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n541_), .B(new_n583_), .ZN(new_n584_));
  XNOR2_X1  g383(.A(new_n584_), .B(new_n245_), .ZN(new_n585_));
  NAND2_X1  g384(.A1(new_n585_), .A2(new_n581_), .ZN(new_n586_));
  INV_X1    g385(.A(new_n586_), .ZN(new_n587_));
  OAI21_X1  g386(.A(new_n582_), .B1(new_n587_), .B2(new_n580_), .ZN(new_n588_));
  INV_X1    g387(.A(KEYINPUT80), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n588_), .A2(new_n589_), .A3(new_n585_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n585_), .A2(new_n589_), .ZN(new_n591_));
  OAI211_X1 g390(.A(new_n591_), .B(new_n582_), .C1(new_n587_), .C2(new_n580_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n590_), .A2(new_n592_), .ZN(new_n593_));
  NOR3_X1   g392(.A1(new_n529_), .A2(new_n575_), .A3(new_n593_), .ZN(new_n594_));
  NAND2_X1  g393(.A1(new_n455_), .A2(new_n594_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n595_), .A2(KEYINPUT104), .ZN(new_n596_));
  INV_X1    g395(.A(new_n596_), .ZN(new_n597_));
  NOR2_X1   g396(.A1(new_n595_), .A2(KEYINPUT104), .ZN(new_n598_));
  OAI21_X1  g397(.A(new_n202_), .B1(new_n597_), .B2(new_n598_), .ZN(new_n599_));
  OR2_X1    g398(.A1(new_n595_), .A2(KEYINPUT104), .ZN(new_n600_));
  NAND3_X1  g399(.A1(new_n600_), .A2(KEYINPUT105), .A3(new_n596_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n453_), .A2(new_n211_), .ZN(new_n602_));
  NAND3_X1  g401(.A1(new_n599_), .A2(new_n601_), .A3(new_n602_), .ZN(new_n603_));
  INV_X1    g402(.A(KEYINPUT38), .ZN(new_n604_));
  OR2_X1    g403(.A1(new_n603_), .A2(new_n604_), .ZN(new_n605_));
  NOR2_X1   g404(.A1(new_n521_), .A2(new_n525_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT106), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n607_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n262_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n574_), .A2(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n610_), .A2(new_n593_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(G1gat), .B1(new_n613_), .B2(new_n453_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n603_), .A2(new_n604_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n605_), .A2(new_n614_), .A3(new_n615_), .ZN(G1324gat));
  INV_X1    g415(.A(new_n449_), .ZN(new_n617_));
  NAND4_X1  g416(.A1(new_n599_), .A2(new_n601_), .A3(new_n617_), .A4(new_n218_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n608_), .A2(new_n617_), .A3(new_n611_), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n619_), .A2(G8gat), .ZN(new_n620_));
  XNOR2_X1  g419(.A(new_n620_), .B(KEYINPUT39), .ZN(new_n621_));
  NAND2_X1  g420(.A1(new_n618_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT40), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n622_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n618_), .A2(KEYINPUT40), .A3(new_n621_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(G1325gat));
  INV_X1    g425(.A(G15gat), .ZN(new_n627_));
  AOI21_X1  g426(.A(new_n627_), .B1(new_n612_), .B2(new_n305_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT41), .ZN(new_n629_));
  NOR2_X1   g428(.A1(new_n597_), .A2(new_n598_), .ZN(new_n630_));
  NAND3_X1  g429(.A1(new_n630_), .A2(new_n627_), .A3(new_n305_), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n629_), .A2(new_n631_), .ZN(G1326gat));
  INV_X1    g431(.A(G22gat), .ZN(new_n633_));
  AOI21_X1  g432(.A(new_n633_), .B1(new_n612_), .B2(new_n366_), .ZN(new_n634_));
  XOR2_X1   g433(.A(new_n634_), .B(KEYINPUT42), .Z(new_n635_));
  NAND3_X1  g434(.A1(new_n630_), .A2(new_n633_), .A3(new_n366_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n635_), .A2(new_n636_), .ZN(G1327gat));
  INV_X1    g436(.A(new_n606_), .ZN(new_n638_));
  INV_X1    g437(.A(new_n593_), .ZN(new_n639_));
  NOR3_X1   g438(.A1(new_n575_), .A2(new_n638_), .A3(new_n639_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n455_), .A2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  AOI21_X1  g441(.A(G29gat), .B1(new_n642_), .B2(new_n416_), .ZN(new_n643_));
  NOR2_X1   g442(.A1(new_n610_), .A2(new_n639_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n529_), .ZN(new_n645_));
  AOI211_X1 g444(.A(KEYINPUT43), .B(new_n645_), .C1(new_n452_), .C2(new_n454_), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT43), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n423_), .A2(new_n424_), .ZN(new_n648_));
  NAND2_X1  g447(.A1(new_n427_), .A2(new_n433_), .ZN(new_n649_));
  NAND3_X1  g448(.A1(new_n648_), .A2(new_n435_), .A3(new_n649_), .ZN(new_n650_));
  AOI22_X1  g449(.A1(new_n650_), .A2(new_n365_), .B1(new_n450_), .B2(new_n449_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n454_), .B1(new_n651_), .B2(new_n305_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n647_), .B1(new_n652_), .B2(new_n529_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n644_), .B1(new_n646_), .B2(new_n653_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  OAI211_X1 g455(.A(KEYINPUT44), .B(new_n644_), .C1(new_n646_), .C2(new_n653_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  AND2_X1   g457(.A1(new_n416_), .A2(G29gat), .ZN(new_n659_));
  AOI21_X1  g458(.A(new_n643_), .B1(new_n658_), .B2(new_n659_), .ZN(G1328gat));
  NAND3_X1  g459(.A1(new_n656_), .A2(new_n617_), .A3(new_n657_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(G36gat), .ZN(new_n662_));
  NOR3_X1   g461(.A1(new_n641_), .A2(G36gat), .A3(new_n449_), .ZN(new_n663_));
  INV_X1    g462(.A(KEYINPUT45), .ZN(new_n664_));
  XNOR2_X1  g463(.A(new_n663_), .B(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n662_), .A2(new_n665_), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT46), .ZN(new_n667_));
  NAND2_X1  g466(.A1(new_n666_), .A2(new_n667_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n662_), .A2(new_n665_), .A3(KEYINPUT46), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n668_), .A2(new_n669_), .ZN(G1329gat));
  NAND4_X1  g469(.A1(new_n656_), .A2(G43gat), .A3(new_n305_), .A4(new_n657_), .ZN(new_n671_));
  NOR2_X1   g470(.A1(new_n641_), .A2(new_n306_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(G43gat), .B2(new_n672_), .ZN(new_n673_));
  XNOR2_X1  g472(.A(new_n673_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g473(.A(G50gat), .B1(new_n642_), .B2(new_n366_), .ZN(new_n675_));
  AND2_X1   g474(.A1(new_n366_), .A2(G50gat), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n675_), .B1(new_n658_), .B2(new_n676_), .ZN(G1331gat));
  INV_X1    g476(.A(G57gat), .ZN(new_n678_));
  AOI21_X1  g477(.A(new_n609_), .B1(new_n452_), .B2(new_n454_), .ZN(new_n679_));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n679_), .B(new_n680_), .ZN(new_n681_));
  NOR2_X1   g480(.A1(new_n574_), .A2(new_n593_), .ZN(new_n682_));
  INV_X1    g481(.A(new_n682_), .ZN(new_n683_));
  NOR2_X1   g482(.A1(new_n683_), .A2(new_n529_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n684_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n678_), .B1(new_n685_), .B2(new_n453_), .ZN(new_n686_));
  OR2_X1    g485(.A1(new_n686_), .A2(KEYINPUT108), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n686_), .A2(KEYINPUT108), .ZN(new_n688_));
  INV_X1    g487(.A(new_n607_), .ZN(new_n689_));
  AND4_X1   g488(.A1(new_n652_), .A2(new_n262_), .A3(new_n689_), .A4(new_n682_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(KEYINPUT109), .B(G57gat), .ZN(new_n691_));
  NOR2_X1   g490(.A1(new_n453_), .A2(new_n691_), .ZN(new_n692_));
  AOI22_X1  g491(.A1(new_n687_), .A2(new_n688_), .B1(new_n690_), .B2(new_n692_), .ZN(G1332gat));
  INV_X1    g492(.A(G64gat), .ZN(new_n694_));
  AOI21_X1  g493(.A(new_n694_), .B1(new_n690_), .B2(new_n617_), .ZN(new_n695_));
  XOR2_X1   g494(.A(new_n695_), .B(KEYINPUT48), .Z(new_n696_));
  NAND2_X1  g495(.A1(new_n617_), .A2(new_n694_), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n696_), .B1(new_n685_), .B2(new_n697_), .ZN(G1333gat));
  NAND2_X1  g497(.A1(new_n690_), .A2(new_n305_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n699_), .A2(G71gat), .ZN(new_n700_));
  OR2_X1    g499(.A1(new_n700_), .A2(KEYINPUT110), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(KEYINPUT110), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n701_), .A2(new_n702_), .ZN(new_n703_));
  INV_X1    g502(.A(KEYINPUT49), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n703_), .A2(new_n704_), .ZN(new_n705_));
  OR3_X1    g504(.A1(new_n685_), .A2(G71gat), .A3(new_n306_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n701_), .A2(KEYINPUT49), .A3(new_n702_), .ZN(new_n707_));
  NAND3_X1  g506(.A1(new_n705_), .A2(new_n706_), .A3(new_n707_), .ZN(G1334gat));
  INV_X1    g507(.A(KEYINPUT50), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n690_), .A2(new_n366_), .ZN(new_n710_));
  AOI21_X1  g509(.A(new_n709_), .B1(new_n710_), .B2(G78gat), .ZN(new_n711_));
  INV_X1    g510(.A(G78gat), .ZN(new_n712_));
  AOI211_X1 g511(.A(KEYINPUT50), .B(new_n712_), .C1(new_n690_), .C2(new_n366_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n366_), .A2(new_n712_), .ZN(new_n714_));
  OAI22_X1  g513(.A1(new_n711_), .A2(new_n713_), .B1(new_n685_), .B2(new_n714_), .ZN(new_n715_));
  XOR2_X1   g514(.A(new_n715_), .B(KEYINPUT111), .Z(G1335gat));
  NOR2_X1   g515(.A1(new_n646_), .A2(new_n653_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n575_), .A2(new_n593_), .ZN(new_n718_));
  NOR3_X1   g517(.A1(new_n717_), .A2(new_n609_), .A3(new_n718_), .ZN(new_n719_));
  AOI21_X1  g518(.A(new_n457_), .B1(new_n719_), .B2(new_n416_), .ZN(new_n720_));
  NOR2_X1   g519(.A1(new_n718_), .A2(new_n638_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n681_), .A2(new_n721_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n722_), .A2(G85gat), .A3(new_n453_), .ZN(new_n723_));
  OR2_X1    g522(.A1(new_n720_), .A2(new_n723_), .ZN(G1336gat));
  AOI21_X1  g523(.A(new_n458_), .B1(new_n719_), .B2(new_n617_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n722_), .A2(G92gat), .A3(new_n449_), .ZN(new_n726_));
  OR2_X1    g525(.A1(new_n725_), .A2(new_n726_), .ZN(G1337gat));
  NOR2_X1   g526(.A1(new_n718_), .A2(new_n609_), .ZN(new_n728_));
  OAI211_X1 g527(.A(new_n305_), .B(new_n728_), .C1(new_n646_), .C2(new_n653_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT112), .ZN(new_n730_));
  AND3_X1   g529(.A1(new_n729_), .A2(new_n730_), .A3(G99gat), .ZN(new_n731_));
  AOI21_X1  g530(.A(new_n730_), .B1(new_n729_), .B2(G99gat), .ZN(new_n732_));
  NAND2_X1  g531(.A1(new_n305_), .A2(new_n469_), .ZN(new_n733_));
  OAI22_X1  g532(.A1(new_n731_), .A2(new_n732_), .B1(new_n722_), .B2(new_n733_), .ZN(new_n734_));
  XNOR2_X1  g533(.A(new_n734_), .B(KEYINPUT51), .ZN(G1338gat));
  OAI211_X1 g534(.A(new_n366_), .B(new_n728_), .C1(new_n646_), .C2(new_n653_), .ZN(new_n736_));
  AND3_X1   g535(.A1(new_n736_), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n737_));
  AOI21_X1  g536(.A(KEYINPUT113), .B1(new_n736_), .B2(G106gat), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n737_), .A2(new_n738_), .A3(new_n739_), .ZN(new_n740_));
  NAND2_X1  g539(.A1(new_n736_), .A2(G106gat), .ZN(new_n741_));
  INV_X1    g540(.A(KEYINPUT113), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n741_), .A2(new_n742_), .A3(new_n739_), .ZN(new_n743_));
  NAND4_X1  g542(.A1(new_n681_), .A2(new_n470_), .A3(new_n366_), .A4(new_n721_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n743_), .A2(new_n744_), .ZN(new_n745_));
  OAI21_X1  g544(.A(KEYINPUT53), .B1(new_n740_), .B2(new_n745_), .ZN(new_n746_));
  INV_X1    g545(.A(new_n738_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n736_), .A2(KEYINPUT113), .A3(G106gat), .ZN(new_n748_));
  NAND3_X1  g547(.A1(new_n747_), .A2(KEYINPUT52), .A3(new_n748_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT53), .ZN(new_n750_));
  NAND4_X1  g549(.A1(new_n749_), .A2(new_n750_), .A3(new_n743_), .A4(new_n744_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n746_), .A2(new_n751_), .ZN(G1339gat));
  AOI21_X1  g551(.A(new_n552_), .B1(new_n560_), .B2(new_n564_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT55), .ZN(new_n754_));
  OAI21_X1  g553(.A(new_n565_), .B1(new_n753_), .B2(new_n754_), .ZN(new_n755_));
  NAND4_X1  g554(.A1(new_n560_), .A2(new_n564_), .A3(KEYINPUT55), .A4(new_n552_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n755_), .A2(new_n756_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n757_), .A2(KEYINPUT115), .A3(new_n533_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT116), .ZN(new_n759_));
  AOI21_X1  g558(.A(KEYINPUT56), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n568_), .B1(new_n755_), .B2(new_n756_), .ZN(new_n761_));
  INV_X1    g560(.A(KEYINPUT115), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n762_), .B1(new_n759_), .B2(KEYINPUT56), .ZN(new_n763_));
  AND2_X1   g562(.A1(new_n569_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n261_), .B(new_n260_), .C1(new_n761_), .C2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(KEYINPUT117), .B1(new_n760_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT56), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n762_), .B(new_n568_), .C1(new_n755_), .C2(new_n756_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n767_), .B1(new_n768_), .B2(KEYINPUT116), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT117), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n757_), .A2(new_n533_), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n569_), .A2(new_n763_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n262_), .B1(new_n771_), .B2(new_n772_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n769_), .A2(new_n770_), .A3(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n234_), .ZN(new_n775_));
  OAI211_X1 g574(.A(new_n233_), .B(new_n775_), .C1(new_n253_), .C2(new_n254_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n249_), .A2(new_n233_), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n257_), .B1(new_n777_), .B2(new_n234_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n776_), .A2(new_n778_), .ZN(new_n779_));
  AND2_X1   g578(.A1(new_n258_), .A2(new_n779_), .ZN(new_n780_));
  NAND2_X1  g579(.A1(new_n570_), .A2(new_n780_), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n766_), .A2(new_n774_), .A3(new_n781_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n782_), .A2(new_n638_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT57), .ZN(new_n784_));
  AOI21_X1  g583(.A(KEYINPUT118), .B1(new_n783_), .B2(new_n784_), .ZN(new_n785_));
  INV_X1    g584(.A(KEYINPUT118), .ZN(new_n786_));
  AOI211_X1 g585(.A(new_n786_), .B(KEYINPUT57), .C1(new_n782_), .C2(new_n638_), .ZN(new_n787_));
  NOR2_X1   g586(.A1(new_n785_), .A2(new_n787_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n606_), .A2(new_n784_), .ZN(new_n789_));
  AND3_X1   g588(.A1(new_n782_), .A2(KEYINPUT119), .A3(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(KEYINPUT119), .B1(new_n782_), .B2(new_n789_), .ZN(new_n791_));
  NAND2_X1  g590(.A1(new_n780_), .A2(new_n569_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n792_), .B1(new_n767_), .B2(new_n761_), .ZN(new_n793_));
  OAI211_X1 g592(.A(new_n793_), .B(KEYINPUT58), .C1(new_n767_), .C2(new_n761_), .ZN(new_n794_));
  INV_X1    g593(.A(KEYINPUT58), .ZN(new_n795_));
  OAI211_X1 g594(.A(new_n569_), .B(new_n780_), .C1(new_n771_), .C2(KEYINPUT56), .ZN(new_n796_));
  NOR2_X1   g595(.A1(new_n761_), .A2(new_n767_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n795_), .B1(new_n796_), .B2(new_n797_), .ZN(new_n798_));
  AND3_X1   g597(.A1(new_n529_), .A2(new_n794_), .A3(new_n798_), .ZN(new_n799_));
  NOR3_X1   g598(.A1(new_n790_), .A2(new_n791_), .A3(new_n799_), .ZN(new_n800_));
  AOI21_X1  g599(.A(new_n639_), .B1(new_n788_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n594_), .A2(new_n262_), .ZN(new_n802_));
  XNOR2_X1  g601(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n803_));
  XOR2_X1   g602(.A(new_n802_), .B(new_n803_), .Z(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT120), .B1(new_n801_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(new_n781_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n769_), .A2(new_n773_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(KEYINPUT117), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n606_), .B1(new_n808_), .B2(new_n774_), .ZN(new_n809_));
  OAI21_X1  g608(.A(new_n786_), .B1(new_n809_), .B2(KEYINPUT57), .ZN(new_n810_));
  NAND2_X1  g609(.A1(new_n782_), .A2(new_n789_), .ZN(new_n811_));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n799_), .B1(new_n811_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n790_), .ZN(new_n814_));
  NAND3_X1  g613(.A1(new_n783_), .A2(KEYINPUT118), .A3(new_n784_), .ZN(new_n815_));
  NAND4_X1  g614(.A1(new_n810_), .A2(new_n813_), .A3(new_n814_), .A4(new_n815_), .ZN(new_n816_));
  NAND2_X1  g615(.A1(new_n816_), .A2(new_n593_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT120), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n802_), .B(new_n803_), .ZN(new_n819_));
  NAND3_X1  g618(.A1(new_n817_), .A2(new_n818_), .A3(new_n819_), .ZN(new_n820_));
  NOR4_X1   g619(.A1(new_n306_), .A2(new_n617_), .A3(new_n453_), .A4(new_n366_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n805_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(G113gat), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n609_), .ZN(new_n825_));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n821_), .A2(new_n826_), .ZN(new_n827_));
  OAI211_X1 g626(.A(new_n813_), .B(new_n814_), .C1(KEYINPUT57), .C2(new_n809_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n828_), .A2(new_n593_), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n827_), .B1(new_n829_), .B2(new_n819_), .ZN(new_n830_));
  AOI211_X1 g629(.A(new_n262_), .B(new_n830_), .C1(new_n822_), .C2(KEYINPUT59), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n825_), .B1(new_n831_), .B2(new_n824_), .ZN(G1340gat));
  AOI211_X1 g631(.A(new_n574_), .B(new_n830_), .C1(new_n822_), .C2(KEYINPUT59), .ZN(new_n833_));
  INV_X1    g632(.A(G120gat), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n834_), .B1(new_n574_), .B2(KEYINPUT60), .ZN(new_n835_));
  OAI21_X1  g634(.A(new_n835_), .B1(KEYINPUT60), .B2(new_n834_), .ZN(new_n836_));
  OAI22_X1  g635(.A1(new_n833_), .A2(new_n834_), .B1(new_n822_), .B2(new_n836_), .ZN(G1341gat));
  INV_X1    g636(.A(G127gat), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n593_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  AOI211_X1 g639(.A(new_n830_), .B(new_n840_), .C1(new_n822_), .C2(KEYINPUT59), .ZN(new_n841_));
  NAND4_X1  g640(.A1(new_n805_), .A2(new_n820_), .A3(new_n639_), .A4(new_n821_), .ZN(new_n842_));
  NAND2_X1  g641(.A1(new_n842_), .A2(new_n838_), .ZN(new_n843_));
  INV_X1    g642(.A(new_n843_), .ZN(new_n844_));
  OAI21_X1  g643(.A(KEYINPUT121), .B1(new_n841_), .B2(new_n844_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n822_), .A2(KEYINPUT59), .ZN(new_n846_));
  INV_X1    g645(.A(new_n830_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n847_), .A3(new_n839_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n843_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n845_), .A2(new_n850_), .ZN(G1342gat));
  INV_X1    g650(.A(G134gat), .ZN(new_n852_));
  NAND3_X1  g651(.A1(new_n823_), .A2(new_n852_), .A3(new_n607_), .ZN(new_n853_));
  AOI211_X1 g652(.A(new_n645_), .B(new_n830_), .C1(new_n822_), .C2(KEYINPUT59), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n854_), .B2(new_n852_), .ZN(G1343gat));
  AND2_X1   g654(.A1(new_n805_), .A2(new_n820_), .ZN(new_n856_));
  NAND4_X1  g655(.A1(new_n306_), .A2(new_n416_), .A3(new_n366_), .A4(new_n449_), .ZN(new_n857_));
  INV_X1    g656(.A(new_n857_), .ZN(new_n858_));
  NAND3_X1  g657(.A1(new_n856_), .A2(new_n609_), .A3(new_n858_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(KEYINPUT122), .B(G141gat), .ZN(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1344gat));
  NAND3_X1  g660(.A1(new_n856_), .A2(new_n575_), .A3(new_n858_), .ZN(new_n862_));
  XOR2_X1   g661(.A(KEYINPUT123), .B(G148gat), .Z(new_n863_));
  XNOR2_X1  g662(.A(new_n862_), .B(new_n863_), .ZN(G1345gat));
  NAND3_X1  g663(.A1(new_n856_), .A2(new_n639_), .A3(new_n858_), .ZN(new_n865_));
  XNOR2_X1  g664(.A(KEYINPUT61), .B(G155gat), .ZN(new_n866_));
  XNOR2_X1  g665(.A(new_n865_), .B(new_n866_), .ZN(G1346gat));
  NAND2_X1  g666(.A1(new_n856_), .A2(new_n858_), .ZN(new_n868_));
  OAI21_X1  g667(.A(G162gat), .B1(new_n868_), .B2(new_n645_), .ZN(new_n869_));
  OR2_X1    g668(.A1(new_n689_), .A2(G162gat), .ZN(new_n870_));
  OAI21_X1  g669(.A(new_n869_), .B1(new_n868_), .B2(new_n870_), .ZN(G1347gat));
  NAND2_X1  g670(.A1(new_n829_), .A2(new_n819_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n306_), .A2(new_n416_), .A3(new_n449_), .ZN(new_n873_));
  NAND3_X1  g672(.A1(new_n872_), .A2(new_n365_), .A3(new_n873_), .ZN(new_n874_));
  INV_X1    g673(.A(new_n874_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(KEYINPUT22), .B(G169gat), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n875_), .A2(new_n609_), .A3(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n873_), .A2(new_n609_), .ZN(new_n878_));
  XOR2_X1   g677(.A(new_n878_), .B(KEYINPUT124), .Z(new_n879_));
  NAND3_X1  g678(.A1(new_n879_), .A2(new_n872_), .A3(new_n365_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n881_));
  NAND3_X1  g680(.A1(new_n880_), .A2(new_n881_), .A3(G169gat), .ZN(new_n882_));
  INV_X1    g681(.A(new_n882_), .ZN(new_n883_));
  AOI21_X1  g682(.A(new_n881_), .B1(new_n880_), .B2(G169gat), .ZN(new_n884_));
  OAI21_X1  g683(.A(new_n877_), .B1(new_n883_), .B2(new_n884_), .ZN(G1348gat));
  AOI21_X1  g684(.A(G176gat), .B1(new_n875_), .B2(new_n575_), .ZN(new_n886_));
  AND2_X1   g685(.A1(new_n856_), .A2(new_n365_), .ZN(new_n887_));
  AND3_X1   g686(.A1(new_n873_), .A2(G176gat), .A3(new_n575_), .ZN(new_n888_));
  AOI21_X1  g687(.A(new_n886_), .B1(new_n887_), .B2(new_n888_), .ZN(G1349gat));
  NOR3_X1   g688(.A1(new_n874_), .A2(new_n271_), .A3(new_n593_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n887_), .A2(new_n639_), .A3(new_n873_), .ZN(new_n891_));
  INV_X1    g690(.A(G183gat), .ZN(new_n892_));
  AOI21_X1  g691(.A(new_n890_), .B1(new_n891_), .B2(new_n892_), .ZN(G1350gat));
  OAI21_X1  g692(.A(G190gat), .B1(new_n874_), .B2(new_n645_), .ZN(new_n894_));
  NAND2_X1  g693(.A1(new_n607_), .A2(new_n272_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n874_), .B2(new_n895_), .ZN(G1351gat));
  NOR4_X1   g695(.A1(new_n305_), .A2(new_n449_), .A3(new_n416_), .A4(new_n365_), .ZN(new_n897_));
  NAND3_X1  g696(.A1(new_n856_), .A2(new_n609_), .A3(new_n897_), .ZN(new_n898_));
  XNOR2_X1  g697(.A(new_n898_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g698(.A1(new_n856_), .A2(new_n575_), .A3(new_n897_), .ZN(new_n900_));
  XNOR2_X1  g699(.A(new_n900_), .B(G204gat), .ZN(G1353gat));
  AOI21_X1  g700(.A(new_n593_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n902_));
  XOR2_X1   g701(.A(new_n902_), .B(KEYINPUT125), .Z(new_n903_));
  NAND3_X1  g702(.A1(new_n856_), .A2(new_n897_), .A3(new_n903_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n905_));
  AND2_X1   g704(.A1(new_n905_), .A2(KEYINPUT126), .ZN(new_n906_));
  NOR2_X1   g705(.A1(new_n904_), .A2(new_n906_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n905_), .B(KEYINPUT126), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n907_), .B1(new_n904_), .B2(new_n908_), .ZN(G1354gat));
  NAND4_X1  g708(.A1(new_n805_), .A2(new_n820_), .A3(new_n529_), .A4(new_n897_), .ZN(new_n910_));
  NAND2_X1  g709(.A1(new_n910_), .A2(G218gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n856_), .A2(new_n897_), .ZN(new_n912_));
  OR2_X1    g711(.A1(new_n689_), .A2(G218gat), .ZN(new_n913_));
  OAI21_X1  g712(.A(new_n911_), .B1(new_n912_), .B2(new_n913_), .ZN(new_n914_));
  INV_X1    g713(.A(KEYINPUT127), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n914_), .A2(new_n915_), .ZN(new_n916_));
  OAI211_X1 g715(.A(KEYINPUT127), .B(new_n911_), .C1(new_n912_), .C2(new_n913_), .ZN(new_n917_));
  NAND2_X1  g716(.A1(new_n916_), .A2(new_n917_), .ZN(G1355gat));
endmodule


