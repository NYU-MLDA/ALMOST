//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:29:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n655_, new_n656_, new_n657_, new_n658_, new_n659_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n714_, new_n715_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n729_, new_n730_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n762_, new_n763_, new_n765_, new_n766_, new_n767_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n785_, new_n786_,
    new_n787_, new_n788_, new_n789_, new_n790_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n860_, new_n861_,
    new_n862_, new_n864_, new_n865_, new_n866_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n872_, new_n873_, new_n875_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n882_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n896_, new_n897_, new_n898_,
    new_n900_, new_n901_, new_n902_, new_n903_, new_n904_, new_n906_,
    new_n907_, new_n908_, new_n909_, new_n910_, new_n911_, new_n912_,
    new_n913_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n922_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n930_, new_n931_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XOR2_X1   g001(.A(G85gat), .B(G92gat), .Z(new_n203_));
  NOR3_X1   g002(.A1(KEYINPUT7), .A2(G99gat), .A3(G106gat), .ZN(new_n204_));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NAND2_X1  g005(.A1(G99gat), .A2(G106gat), .ZN(new_n207_));
  XNOR2_X1  g006(.A(new_n207_), .B(KEYINPUT6), .ZN(new_n208_));
  OAI21_X1  g007(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n208_), .A2(new_n209_), .ZN(new_n210_));
  OAI21_X1  g009(.A(new_n203_), .B1(new_n206_), .B2(new_n210_), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT8), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n211_), .A2(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(KEYINPUT10), .B(G99gat), .Z(new_n214_));
  INV_X1    g013(.A(G106gat), .ZN(new_n215_));
  NAND2_X1  g014(.A1(new_n214_), .A2(new_n215_), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n203_), .A2(KEYINPUT9), .ZN(new_n217_));
  INV_X1    g016(.A(KEYINPUT9), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n218_), .A2(G85gat), .A3(G92gat), .ZN(new_n219_));
  NAND4_X1  g018(.A1(new_n216_), .A2(new_n217_), .A3(new_n208_), .A4(new_n219_), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n213_), .A2(new_n220_), .ZN(new_n221_));
  NOR2_X1   g020(.A1(new_n211_), .A2(new_n212_), .ZN(new_n222_));
  OR3_X1    g021(.A1(new_n221_), .A2(KEYINPUT67), .A3(new_n222_), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n211_), .A2(new_n212_), .ZN(new_n224_));
  NAND3_X1  g023(.A1(new_n224_), .A2(new_n220_), .A3(new_n213_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(KEYINPUT67), .ZN(new_n226_));
  XNOR2_X1  g025(.A(G57gat), .B(G64gat), .ZN(new_n227_));
  XOR2_X1   g026(.A(new_n227_), .B(KEYINPUT11), .Z(new_n228_));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(G71gat), .ZN(new_n229_));
  XNOR2_X1  g028(.A(new_n229_), .B(G78gat), .ZN(new_n230_));
  OR2_X1    g029(.A1(new_n228_), .A2(new_n230_), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n227_), .A2(KEYINPUT11), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n230_), .A2(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n223_), .A2(new_n226_), .A3(KEYINPUT12), .A4(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n225_), .A2(new_n234_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT12), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  AND2_X1   g037(.A1(new_n235_), .A2(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(new_n221_), .A2(new_n222_), .ZN(new_n240_));
  NAND3_X1  g039(.A1(new_n240_), .A2(new_n231_), .A3(new_n233_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G230gat), .A2(G233gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  AND2_X1   g042(.A1(new_n243_), .A2(KEYINPUT68), .ZN(new_n244_));
  NOR2_X1   g043(.A1(new_n243_), .A2(KEYINPUT68), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n239_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n241_), .A2(KEYINPUT66), .A3(new_n236_), .ZN(new_n247_));
  INV_X1    g046(.A(new_n242_), .ZN(new_n248_));
  OAI211_X1 g047(.A(new_n247_), .B(new_n248_), .C1(KEYINPUT66), .C2(new_n241_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n246_), .A2(new_n249_), .ZN(new_n250_));
  XNOR2_X1  g049(.A(G120gat), .B(G148gat), .ZN(new_n251_));
  XNOR2_X1  g050(.A(new_n251_), .B(KEYINPUT5), .ZN(new_n252_));
  XNOR2_X1  g051(.A(G176gat), .B(G204gat), .ZN(new_n253_));
  XOR2_X1   g052(.A(new_n252_), .B(new_n253_), .Z(new_n254_));
  NAND2_X1  g053(.A1(new_n250_), .A2(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(new_n254_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n246_), .A2(new_n249_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(KEYINPUT13), .ZN(new_n259_));
  NAND2_X1  g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  NAND3_X1  g059(.A1(new_n255_), .A2(KEYINPUT13), .A3(new_n257_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  XNOR2_X1  g062(.A(G1gat), .B(G8gat), .ZN(new_n264_));
  XNOR2_X1  g063(.A(new_n264_), .B(KEYINPUT72), .ZN(new_n265_));
  INV_X1    g064(.A(G15gat), .ZN(new_n266_));
  INV_X1    g065(.A(G22gat), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(G15gat), .A2(G22gat), .ZN(new_n269_));
  NAND2_X1  g068(.A1(G1gat), .A2(G8gat), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n268_), .A2(new_n269_), .B1(KEYINPUT14), .B2(new_n270_), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n265_), .B(new_n271_), .ZN(new_n272_));
  XOR2_X1   g071(.A(G29gat), .B(G36gat), .Z(new_n273_));
  XOR2_X1   g072(.A(G43gat), .B(G50gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(new_n273_), .B(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n272_), .A2(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT15), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n275_), .B(new_n277_), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n276_), .B1(new_n278_), .B2(new_n272_), .ZN(new_n279_));
  INV_X1    g078(.A(KEYINPUT76), .ZN(new_n280_));
  NAND2_X1  g079(.A1(G229gat), .A2(G233gat), .ZN(new_n281_));
  INV_X1    g080(.A(new_n281_), .ZN(new_n282_));
  OR3_X1    g081(.A1(new_n279_), .A2(new_n280_), .A3(new_n282_), .ZN(new_n283_));
  AOI21_X1  g082(.A(KEYINPUT75), .B1(new_n272_), .B2(new_n275_), .ZN(new_n284_));
  OAI21_X1  g083(.A(new_n284_), .B1(new_n275_), .B2(new_n272_), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n265_), .B(new_n271_), .Z(new_n286_));
  INV_X1    g085(.A(new_n275_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n286_), .A2(KEYINPUT75), .A3(new_n287_), .ZN(new_n288_));
  NAND3_X1  g087(.A1(new_n285_), .A2(new_n282_), .A3(new_n288_), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n280_), .B1(new_n279_), .B2(new_n282_), .ZN(new_n290_));
  NAND3_X1  g089(.A1(new_n283_), .A2(new_n289_), .A3(new_n290_), .ZN(new_n291_));
  XOR2_X1   g090(.A(G113gat), .B(G141gat), .Z(new_n292_));
  XNOR2_X1  g091(.A(new_n292_), .B(KEYINPUT77), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G169gat), .B(G197gat), .ZN(new_n294_));
  XOR2_X1   g093(.A(new_n293_), .B(new_n294_), .Z(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n291_), .A2(new_n296_), .ZN(new_n297_));
  NAND4_X1  g096(.A1(new_n283_), .A2(new_n289_), .A3(new_n290_), .A4(new_n295_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n297_), .A2(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G231gat), .A2(G233gat), .ZN(new_n300_));
  XNOR2_X1  g099(.A(new_n234_), .B(new_n300_), .ZN(new_n301_));
  XNOR2_X1  g100(.A(new_n301_), .B(new_n286_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n302_), .ZN(new_n303_));
  XOR2_X1   g102(.A(G127gat), .B(G155gat), .Z(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(KEYINPUT16), .ZN(new_n305_));
  XNOR2_X1  g104(.A(G183gat), .B(G211gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n305_), .B(new_n306_), .ZN(new_n307_));
  XOR2_X1   g106(.A(KEYINPUT73), .B(KEYINPUT17), .Z(new_n308_));
  OR3_X1    g107(.A1(new_n303_), .A2(new_n307_), .A3(new_n308_), .ZN(new_n309_));
  OR2_X1    g108(.A1(new_n309_), .A2(KEYINPUT74), .ZN(new_n310_));
  XNOR2_X1  g109(.A(new_n307_), .B(KEYINPUT17), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n303_), .A2(new_n311_), .ZN(new_n312_));
  NAND2_X1  g111(.A1(new_n309_), .A2(KEYINPUT74), .ZN(new_n313_));
  AND3_X1   g112(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n263_), .A2(new_n299_), .A3(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(new_n315_), .B(KEYINPUT99), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G127gat), .B(G134gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(G113gat), .B(G120gat), .ZN(new_n318_));
  XOR2_X1   g117(.A(new_n317_), .B(new_n318_), .Z(new_n319_));
  XNOR2_X1  g118(.A(new_n319_), .B(KEYINPUT31), .ZN(new_n320_));
  XNOR2_X1  g119(.A(KEYINPUT26), .B(G190gat), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT25), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G183gat), .ZN(new_n323_));
  INV_X1    g122(.A(KEYINPUT78), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n323_), .A2(new_n324_), .ZN(new_n325_));
  XNOR2_X1  g124(.A(KEYINPUT25), .B(G183gat), .ZN(new_n326_));
  OAI211_X1 g125(.A(new_n321_), .B(new_n325_), .C1(new_n326_), .C2(new_n324_), .ZN(new_n327_));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n328_));
  NAND3_X1  g127(.A1(new_n328_), .A2(G183gat), .A3(G190gat), .ZN(new_n329_));
  NAND2_X1  g128(.A1(G183gat), .A2(G190gat), .ZN(new_n330_));
  AND3_X1   g129(.A1(new_n330_), .A2(KEYINPUT79), .A3(KEYINPUT23), .ZN(new_n331_));
  AOI21_X1  g130(.A(KEYINPUT79), .B1(new_n330_), .B2(KEYINPUT23), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n329_), .B1(new_n331_), .B2(new_n332_), .ZN(new_n333_));
  NOR3_X1   g132(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n334_));
  NAND2_X1  g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n335_), .A2(KEYINPUT24), .ZN(new_n336_));
  OR2_X1    g135(.A1(G169gat), .A2(G176gat), .ZN(new_n337_));
  AOI21_X1  g136(.A(new_n334_), .B1(new_n336_), .B2(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n327_), .A2(new_n333_), .A3(new_n338_), .ZN(new_n339_));
  NOR2_X1   g138(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n340_));
  XNOR2_X1  g139(.A(new_n340_), .B(G169gat), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n330_), .A2(KEYINPUT23), .ZN(new_n342_));
  AND2_X1   g141(.A1(new_n342_), .A2(new_n329_), .ZN(new_n343_));
  NOR2_X1   g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(new_n341_), .B1(new_n343_), .B2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n339_), .A2(new_n345_), .ZN(new_n346_));
  XNOR2_X1  g145(.A(new_n346_), .B(KEYINPUT30), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT80), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  XNOR2_X1  g148(.A(G71gat), .B(G99gat), .ZN(new_n350_));
  XNOR2_X1  g149(.A(new_n350_), .B(G43gat), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G227gat), .A2(G233gat), .ZN(new_n352_));
  XNOR2_X1  g151(.A(new_n352_), .B(new_n266_), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n351_), .B(new_n353_), .ZN(new_n354_));
  OR2_X1    g153(.A1(new_n349_), .A2(new_n354_), .ZN(new_n355_));
  INV_X1    g154(.A(KEYINPUT30), .ZN(new_n356_));
  XNOR2_X1  g155(.A(new_n346_), .B(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(KEYINPUT80), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n349_), .A2(new_n358_), .A3(new_n354_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n355_), .A2(new_n359_), .ZN(new_n360_));
  AOI21_X1  g159(.A(new_n320_), .B1(new_n360_), .B2(KEYINPUT81), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n361_), .B1(KEYINPUT81), .B2(new_n360_), .ZN(new_n362_));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n363_));
  NAND4_X1  g162(.A1(new_n355_), .A2(new_n363_), .A3(new_n359_), .A4(new_n320_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  XNOR2_X1  g164(.A(G141gat), .B(G148gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(G155gat), .A2(G162gat), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n367_), .A2(KEYINPUT1), .ZN(new_n368_));
  NOR2_X1   g167(.A1(G155gat), .A2(G162gat), .ZN(new_n369_));
  OAI21_X1  g168(.A(new_n367_), .B1(new_n369_), .B2(KEYINPUT1), .ZN(new_n370_));
  AOI21_X1  g169(.A(new_n368_), .B1(new_n370_), .B2(KEYINPUT82), .ZN(new_n371_));
  INV_X1    g170(.A(KEYINPUT1), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n372_), .B1(G155gat), .B2(G162gat), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(new_n374_), .A3(new_n367_), .ZN(new_n375_));
  AOI21_X1  g174(.A(new_n366_), .B1(new_n371_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(new_n367_), .ZN(new_n377_));
  NOR2_X1   g176(.A1(new_n377_), .A2(new_n369_), .ZN(new_n378_));
  INV_X1    g177(.A(new_n378_), .ZN(new_n379_));
  NAND2_X1  g178(.A1(G141gat), .A2(G148gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT2), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n380_), .A2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n382_), .A2(KEYINPUT83), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT83), .ZN(new_n384_));
  NAND3_X1  g183(.A1(new_n380_), .A2(new_n384_), .A3(new_n381_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387_));
  INV_X1    g186(.A(G141gat), .ZN(new_n388_));
  INV_X1    g187(.A(G148gat), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n387_), .A2(new_n388_), .A3(new_n389_), .ZN(new_n390_));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n391_));
  NAND3_X1  g190(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n379_), .B1(new_n386_), .B2(new_n393_), .ZN(new_n394_));
  OAI21_X1  g193(.A(new_n319_), .B1(new_n376_), .B2(new_n394_), .ZN(new_n395_));
  AND3_X1   g194(.A1(new_n380_), .A2(new_n384_), .A3(new_n381_), .ZN(new_n396_));
  AOI21_X1  g195(.A(new_n384_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n396_), .A2(new_n397_), .ZN(new_n398_));
  NAND3_X1  g197(.A1(new_n390_), .A2(new_n391_), .A3(new_n392_), .ZN(new_n399_));
  OAI21_X1  g198(.A(new_n378_), .B1(new_n398_), .B2(new_n399_), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n317_), .B(new_n318_), .ZN(new_n401_));
  AND3_X1   g200(.A1(new_n373_), .A2(new_n374_), .A3(new_n367_), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n374_), .B1(new_n373_), .B2(new_n367_), .ZN(new_n403_));
  NOR3_X1   g202(.A1(new_n402_), .A2(new_n403_), .A3(new_n368_), .ZN(new_n404_));
  OAI211_X1 g203(.A(new_n400_), .B(new_n401_), .C1(new_n404_), .C2(new_n366_), .ZN(new_n405_));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406_));
  NAND3_X1  g205(.A1(new_n395_), .A2(new_n405_), .A3(new_n406_), .ZN(new_n407_));
  AND3_X1   g206(.A1(new_n395_), .A2(new_n405_), .A3(KEYINPUT4), .ZN(new_n408_));
  INV_X1    g207(.A(new_n406_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n409_), .B1(new_n395_), .B2(KEYINPUT4), .ZN(new_n410_));
  OAI21_X1  g209(.A(new_n407_), .B1(new_n408_), .B2(new_n410_), .ZN(new_n411_));
  XNOR2_X1  g210(.A(G1gat), .B(G29gat), .ZN(new_n412_));
  XNOR2_X1  g211(.A(new_n412_), .B(G85gat), .ZN(new_n413_));
  XNOR2_X1  g212(.A(KEYINPUT0), .B(G57gat), .ZN(new_n414_));
  XOR2_X1   g213(.A(new_n413_), .B(new_n414_), .Z(new_n415_));
  INV_X1    g214(.A(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n411_), .A2(new_n416_), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT96), .ZN(new_n418_));
  OAI211_X1 g217(.A(new_n407_), .B(new_n415_), .C1(new_n408_), .C2(new_n410_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n417_), .A2(new_n418_), .A3(new_n419_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n411_), .A2(KEYINPUT96), .A3(new_n416_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  INV_X1    g221(.A(new_n422_), .ZN(new_n423_));
  XOR2_X1   g222(.A(KEYINPUT84), .B(KEYINPUT28), .Z(new_n424_));
  OAI21_X1  g223(.A(new_n400_), .B1(new_n404_), .B2(new_n366_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n424_), .B1(new_n425_), .B2(KEYINPUT29), .ZN(new_n426_));
  NOR2_X1   g225(.A1(new_n376_), .A2(new_n394_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT29), .ZN(new_n428_));
  INV_X1    g227(.A(new_n424_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n427_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n426_), .A2(new_n430_), .ZN(new_n431_));
  XOR2_X1   g230(.A(G22gat), .B(G50gat), .Z(new_n432_));
  XNOR2_X1  g231(.A(new_n431_), .B(new_n432_), .ZN(new_n433_));
  XNOR2_X1  g232(.A(G78gat), .B(G106gat), .ZN(new_n434_));
  XOR2_X1   g233(.A(new_n434_), .B(KEYINPUT89), .Z(new_n435_));
  INV_X1    g234(.A(new_n435_), .ZN(new_n436_));
  INV_X1    g235(.A(G204gat), .ZN(new_n437_));
  OAI21_X1  g236(.A(KEYINPUT86), .B1(new_n437_), .B2(G197gat), .ZN(new_n438_));
  INV_X1    g237(.A(KEYINPUT86), .ZN(new_n439_));
  INV_X1    g238(.A(G197gat), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n439_), .A2(new_n440_), .A3(G204gat), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n437_), .A2(G197gat), .ZN(new_n442_));
  NAND3_X1  g241(.A1(new_n438_), .A2(new_n441_), .A3(new_n442_), .ZN(new_n443_));
  INV_X1    g242(.A(G218gat), .ZN(new_n444_));
  NAND2_X1  g243(.A1(new_n444_), .A2(G211gat), .ZN(new_n445_));
  INV_X1    g244(.A(G211gat), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n446_), .A2(G218gat), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n445_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n443_), .A2(KEYINPUT21), .A3(new_n448_), .ZN(new_n449_));
  INV_X1    g248(.A(KEYINPUT21), .ZN(new_n450_));
  AOI21_X1  g249(.A(KEYINPUT85), .B1(new_n440_), .B2(G204gat), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n440_), .A2(G204gat), .ZN(new_n452_));
  NOR2_X1   g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND3_X1  g252(.A1(new_n440_), .A2(KEYINPUT85), .A3(G204gat), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n450_), .B1(new_n453_), .B2(new_n454_), .ZN(new_n455_));
  NAND4_X1  g254(.A1(new_n438_), .A2(new_n441_), .A3(new_n450_), .A4(new_n442_), .ZN(new_n456_));
  INV_X1    g255(.A(new_n448_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n456_), .A2(new_n457_), .ZN(new_n458_));
  OAI21_X1  g257(.A(new_n449_), .B1(new_n455_), .B2(new_n458_), .ZN(new_n459_));
  INV_X1    g258(.A(KEYINPUT87), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n459_), .A2(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(KEYINPUT85), .ZN(new_n462_));
  OAI21_X1  g261(.A(new_n462_), .B1(new_n437_), .B2(G197gat), .ZN(new_n463_));
  NAND3_X1  g262(.A1(new_n463_), .A2(new_n454_), .A3(new_n442_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n464_), .A2(KEYINPUT21), .ZN(new_n465_));
  NAND3_X1  g264(.A1(new_n465_), .A2(new_n456_), .A3(new_n457_), .ZN(new_n466_));
  NAND3_X1  g265(.A1(new_n466_), .A2(KEYINPUT87), .A3(new_n449_), .ZN(new_n467_));
  AOI22_X1  g266(.A1(new_n461_), .A2(new_n467_), .B1(new_n425_), .B2(KEYINPUT29), .ZN(new_n468_));
  INV_X1    g267(.A(G228gat), .ZN(new_n469_));
  INV_X1    g268(.A(G233gat), .ZN(new_n470_));
  NOR2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  OAI21_X1  g271(.A(KEYINPUT88), .B1(new_n468_), .B2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT29), .B1(new_n376_), .B2(new_n394_), .ZN(new_n474_));
  AND3_X1   g273(.A1(new_n466_), .A2(KEYINPUT87), .A3(new_n449_), .ZN(new_n475_));
  AOI21_X1  g274(.A(KEYINPUT87), .B1(new_n466_), .B2(new_n449_), .ZN(new_n476_));
  OAI21_X1  g275(.A(new_n474_), .B1(new_n475_), .B2(new_n476_), .ZN(new_n477_));
  INV_X1    g276(.A(KEYINPUT88), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n477_), .A2(new_n478_), .A3(new_n471_), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n473_), .A2(new_n479_), .ZN(new_n480_));
  NAND3_X1  g279(.A1(new_n474_), .A2(new_n472_), .A3(new_n459_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n436_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  INV_X1    g281(.A(new_n481_), .ZN(new_n483_));
  AOI211_X1 g282(.A(new_n435_), .B(new_n483_), .C1(new_n473_), .C2(new_n479_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n433_), .B1(new_n482_), .B2(new_n484_), .ZN(new_n485_));
  NOR3_X1   g284(.A1(new_n468_), .A2(KEYINPUT88), .A3(new_n472_), .ZN(new_n486_));
  AOI21_X1  g285(.A(new_n478_), .B1(new_n477_), .B2(new_n471_), .ZN(new_n487_));
  OAI21_X1  g286(.A(new_n481_), .B1(new_n486_), .B2(new_n487_), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(new_n435_), .ZN(new_n489_));
  INV_X1    g288(.A(new_n433_), .ZN(new_n490_));
  NAND3_X1  g289(.A1(new_n480_), .A2(new_n436_), .A3(new_n481_), .ZN(new_n491_));
  NAND3_X1  g290(.A1(new_n489_), .A2(new_n490_), .A3(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n485_), .A2(new_n492_), .ZN(new_n493_));
  INV_X1    g292(.A(KEYINPUT27), .ZN(new_n494_));
  XNOR2_X1  g293(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n495_));
  XNOR2_X1  g294(.A(new_n495_), .B(KEYINPUT93), .ZN(new_n496_));
  XNOR2_X1  g295(.A(G8gat), .B(G36gat), .ZN(new_n497_));
  AND2_X1   g296(.A1(new_n496_), .A2(new_n497_), .ZN(new_n498_));
  NOR2_X1   g297(.A1(new_n496_), .A2(new_n497_), .ZN(new_n499_));
  NOR2_X1   g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  XNOR2_X1  g299(.A(G64gat), .B(G92gat), .ZN(new_n501_));
  NAND2_X1  g300(.A1(new_n500_), .A2(new_n501_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n496_), .B(new_n497_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n501_), .ZN(new_n504_));
  NAND2_X1  g303(.A1(new_n503_), .A2(new_n504_), .ZN(new_n505_));
  NAND2_X1  g304(.A1(new_n502_), .A2(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT20), .ZN(new_n507_));
  NOR2_X1   g306(.A1(new_n343_), .A2(new_n334_), .ZN(new_n508_));
  INV_X1    g307(.A(G183gat), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(KEYINPUT25), .ZN(new_n510_));
  INV_X1    g309(.A(G190gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n511_), .A2(KEYINPUT26), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT26), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n513_), .A2(G190gat), .ZN(new_n514_));
  NAND4_X1  g313(.A1(new_n323_), .A2(new_n510_), .A3(new_n512_), .A4(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(KEYINPUT90), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n337_), .A2(KEYINPUT24), .A3(new_n335_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n515_), .A2(new_n516_), .A3(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n516_), .B1(new_n515_), .B2(new_n517_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n508_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n333_), .B1(G183gat), .B2(G190gat), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n335_), .A2(KEYINPUT91), .ZN(new_n522_));
  OR2_X1    g321(.A1(new_n335_), .A2(KEYINPUT91), .ZN(new_n523_));
  XNOR2_X1  g322(.A(KEYINPUT22), .B(G169gat), .ZN(new_n524_));
  INV_X1    g323(.A(G176gat), .ZN(new_n525_));
  AOI22_X1  g324(.A1(new_n522_), .A2(new_n523_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n521_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n520_), .A2(new_n527_), .ZN(new_n528_));
  AOI21_X1  g327(.A(new_n507_), .B1(new_n528_), .B2(new_n459_), .ZN(new_n529_));
  NOR2_X1   g328(.A1(new_n346_), .A2(new_n459_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(new_n529_), .A2(new_n531_), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G226gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n533_), .B(KEYINPUT19), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n532_), .A2(new_n534_), .ZN(new_n535_));
  NAND4_X1  g334(.A1(new_n520_), .A2(new_n527_), .A3(new_n466_), .A4(new_n449_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n507_), .B1(new_n346_), .B2(new_n459_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n534_), .ZN(new_n538_));
  NAND3_X1  g337(.A1(new_n536_), .A2(new_n537_), .A3(new_n538_), .ZN(new_n539_));
  AOI21_X1  g338(.A(new_n506_), .B1(new_n535_), .B2(new_n539_), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n538_), .B1(new_n529_), .B2(new_n531_), .ZN(new_n541_));
  AND2_X1   g340(.A1(new_n502_), .A2(new_n505_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n539_), .ZN(new_n543_));
  NOR3_X1   g342(.A1(new_n541_), .A2(new_n542_), .A3(new_n543_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n494_), .B1(new_n540_), .B2(new_n544_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n529_), .A2(new_n538_), .A3(new_n531_), .ZN(new_n546_));
  NAND4_X1  g345(.A1(new_n461_), .A2(new_n467_), .A3(new_n527_), .A4(new_n520_), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n547_), .A2(new_n537_), .ZN(new_n548_));
  OAI21_X1  g347(.A(new_n546_), .B1(new_n548_), .B2(new_n538_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n549_), .A2(new_n542_), .ZN(new_n550_));
  NAND3_X1  g349(.A1(new_n535_), .A2(new_n506_), .A3(new_n539_), .ZN(new_n551_));
  NAND3_X1  g350(.A1(new_n550_), .A2(KEYINPUT27), .A3(new_n551_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n545_), .A2(new_n552_), .ZN(new_n553_));
  NOR4_X1   g352(.A1(new_n365_), .A2(new_n423_), .A3(new_n493_), .A4(new_n553_), .ZN(new_n554_));
  INV_X1    g353(.A(KEYINPUT97), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT32), .ZN(new_n556_));
  AOI21_X1  g355(.A(new_n556_), .B1(new_n502_), .B2(new_n505_), .ZN(new_n557_));
  INV_X1    g356(.A(new_n557_), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n558_), .A2(new_n535_), .A3(new_n539_), .ZN(new_n559_));
  AND3_X1   g358(.A1(new_n420_), .A2(new_n421_), .A3(new_n559_), .ZN(new_n560_));
  AOI22_X1  g359(.A1(new_n520_), .A2(new_n527_), .B1(new_n466_), .B2(new_n449_), .ZN(new_n561_));
  NOR4_X1   g360(.A1(new_n561_), .A2(new_n530_), .A3(new_n507_), .A4(new_n534_), .ZN(new_n562_));
  AOI21_X1  g361(.A(new_n538_), .B1(new_n547_), .B2(new_n537_), .ZN(new_n563_));
  OAI21_X1  g362(.A(new_n557_), .B1(new_n562_), .B2(new_n563_), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n564_), .A2(KEYINPUT95), .ZN(new_n565_));
  INV_X1    g364(.A(KEYINPUT95), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n566_), .B(new_n557_), .C1(new_n562_), .C2(new_n563_), .ZN(new_n567_));
  NAND2_X1  g366(.A1(new_n565_), .A2(new_n567_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n542_), .B1(new_n541_), .B2(new_n543_), .ZN(new_n569_));
  NAND3_X1  g368(.A1(new_n395_), .A2(new_n405_), .A3(new_n409_), .ZN(new_n570_));
  OAI21_X1  g369(.A(new_n406_), .B1(new_n395_), .B2(KEYINPUT4), .ZN(new_n571_));
  OAI211_X1 g370(.A(new_n570_), .B(new_n416_), .C1(new_n408_), .C2(new_n571_), .ZN(new_n572_));
  AND3_X1   g371(.A1(new_n551_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n573_));
  NOR2_X1   g372(.A1(KEYINPUT94), .A2(KEYINPUT33), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n419_), .B(new_n574_), .Z(new_n575_));
  AOI22_X1  g374(.A1(new_n560_), .A2(new_n568_), .B1(new_n573_), .B2(new_n575_), .ZN(new_n576_));
  OAI21_X1  g375(.A(new_n555_), .B1(new_n576_), .B2(new_n493_), .ZN(new_n577_));
  NOR3_X1   g376(.A1(new_n482_), .A2(new_n484_), .A3(new_n433_), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n490_), .B1(new_n489_), .B2(new_n491_), .ZN(new_n579_));
  NOR2_X1   g378(.A1(new_n578_), .A2(new_n579_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n545_), .A2(new_n552_), .A3(new_n422_), .ZN(new_n581_));
  OAI21_X1  g380(.A(KEYINPUT98), .B1(new_n580_), .B2(new_n581_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n566_), .B1(new_n549_), .B2(new_n557_), .ZN(new_n583_));
  INV_X1    g382(.A(new_n567_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n583_), .A2(new_n584_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n420_), .A2(new_n421_), .A3(new_n559_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n551_), .A2(new_n569_), .A3(new_n572_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(new_n419_), .B(new_n574_), .ZN(new_n588_));
  OAI22_X1  g387(.A1(new_n585_), .A2(new_n586_), .B1(new_n587_), .B2(new_n588_), .ZN(new_n589_));
  NAND3_X1  g388(.A1(new_n589_), .A2(new_n580_), .A3(KEYINPUT97), .ZN(new_n590_));
  AND2_X1   g389(.A1(new_n545_), .A2(new_n552_), .ZN(new_n591_));
  INV_X1    g390(.A(KEYINPUT98), .ZN(new_n592_));
  NAND4_X1  g391(.A1(new_n591_), .A2(new_n493_), .A3(new_n592_), .A4(new_n422_), .ZN(new_n593_));
  NAND4_X1  g392(.A1(new_n577_), .A2(new_n582_), .A3(new_n590_), .A4(new_n593_), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n554_), .B1(new_n594_), .B2(new_n365_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G190gat), .B(G218gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597_));
  XNOR2_X1  g396(.A(new_n596_), .B(new_n597_), .ZN(new_n598_));
  XOR2_X1   g397(.A(new_n598_), .B(KEYINPUT36), .Z(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT70), .ZN(new_n600_));
  NAND2_X1  g399(.A1(G232gat), .A2(G233gat), .ZN(new_n601_));
  XOR2_X1   g400(.A(new_n601_), .B(KEYINPUT34), .Z(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT69), .B(KEYINPUT35), .ZN(new_n603_));
  AOI22_X1  g402(.A1(new_n240_), .A2(new_n275_), .B1(new_n602_), .B2(new_n603_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n223_), .A2(new_n226_), .ZN(new_n605_));
  OAI21_X1  g404(.A(new_n604_), .B1(new_n605_), .B2(new_n278_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n602_), .A2(new_n603_), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  NOR2_X1   g408(.A1(new_n606_), .A2(new_n607_), .ZN(new_n610_));
  OAI21_X1  g409(.A(new_n600_), .B1(new_n609_), .B2(new_n610_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n606_), .A2(new_n607_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n598_), .A2(KEYINPUT36), .ZN(new_n613_));
  NAND3_X1  g412(.A1(new_n612_), .A2(new_n613_), .A3(new_n608_), .ZN(new_n614_));
  AND2_X1   g413(.A1(new_n611_), .A2(new_n614_), .ZN(new_n615_));
  NOR2_X1   g414(.A1(new_n595_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n316_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT100), .ZN(new_n618_));
  XNOR2_X1  g417(.A(new_n617_), .B(new_n618_), .ZN(new_n619_));
  AOI21_X1  g418(.A(new_n202_), .B1(new_n619_), .B2(new_n423_), .ZN(new_n620_));
  INV_X1    g419(.A(new_n299_), .ZN(new_n621_));
  NOR2_X1   g420(.A1(new_n595_), .A2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT37), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n615_), .A2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(new_n614_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n600_), .B(KEYINPUT71), .ZN(new_n626_));
  AOI21_X1  g425(.A(new_n626_), .B1(new_n612_), .B2(new_n608_), .ZN(new_n627_));
  OAI21_X1  g426(.A(KEYINPUT37), .B1(new_n625_), .B2(new_n627_), .ZN(new_n628_));
  AND2_X1   g427(.A1(new_n624_), .A2(new_n628_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n310_), .A2(new_n312_), .A3(new_n313_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n629_), .A2(new_n630_), .ZN(new_n631_));
  AND3_X1   g430(.A1(new_n622_), .A2(new_n263_), .A3(new_n631_), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n632_), .A2(new_n202_), .A3(new_n423_), .ZN(new_n633_));
  XOR2_X1   g432(.A(new_n633_), .B(KEYINPUT38), .Z(new_n634_));
  OR2_X1    g433(.A1(new_n620_), .A2(new_n634_), .ZN(G1324gat));
  XNOR2_X1  g434(.A(KEYINPUT102), .B(KEYINPUT40), .ZN(new_n636_));
  OAI21_X1  g435(.A(G8gat), .B1(new_n617_), .B2(new_n591_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(new_n637_), .B(KEYINPUT39), .ZN(new_n638_));
  INV_X1    g437(.A(G8gat), .ZN(new_n639_));
  NAND3_X1  g438(.A1(new_n632_), .A2(new_n639_), .A3(new_n553_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT101), .ZN(new_n641_));
  AOI21_X1  g440(.A(new_n636_), .B1(new_n638_), .B2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT39), .ZN(new_n643_));
  OR2_X1    g442(.A1(new_n637_), .A2(new_n643_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n637_), .A2(new_n643_), .ZN(new_n645_));
  AND4_X1   g444(.A1(new_n641_), .A2(new_n644_), .A3(new_n645_), .A4(new_n636_), .ZN(new_n646_));
  NOR2_X1   g445(.A1(new_n642_), .A2(new_n646_), .ZN(G1325gat));
  INV_X1    g446(.A(new_n365_), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n266_), .B1(new_n619_), .B2(new_n648_), .ZN(new_n649_));
  XOR2_X1   g448(.A(KEYINPUT103), .B(KEYINPUT41), .Z(new_n650_));
  OR2_X1    g449(.A1(new_n649_), .A2(new_n650_), .ZN(new_n651_));
  NAND2_X1  g450(.A1(new_n649_), .A2(new_n650_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n632_), .A2(new_n266_), .A3(new_n648_), .ZN(new_n653_));
  NAND3_X1  g452(.A1(new_n651_), .A2(new_n652_), .A3(new_n653_), .ZN(G1326gat));
  NAND3_X1  g453(.A1(new_n632_), .A2(new_n267_), .A3(new_n493_), .ZN(new_n655_));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n619_), .A2(new_n493_), .ZN(new_n657_));
  AOI21_X1  g456(.A(new_n656_), .B1(new_n657_), .B2(G22gat), .ZN(new_n658_));
  AOI211_X1 g457(.A(KEYINPUT42), .B(new_n267_), .C1(new_n619_), .C2(new_n493_), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n655_), .B1(new_n658_), .B2(new_n659_), .ZN(G1327gat));
  INV_X1    g459(.A(new_n615_), .ZN(new_n661_));
  NOR3_X1   g460(.A1(new_n314_), .A2(new_n262_), .A3(new_n661_), .ZN(new_n662_));
  AND2_X1   g461(.A1(new_n622_), .A2(new_n662_), .ZN(new_n663_));
  INV_X1    g462(.A(G29gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(new_n664_), .A3(new_n423_), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n263_), .A2(new_n299_), .A3(new_n630_), .ZN(new_n666_));
  INV_X1    g465(.A(new_n666_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n668_));
  NAND2_X1  g467(.A1(new_n594_), .A2(new_n365_), .ZN(new_n669_));
  INV_X1    g468(.A(new_n554_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n669_), .A2(new_n670_), .ZN(new_n671_));
  AOI21_X1  g470(.A(new_n668_), .B1(new_n671_), .B2(new_n629_), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n624_), .A2(new_n628_), .ZN(new_n673_));
  NOR3_X1   g472(.A1(new_n595_), .A2(KEYINPUT43), .A3(new_n673_), .ZN(new_n674_));
  OAI211_X1 g473(.A(KEYINPUT44), .B(new_n667_), .C1(new_n672_), .C2(new_n674_), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n675_), .A2(new_n676_), .ZN(new_n677_));
  NAND3_X1  g476(.A1(new_n671_), .A2(new_n668_), .A3(new_n629_), .ZN(new_n678_));
  OAI21_X1  g477(.A(KEYINPUT43), .B1(new_n595_), .B2(new_n673_), .ZN(new_n679_));
  AOI21_X1  g478(.A(new_n666_), .B1(new_n678_), .B2(new_n679_), .ZN(new_n680_));
  NAND3_X1  g479(.A1(new_n680_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n681_));
  OAI21_X1  g480(.A(new_n667_), .B1(new_n672_), .B2(new_n674_), .ZN(new_n682_));
  XOR2_X1   g481(.A(KEYINPUT104), .B(KEYINPUT44), .Z(new_n683_));
  AOI22_X1  g482(.A1(new_n677_), .A2(new_n681_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(new_n423_), .ZN(new_n685_));
  AND3_X1   g484(.A1(new_n685_), .A2(KEYINPUT106), .A3(G29gat), .ZN(new_n686_));
  AOI21_X1  g485(.A(KEYINPUT106), .B1(new_n685_), .B2(G29gat), .ZN(new_n687_));
  OAI21_X1  g486(.A(new_n665_), .B1(new_n686_), .B2(new_n687_), .ZN(G1328gat));
  INV_X1    g487(.A(G36gat), .ZN(new_n689_));
  NAND3_X1  g488(.A1(new_n663_), .A2(new_n689_), .A3(new_n553_), .ZN(new_n690_));
  XNOR2_X1  g489(.A(new_n690_), .B(KEYINPUT45), .ZN(new_n691_));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n692_));
  NAND2_X1  g491(.A1(new_n677_), .A2(new_n681_), .ZN(new_n693_));
  AOI21_X1  g492(.A(new_n591_), .B1(new_n682_), .B2(new_n683_), .ZN(new_n694_));
  AOI211_X1 g493(.A(new_n692_), .B(new_n689_), .C1(new_n693_), .C2(new_n694_), .ZN(new_n695_));
  NOR2_X1   g494(.A1(new_n675_), .A2(new_n676_), .ZN(new_n696_));
  AOI21_X1  g495(.A(KEYINPUT105), .B1(new_n680_), .B2(KEYINPUT44), .ZN(new_n697_));
  OAI21_X1  g496(.A(new_n694_), .B1(new_n696_), .B2(new_n697_), .ZN(new_n698_));
  AOI21_X1  g497(.A(KEYINPUT107), .B1(new_n698_), .B2(G36gat), .ZN(new_n699_));
  OAI21_X1  g498(.A(new_n691_), .B1(new_n695_), .B2(new_n699_), .ZN(new_n700_));
  INV_X1    g499(.A(KEYINPUT46), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n700_), .A2(new_n701_), .ZN(new_n702_));
  OAI211_X1 g501(.A(KEYINPUT46), .B(new_n691_), .C1(new_n695_), .C2(new_n699_), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n702_), .A2(new_n703_), .ZN(G1329gat));
  NAND3_X1  g503(.A1(new_n684_), .A2(G43gat), .A3(new_n648_), .ZN(new_n705_));
  AOI21_X1  g504(.A(G43gat), .B1(new_n663_), .B2(new_n648_), .ZN(new_n706_));
  INV_X1    g505(.A(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n705_), .A2(new_n707_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n708_), .A2(new_n710_), .ZN(new_n711_));
  NAND3_X1  g510(.A1(new_n705_), .A2(new_n707_), .A3(new_n709_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n711_), .A2(new_n712_), .ZN(G1330gat));
  AOI21_X1  g512(.A(G50gat), .B1(new_n663_), .B2(new_n493_), .ZN(new_n714_));
  AND2_X1   g513(.A1(new_n493_), .A2(G50gat), .ZN(new_n715_));
  AOI21_X1  g514(.A(new_n714_), .B1(new_n684_), .B2(new_n715_), .ZN(G1331gat));
  AND4_X1   g515(.A1(new_n616_), .A2(new_n621_), .A3(new_n262_), .A4(new_n314_), .ZN(new_n717_));
  NAND3_X1  g516(.A1(new_n717_), .A2(G57gat), .A3(new_n423_), .ZN(new_n718_));
  AOI21_X1  g517(.A(KEYINPUT109), .B1(new_n671_), .B2(new_n621_), .ZN(new_n719_));
  INV_X1    g518(.A(KEYINPUT109), .ZN(new_n720_));
  NOR3_X1   g519(.A1(new_n595_), .A2(new_n720_), .A3(new_n299_), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n719_), .A2(new_n721_), .ZN(new_n722_));
  NOR3_X1   g521(.A1(new_n263_), .A2(new_n629_), .A3(new_n630_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(new_n423_), .A3(new_n723_), .ZN(new_n724_));
  INV_X1    g523(.A(G57gat), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n724_), .A2(new_n725_), .ZN(new_n726_));
  AND2_X1   g525(.A1(new_n726_), .A2(KEYINPUT110), .ZN(new_n727_));
  NOR2_X1   g526(.A1(new_n726_), .A2(KEYINPUT110), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n718_), .B1(new_n727_), .B2(new_n728_), .ZN(new_n729_));
  INV_X1    g528(.A(KEYINPUT111), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n729_), .B(new_n730_), .ZN(G1332gat));
  INV_X1    g530(.A(G64gat), .ZN(new_n732_));
  AOI21_X1  g531(.A(new_n732_), .B1(new_n717_), .B2(new_n553_), .ZN(new_n733_));
  XOR2_X1   g532(.A(new_n733_), .B(KEYINPUT48), .Z(new_n734_));
  NAND2_X1  g533(.A1(new_n722_), .A2(new_n723_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n735_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n736_), .A2(new_n732_), .A3(new_n553_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n734_), .A2(new_n737_), .ZN(G1333gat));
  INV_X1    g537(.A(G71gat), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n739_), .B1(new_n717_), .B2(new_n648_), .ZN(new_n740_));
  XOR2_X1   g539(.A(new_n740_), .B(KEYINPUT49), .Z(new_n741_));
  NAND3_X1  g540(.A1(new_n736_), .A2(new_n739_), .A3(new_n648_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1334gat));
  INV_X1    g542(.A(G78gat), .ZN(new_n744_));
  AOI21_X1  g543(.A(new_n744_), .B1(new_n717_), .B2(new_n493_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n746_));
  XNOR2_X1  g545(.A(new_n745_), .B(new_n746_), .ZN(new_n747_));
  NAND3_X1  g546(.A1(new_n736_), .A2(new_n744_), .A3(new_n493_), .ZN(new_n748_));
  NAND2_X1  g547(.A1(new_n747_), .A2(new_n748_), .ZN(G1335gat));
  NAND2_X1  g548(.A1(new_n678_), .A2(new_n679_), .ZN(new_n750_));
  NOR3_X1   g549(.A1(new_n263_), .A2(new_n314_), .A3(new_n299_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n750_), .A2(new_n751_), .ZN(new_n752_));
  OAI21_X1  g551(.A(G85gat), .B1(new_n752_), .B2(new_n422_), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n263_), .A2(new_n314_), .A3(new_n661_), .ZN(new_n754_));
  NAND3_X1  g553(.A1(new_n722_), .A2(KEYINPUT113), .A3(new_n754_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n754_), .B1(new_n719_), .B2(new_n721_), .ZN(new_n756_));
  INV_X1    g555(.A(KEYINPUT113), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AND2_X1   g557(.A1(new_n755_), .A2(new_n758_), .ZN(new_n759_));
  OR2_X1    g558(.A1(new_n422_), .A2(G85gat), .ZN(new_n760_));
  OAI21_X1  g559(.A(new_n753_), .B1(new_n759_), .B2(new_n760_), .ZN(G1336gat));
  OAI21_X1  g560(.A(G92gat), .B1(new_n752_), .B2(new_n591_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n591_), .A2(G92gat), .ZN(new_n763_));
  OAI21_X1  g562(.A(new_n762_), .B1(new_n759_), .B2(new_n763_), .ZN(G1337gat));
  OAI21_X1  g563(.A(G99gat), .B1(new_n752_), .B2(new_n365_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n648_), .A2(new_n214_), .ZN(new_n766_));
  OAI21_X1  g565(.A(new_n765_), .B1(new_n759_), .B2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g567(.A(KEYINPUT114), .ZN(new_n769_));
  NOR2_X1   g568(.A1(new_n580_), .A2(G106gat), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  OAI21_X1  g570(.A(new_n769_), .B1(new_n759_), .B2(new_n771_), .ZN(new_n772_));
  NAND2_X1  g571(.A1(new_n755_), .A2(new_n758_), .ZN(new_n773_));
  NAND3_X1  g572(.A1(new_n773_), .A2(KEYINPUT114), .A3(new_n770_), .ZN(new_n774_));
  NAND2_X1  g573(.A1(new_n772_), .A2(new_n774_), .ZN(new_n775_));
  NAND3_X1  g574(.A1(new_n750_), .A2(new_n493_), .A3(new_n751_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n776_), .A2(G106gat), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n777_), .A2(new_n778_), .A3(new_n779_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n779_), .B1(new_n777_), .B2(new_n778_), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n781_), .B1(new_n778_), .B2(new_n777_), .ZN(new_n782_));
  XNOR2_X1  g581(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n775_), .A2(new_n780_), .A3(new_n782_), .A4(new_n783_), .ZN(new_n784_));
  INV_X1    g583(.A(new_n783_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n782_), .A2(new_n780_), .ZN(new_n786_));
  AOI21_X1  g585(.A(KEYINPUT114), .B1(new_n773_), .B2(new_n770_), .ZN(new_n787_));
  AOI211_X1 g586(.A(new_n769_), .B(new_n771_), .C1(new_n755_), .C2(new_n758_), .ZN(new_n788_));
  NOR2_X1   g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  OAI21_X1  g588(.A(new_n785_), .B1(new_n786_), .B2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n784_), .A2(new_n790_), .ZN(G1339gat));
  NAND4_X1  g590(.A1(new_n263_), .A2(new_n314_), .A3(new_n621_), .A4(new_n673_), .ZN(new_n792_));
  XOR2_X1   g591(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n792_), .A2(new_n794_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n631_), .A2(new_n263_), .A3(new_n621_), .A4(new_n793_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n795_), .A2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n257_), .A2(new_n299_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n799_));
  NAND2_X1  g598(.A1(new_n246_), .A2(new_n799_), .ZN(new_n800_));
  OAI211_X1 g599(.A(new_n239_), .B(KEYINPUT55), .C1(new_n244_), .C2(new_n245_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n239_), .A2(new_n241_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(new_n248_), .ZN(new_n803_));
  NAND3_X1  g602(.A1(new_n800_), .A2(new_n801_), .A3(new_n803_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n804_), .A2(new_n254_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT56), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n805_), .A2(new_n806_), .ZN(new_n807_));
  NAND3_X1  g606(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n254_), .ZN(new_n808_));
  AOI21_X1  g607(.A(new_n798_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n258_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n285_), .A2(new_n281_), .A3(new_n288_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n811_), .A2(KEYINPUT118), .A3(new_n296_), .ZN(new_n812_));
  OAI21_X1  g611(.A(new_n812_), .B1(new_n281_), .B2(new_n279_), .ZN(new_n813_));
  AOI21_X1  g612(.A(KEYINPUT118), .B1(new_n811_), .B2(new_n296_), .ZN(new_n814_));
  OAI21_X1  g613(.A(new_n298_), .B1(new_n813_), .B2(new_n814_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(new_n815_), .B(KEYINPUT119), .ZN(new_n816_));
  NOR2_X1   g615(.A1(new_n810_), .A2(new_n816_), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n661_), .B1(new_n809_), .B2(new_n817_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(KEYINPUT120), .A2(KEYINPUT57), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n818_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n257_), .ZN(new_n821_));
  INV_X1    g620(.A(KEYINPUT119), .ZN(new_n822_));
  OR2_X1    g621(.A1(new_n815_), .A2(new_n822_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n815_), .A2(new_n822_), .ZN(new_n824_));
  AOI21_X1  g623(.A(new_n821_), .B1(new_n823_), .B2(new_n824_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n804_), .A2(KEYINPUT56), .A3(new_n254_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT56), .B1(new_n804_), .B2(new_n254_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n825_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT58), .ZN(new_n829_));
  AOI21_X1  g628(.A(new_n673_), .B1(new_n828_), .B2(new_n829_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n825_), .B(KEYINPUT58), .C1(new_n826_), .C2(new_n827_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n819_), .ZN(new_n833_));
  OAI211_X1 g632(.A(new_n661_), .B(new_n833_), .C1(new_n809_), .C2(new_n817_), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n820_), .A2(new_n832_), .A3(new_n834_), .ZN(new_n835_));
  AOI21_X1  g634(.A(new_n797_), .B1(new_n835_), .B2(new_n630_), .ZN(new_n836_));
  NOR4_X1   g635(.A1(new_n365_), .A2(new_n422_), .A3(new_n493_), .A4(new_n553_), .ZN(new_n837_));
  XOR2_X1   g636(.A(new_n837_), .B(KEYINPUT121), .Z(new_n838_));
  INV_X1    g637(.A(new_n838_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n836_), .A2(new_n839_), .ZN(new_n840_));
  INV_X1    g639(.A(G113gat), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n840_), .A2(new_n841_), .A3(new_n299_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT59), .ZN(new_n843_));
  OAI21_X1  g642(.A(new_n843_), .B1(new_n836_), .B2(new_n839_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n817_), .ZN(new_n845_));
  OAI211_X1 g644(.A(new_n299_), .B(new_n257_), .C1(new_n826_), .C2(new_n827_), .ZN(new_n846_));
  AOI21_X1  g645(.A(new_n615_), .B1(new_n845_), .B2(new_n846_), .ZN(new_n847_));
  AOI22_X1  g646(.A1(new_n847_), .A2(new_n833_), .B1(new_n830_), .B2(new_n831_), .ZN(new_n848_));
  AOI21_X1  g647(.A(new_n314_), .B1(new_n848_), .B2(new_n820_), .ZN(new_n849_));
  OAI211_X1 g648(.A(KEYINPUT59), .B(new_n838_), .C1(new_n849_), .C2(new_n797_), .ZN(new_n850_));
  AND3_X1   g649(.A1(new_n844_), .A2(new_n850_), .A3(KEYINPUT122), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT122), .B1(new_n844_), .B2(new_n850_), .ZN(new_n852_));
  NOR3_X1   g651(.A1(new_n851_), .A2(new_n852_), .A3(new_n621_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n842_), .B1(new_n853_), .B2(new_n841_), .ZN(G1340gat));
  INV_X1    g653(.A(G120gat), .ZN(new_n855_));
  OAI21_X1  g654(.A(new_n855_), .B1(new_n263_), .B2(KEYINPUT60), .ZN(new_n856_));
  OAI211_X1 g655(.A(new_n840_), .B(new_n856_), .C1(KEYINPUT60), .C2(new_n855_), .ZN(new_n857_));
  AOI21_X1  g656(.A(new_n263_), .B1(new_n844_), .B2(new_n850_), .ZN(new_n858_));
  OAI21_X1  g657(.A(new_n857_), .B1(new_n858_), .B2(new_n855_), .ZN(G1341gat));
  INV_X1    g658(.A(G127gat), .ZN(new_n860_));
  NAND3_X1  g659(.A1(new_n840_), .A2(new_n860_), .A3(new_n314_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n851_), .A2(new_n852_), .A3(new_n630_), .ZN(new_n862_));
  OAI21_X1  g661(.A(new_n861_), .B1(new_n862_), .B2(new_n860_), .ZN(G1342gat));
  INV_X1    g662(.A(G134gat), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n840_), .A2(new_n864_), .A3(new_n615_), .ZN(new_n865_));
  NOR3_X1   g664(.A1(new_n851_), .A2(new_n852_), .A3(new_n673_), .ZN(new_n866_));
  OAI21_X1  g665(.A(new_n865_), .B1(new_n866_), .B2(new_n864_), .ZN(G1343gat));
  NAND2_X1  g666(.A1(new_n835_), .A2(new_n630_), .ZN(new_n868_));
  INV_X1    g667(.A(new_n797_), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n868_), .A2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n648_), .A2(new_n580_), .ZN(new_n871_));
  AND4_X1   g670(.A1(new_n423_), .A2(new_n870_), .A3(new_n591_), .A4(new_n871_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n872_), .A2(new_n299_), .ZN(new_n873_));
  XNOR2_X1  g672(.A(new_n873_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g673(.A1(new_n872_), .A2(new_n262_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g675(.A1(new_n872_), .A2(new_n314_), .ZN(new_n877_));
  XNOR2_X1  g676(.A(KEYINPUT61), .B(G155gat), .ZN(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  AOI21_X1  g678(.A(G162gat), .B1(new_n872_), .B2(new_n615_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n629_), .A2(G162gat), .ZN(new_n881_));
  XOR2_X1   g680(.A(new_n881_), .B(KEYINPUT123), .Z(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n872_), .B2(new_n882_), .ZN(G1347gat));
  NOR4_X1   g682(.A1(new_n365_), .A2(new_n591_), .A3(new_n493_), .A4(new_n423_), .ZN(new_n884_));
  INV_X1    g683(.A(new_n884_), .ZN(new_n885_));
  OAI21_X1  g684(.A(KEYINPUT124), .B1(new_n836_), .B2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887_));
  OAI211_X1 g686(.A(new_n887_), .B(new_n884_), .C1(new_n849_), .C2(new_n797_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n886_), .A2(new_n888_), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n889_), .A2(new_n524_), .A3(new_n299_), .ZN(new_n890_));
  NAND3_X1  g689(.A1(new_n870_), .A2(new_n299_), .A3(new_n884_), .ZN(new_n891_));
  INV_X1    g690(.A(KEYINPUT62), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n891_), .A2(new_n892_), .A3(G169gat), .ZN(new_n893_));
  AOI21_X1  g692(.A(new_n892_), .B1(new_n891_), .B2(G169gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n890_), .B1(new_n893_), .B2(new_n894_), .ZN(G1348gat));
  NAND3_X1  g694(.A1(new_n889_), .A2(new_n525_), .A3(new_n262_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n870_), .A2(new_n884_), .ZN(new_n897_));
  OAI21_X1  g696(.A(G176gat), .B1(new_n897_), .B2(new_n263_), .ZN(new_n898_));
  NAND2_X1  g697(.A1(new_n896_), .A2(new_n898_), .ZN(G1349gat));
  OAI21_X1  g698(.A(new_n509_), .B1(new_n897_), .B2(new_n630_), .ZN(new_n900_));
  OR2_X1    g699(.A1(new_n630_), .A2(new_n326_), .ZN(new_n901_));
  AOI21_X1  g700(.A(new_n901_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n903_));
  OAI21_X1  g702(.A(new_n900_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(new_n904_), .B1(new_n903_), .B2(new_n902_), .ZN(G1350gat));
  INV_X1    g704(.A(KEYINPUT126), .ZN(new_n906_));
  AOI21_X1  g705(.A(new_n511_), .B1(new_n889_), .B2(new_n629_), .ZN(new_n907_));
  NAND2_X1  g706(.A1(new_n615_), .A2(new_n321_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n906_), .B1(new_n907_), .B2(new_n909_), .ZN(new_n910_));
  INV_X1    g709(.A(new_n909_), .ZN(new_n911_));
  AOI21_X1  g710(.A(new_n673_), .B1(new_n886_), .B2(new_n888_), .ZN(new_n912_));
  OAI211_X1 g711(.A(new_n911_), .B(KEYINPUT126), .C1(new_n511_), .C2(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n910_), .A2(new_n913_), .ZN(G1351gat));
  NOR2_X1   g713(.A1(new_n591_), .A2(new_n423_), .ZN(new_n915_));
  OAI211_X1 g714(.A(new_n871_), .B(new_n915_), .C1(new_n849_), .C2(new_n797_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(KEYINPUT127), .ZN(new_n917_));
  INV_X1    g716(.A(KEYINPUT127), .ZN(new_n918_));
  NAND4_X1  g717(.A1(new_n870_), .A2(new_n918_), .A3(new_n871_), .A4(new_n915_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n621_), .B1(new_n917_), .B2(new_n919_), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(new_n440_), .ZN(G1352gat));
  AOI21_X1  g720(.A(new_n263_), .B1(new_n917_), .B2(new_n919_), .ZN(new_n922_));
  XNOR2_X1  g721(.A(new_n922_), .B(new_n437_), .ZN(G1353gat));
  XNOR2_X1  g722(.A(KEYINPUT63), .B(G211gat), .ZN(new_n924_));
  AOI211_X1 g723(.A(new_n630_), .B(new_n924_), .C1(new_n917_), .C2(new_n919_), .ZN(new_n925_));
  NAND2_X1  g724(.A1(new_n917_), .A2(new_n919_), .ZN(new_n926_));
  NAND2_X1  g725(.A1(new_n926_), .A2(new_n314_), .ZN(new_n927_));
  NOR2_X1   g726(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n928_));
  AOI21_X1  g727(.A(new_n925_), .B1(new_n927_), .B2(new_n928_), .ZN(G1354gat));
  NAND3_X1  g728(.A1(new_n926_), .A2(new_n444_), .A3(new_n615_), .ZN(new_n930_));
  AOI21_X1  g729(.A(new_n673_), .B1(new_n917_), .B2(new_n919_), .ZN(new_n931_));
  OAI21_X1  g730(.A(new_n930_), .B1(new_n444_), .B2(new_n931_), .ZN(G1355gat));
endmodule


