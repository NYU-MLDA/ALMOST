//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n725_,
    new_n726_, new_n727_, new_n728_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n823_, new_n824_, new_n825_, new_n826_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n836_, new_n837_, new_n838_, new_n839_, new_n840_,
    new_n841_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n862_,
    new_n863_, new_n865_, new_n866_, new_n867_, new_n868_, new_n869_,
    new_n870_, new_n871_, new_n873_, new_n874_, new_n875_, new_n876_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n903_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n908_, new_n909_, new_n910_, new_n911_, new_n912_, new_n913_,
    new_n914_, new_n915_, new_n916_, new_n917_, new_n918_, new_n919_,
    new_n920_, new_n921_, new_n922_, new_n923_, new_n924_, new_n925_,
    new_n926_, new_n927_, new_n928_, new_n929_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n951_, new_n952_, new_n953_,
    new_n954_, new_n955_, new_n957_, new_n958_, new_n960_, new_n961_,
    new_n962_, new_n964_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n986_, new_n987_, new_n989_, new_n990_,
    new_n992_, new_n993_, new_n994_, new_n996_, new_n997_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1004_, new_n1005_, new_n1006_;
  NAND2_X1  g000(.A1(G230gat), .A2(G233gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT65), .ZN(new_n203_));
  INV_X1    g002(.A(G57gat), .ZN(new_n204_));
  NOR2_X1   g003(.A1(new_n204_), .A2(G64gat), .ZN(new_n205_));
  INV_X1    g004(.A(G64gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(G57gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n203_), .B1(new_n205_), .B2(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n209_));
  NAND2_X1  g008(.A1(new_n206_), .A2(G57gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n204_), .A2(G64gat), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT65), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n208_), .A2(new_n209_), .A3(new_n212_), .ZN(new_n213_));
  XOR2_X1   g012(.A(G71gat), .B(G78gat), .Z(new_n214_));
  NAND2_X1  g013(.A1(new_n213_), .A2(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n208_), .A2(new_n212_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n216_), .B1(new_n217_), .B2(KEYINPUT11), .ZN(new_n218_));
  AOI211_X1 g017(.A(KEYINPUT66), .B(new_n209_), .C1(new_n208_), .C2(new_n212_), .ZN(new_n219_));
  OAI21_X1  g018(.A(new_n215_), .B1(new_n218_), .B2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(new_n214_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n210_), .A2(new_n211_), .A3(KEYINPUT65), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT65), .B1(new_n210_), .B2(new_n211_), .ZN(new_n223_));
  NOR2_X1   g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n221_), .B1(new_n224_), .B2(new_n209_), .ZN(new_n225_));
  OAI21_X1  g024(.A(KEYINPUT11), .B1(new_n222_), .B2(new_n223_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(new_n226_), .A2(KEYINPUT66), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n217_), .A2(new_n216_), .A3(KEYINPUT11), .ZN(new_n228_));
  NAND3_X1  g027(.A1(new_n225_), .A2(new_n227_), .A3(new_n228_), .ZN(new_n229_));
  INV_X1    g028(.A(KEYINPUT7), .ZN(new_n230_));
  INV_X1    g029(.A(G99gat), .ZN(new_n231_));
  INV_X1    g030(.A(G106gat), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n230_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(G99gat), .A2(G106gat), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT6), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n237_));
  OAI21_X1  g036(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n238_));
  NAND4_X1  g037(.A1(new_n233_), .A2(new_n236_), .A3(new_n237_), .A4(new_n238_), .ZN(new_n239_));
  XOR2_X1   g038(.A(G85gat), .B(G92gat), .Z(new_n240_));
  NAND2_X1  g039(.A1(new_n239_), .A2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT8), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT8), .ZN(new_n243_));
  NAND3_X1  g042(.A1(new_n239_), .A2(new_n243_), .A3(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n236_), .A2(new_n237_), .ZN(new_n245_));
  XOR2_X1   g044(.A(KEYINPUT10), .B(G99gat), .Z(new_n246_));
  AOI21_X1  g045(.A(new_n245_), .B1(new_n246_), .B2(new_n232_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(KEYINPUT9), .A2(G85gat), .A3(G92gat), .ZN(new_n248_));
  INV_X1    g047(.A(G85gat), .ZN(new_n249_));
  OR2_X1    g048(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n250_));
  NAND2_X1  g049(.A1(KEYINPUT64), .A2(G92gat), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n249_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  OAI21_X1  g051(.A(KEYINPUT9), .B1(G85gat), .B2(G92gat), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  OAI21_X1  g053(.A(new_n248_), .B1(new_n252_), .B2(new_n254_), .ZN(new_n255_));
  AOI22_X1  g054(.A1(new_n242_), .A2(new_n244_), .B1(new_n247_), .B2(new_n255_), .ZN(new_n256_));
  NAND3_X1  g055(.A1(new_n220_), .A2(new_n229_), .A3(new_n256_), .ZN(new_n257_));
  NAND2_X1  g056(.A1(new_n257_), .A2(KEYINPUT12), .ZN(new_n258_));
  AOI21_X1  g057(.A(new_n256_), .B1(new_n220_), .B2(new_n229_), .ZN(new_n259_));
  NOR2_X1   g058(.A1(new_n258_), .A2(new_n259_), .ZN(new_n260_));
  AOI211_X1 g059(.A(KEYINPUT12), .B(new_n256_), .C1(new_n220_), .C2(new_n229_), .ZN(new_n261_));
  OAI21_X1  g060(.A(new_n202_), .B1(new_n260_), .B2(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n256_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n225_), .B1(new_n227_), .B2(new_n228_), .ZN(new_n264_));
  NOR3_X1   g063(.A1(new_n218_), .A2(new_n219_), .A3(new_n215_), .ZN(new_n265_));
  OAI21_X1  g064(.A(new_n263_), .B1(new_n264_), .B2(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n202_), .B1(new_n266_), .B2(new_n257_), .ZN(new_n267_));
  INV_X1    g066(.A(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n262_), .A2(new_n268_), .ZN(new_n269_));
  XNOR2_X1  g068(.A(G120gat), .B(G148gat), .ZN(new_n270_));
  INV_X1    g069(.A(G204gat), .ZN(new_n271_));
  XNOR2_X1  g070(.A(new_n270_), .B(new_n271_), .ZN(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT5), .B(G176gat), .ZN(new_n273_));
  XOR2_X1   g072(.A(new_n272_), .B(new_n273_), .Z(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  NAND2_X1  g074(.A1(new_n269_), .A2(new_n275_), .ZN(new_n276_));
  XOR2_X1   g075(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n277_));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n278_));
  NAND3_X1  g077(.A1(new_n266_), .A2(KEYINPUT12), .A3(new_n257_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n258_), .A2(new_n259_), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n267_), .B1(new_n281_), .B2(new_n202_), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n278_), .B1(new_n282_), .B2(new_n274_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n202_), .ZN(new_n284_));
  AOI21_X1  g083(.A(new_n284_), .B1(new_n279_), .B2(new_n280_), .ZN(new_n285_));
  NOR4_X1   g084(.A1(new_n285_), .A2(KEYINPUT67), .A3(new_n267_), .A4(new_n275_), .ZN(new_n286_));
  OAI211_X1 g085(.A(new_n276_), .B(new_n277_), .C1(new_n283_), .C2(new_n286_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n262_), .A2(new_n268_), .A3(new_n274_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n288_), .A2(KEYINPUT67), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n282_), .A2(new_n278_), .A3(new_n274_), .ZN(new_n290_));
  AOI22_X1  g089(.A1(new_n289_), .A2(new_n290_), .B1(new_n269_), .B2(new_n275_), .ZN(new_n291_));
  INV_X1    g090(.A(KEYINPUT68), .ZN(new_n292_));
  NOR2_X1   g091(.A1(new_n292_), .A2(KEYINPUT13), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n287_), .B1(new_n291_), .B2(new_n293_), .ZN(new_n294_));
  OR2_X1    g093(.A1(new_n294_), .A2(KEYINPUT69), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n294_), .A2(KEYINPUT69), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n295_), .A2(new_n296_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(G226gat), .A2(G233gat), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n299_), .B(KEYINPUT19), .ZN(new_n300_));
  INV_X1    g099(.A(KEYINPUT20), .ZN(new_n301_));
  NOR2_X1   g100(.A1(new_n300_), .A2(new_n301_), .ZN(new_n302_));
  XNOR2_X1  g101(.A(G211gat), .B(G218gat), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n304_), .A2(KEYINPUT21), .ZN(new_n305_));
  INV_X1    g104(.A(G197gat), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(KEYINPUT83), .ZN(new_n307_));
  INV_X1    g106(.A(KEYINPUT83), .ZN(new_n308_));
  NAND2_X1  g107(.A1(new_n308_), .A2(G197gat), .ZN(new_n309_));
  NAND3_X1  g108(.A1(new_n307_), .A2(new_n309_), .A3(G204gat), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT86), .ZN(new_n311_));
  XNOR2_X1  g110(.A(KEYINPUT84), .B(G204gat), .ZN(new_n312_));
  AOI22_X1  g111(.A1(new_n310_), .A2(new_n311_), .B1(new_n312_), .B2(G197gat), .ZN(new_n313_));
  NAND4_X1  g112(.A1(new_n307_), .A2(new_n309_), .A3(KEYINPUT86), .A4(G204gat), .ZN(new_n314_));
  AOI21_X1  g113(.A(new_n305_), .B1(new_n313_), .B2(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  XNOR2_X1  g115(.A(KEYINPUT83), .B(G197gat), .ZN(new_n317_));
  OAI22_X1  g116(.A1(G197gat), .A2(new_n312_), .B1(new_n317_), .B2(G204gat), .ZN(new_n318_));
  AOI21_X1  g117(.A(KEYINPUT85), .B1(new_n318_), .B2(KEYINPUT21), .ZN(new_n319_));
  AOI21_X1  g118(.A(G204gat), .B1(new_n307_), .B2(new_n309_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n271_), .A2(KEYINPUT84), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT84), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n322_), .A2(G204gat), .ZN(new_n323_));
  AOI21_X1  g122(.A(G197gat), .B1(new_n321_), .B2(new_n323_), .ZN(new_n324_));
  OAI211_X1 g123(.A(KEYINPUT85), .B(KEYINPUT21), .C1(new_n320_), .C2(new_n324_), .ZN(new_n325_));
  INV_X1    g124(.A(new_n325_), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n319_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n310_), .A2(new_n311_), .ZN(new_n328_));
  INV_X1    g127(.A(KEYINPUT21), .ZN(new_n329_));
  NAND2_X1  g128(.A1(new_n312_), .A2(G197gat), .ZN(new_n330_));
  NAND4_X1  g129(.A1(new_n328_), .A2(new_n329_), .A3(new_n314_), .A4(new_n330_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n331_), .A2(new_n303_), .ZN(new_n332_));
  OAI21_X1  g131(.A(new_n316_), .B1(new_n327_), .B2(new_n332_), .ZN(new_n333_));
  INV_X1    g132(.A(G183gat), .ZN(new_n334_));
  INV_X1    g133(.A(G190gat), .ZN(new_n335_));
  OAI21_X1  g134(.A(KEYINPUT23), .B1(new_n334_), .B2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT23), .ZN(new_n337_));
  NAND3_X1  g136(.A1(new_n337_), .A2(G183gat), .A3(G190gat), .ZN(new_n338_));
  NAND2_X1  g137(.A1(new_n336_), .A2(new_n338_), .ZN(new_n339_));
  INV_X1    g138(.A(G169gat), .ZN(new_n340_));
  INV_X1    g139(.A(G176gat), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n340_), .A2(new_n341_), .A3(KEYINPUT79), .ZN(new_n342_));
  INV_X1    g141(.A(KEYINPUT79), .ZN(new_n343_));
  OAI21_X1  g142(.A(new_n343_), .B1(G169gat), .B2(G176gat), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n342_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346_));
  AND2_X1   g145(.A1(KEYINPUT88), .A2(KEYINPUT24), .ZN(new_n347_));
  NOR2_X1   g146(.A1(KEYINPUT88), .A2(KEYINPUT24), .ZN(new_n348_));
  OAI21_X1  g147(.A(new_n346_), .B1(new_n347_), .B2(new_n348_), .ZN(new_n349_));
  OAI21_X1  g148(.A(new_n339_), .B1(new_n345_), .B2(new_n349_), .ZN(new_n350_));
  AOI211_X1 g149(.A(new_n348_), .B(new_n347_), .C1(new_n342_), .C2(new_n344_), .ZN(new_n351_));
  NOR2_X1   g150(.A1(new_n350_), .A2(new_n351_), .ZN(new_n352_));
  NAND2_X1  g151(.A1(new_n334_), .A2(KEYINPUT25), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT25), .ZN(new_n354_));
  NAND2_X1  g153(.A1(new_n354_), .A2(G183gat), .ZN(new_n355_));
  AND2_X1   g154(.A1(new_n353_), .A2(new_n355_), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT26), .B(G190gat), .ZN(new_n357_));
  INV_X1    g156(.A(KEYINPUT87), .ZN(new_n358_));
  AND2_X1   g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  NOR2_X1   g158(.A1(new_n357_), .A2(new_n358_), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n356_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n352_), .A2(new_n361_), .ZN(new_n362_));
  INV_X1    g161(.A(new_n346_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G169gat), .ZN(new_n364_));
  AOI21_X1  g163(.A(new_n363_), .B1(new_n364_), .B2(new_n341_), .ZN(new_n365_));
  AOI21_X1  g164(.A(new_n337_), .B1(G183gat), .B2(G190gat), .ZN(new_n366_));
  NAND2_X1  g165(.A1(new_n338_), .A2(KEYINPUT81), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n368_));
  NAND4_X1  g167(.A1(new_n368_), .A2(new_n337_), .A3(G183gat), .A4(G190gat), .ZN(new_n369_));
  AOI21_X1  g168(.A(new_n366_), .B1(new_n367_), .B2(new_n369_), .ZN(new_n370_));
  NOR2_X1   g169(.A1(G183gat), .A2(G190gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n365_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n372_), .A2(KEYINPUT89), .ZN(new_n373_));
  INV_X1    g172(.A(KEYINPUT89), .ZN(new_n374_));
  OAI211_X1 g173(.A(new_n374_), .B(new_n365_), .C1(new_n370_), .C2(new_n371_), .ZN(new_n375_));
  NAND3_X1  g174(.A1(new_n362_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n376_));
  OAI21_X1  g175(.A(new_n302_), .B1(new_n333_), .B2(new_n376_), .ZN(new_n377_));
  NAND4_X1  g176(.A1(new_n342_), .A2(new_n344_), .A3(KEYINPUT24), .A4(new_n346_), .ZN(new_n378_));
  AND2_X1   g177(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n379_));
  NOR2_X1   g178(.A1(KEYINPUT78), .A2(G190gat), .ZN(new_n380_));
  INV_X1    g179(.A(KEYINPUT26), .ZN(new_n381_));
  NOR3_X1   g180(.A1(new_n379_), .A2(new_n380_), .A3(new_n381_), .ZN(new_n382_));
  OAI211_X1 g181(.A(new_n353_), .B(new_n355_), .C1(KEYINPUT26), .C2(new_n335_), .ZN(new_n383_));
  OAI21_X1  g182(.A(new_n378_), .B1(new_n382_), .B2(new_n383_), .ZN(new_n384_));
  INV_X1    g183(.A(KEYINPUT80), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n384_), .A2(new_n385_), .ZN(new_n386_));
  OAI211_X1 g185(.A(new_n378_), .B(KEYINPUT80), .C1(new_n382_), .C2(new_n383_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(new_n367_), .A2(new_n369_), .ZN(new_n388_));
  INV_X1    g187(.A(KEYINPUT24), .ZN(new_n389_));
  AOI22_X1  g188(.A1(new_n388_), .A2(new_n336_), .B1(new_n389_), .B2(new_n345_), .ZN(new_n390_));
  NAND3_X1  g189(.A1(new_n386_), .A2(new_n387_), .A3(new_n390_), .ZN(new_n391_));
  OR2_X1    g190(.A1(new_n379_), .A2(new_n380_), .ZN(new_n392_));
  OAI21_X1  g191(.A(new_n339_), .B1(new_n392_), .B2(G183gat), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n393_), .A2(new_n365_), .ZN(new_n394_));
  AND2_X1   g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n331_), .A2(new_n303_), .ZN(new_n396_));
  OAI21_X1  g195(.A(KEYINPUT21), .B1(new_n320_), .B2(new_n324_), .ZN(new_n397_));
  INV_X1    g196(.A(KEYINPUT85), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  NAND2_X1  g198(.A1(new_n399_), .A2(new_n325_), .ZN(new_n400_));
  AOI21_X1  g199(.A(new_n315_), .B1(new_n396_), .B2(new_n400_), .ZN(new_n401_));
  OAI21_X1  g200(.A(KEYINPUT91), .B1(new_n395_), .B2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT91), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n391_), .A2(new_n394_), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n333_), .A2(new_n403_), .A3(new_n404_), .ZN(new_n405_));
  AOI21_X1  g204(.A(new_n377_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n300_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n301_), .B1(new_n333_), .B2(new_n376_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n396_), .A2(new_n400_), .ZN(new_n410_));
  NAND4_X1  g209(.A1(new_n410_), .A2(new_n394_), .A3(new_n391_), .A4(new_n316_), .ZN(new_n411_));
  AOI211_X1 g210(.A(KEYINPUT90), .B(new_n408_), .C1(new_n409_), .C2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT90), .ZN(new_n413_));
  AOI21_X1  g212(.A(new_n332_), .B1(new_n399_), .B2(new_n325_), .ZN(new_n414_));
  OAI21_X1  g213(.A(new_n376_), .B1(new_n414_), .B2(new_n315_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n415_), .A2(new_n411_), .A3(KEYINPUT20), .ZN(new_n416_));
  AOI21_X1  g215(.A(new_n413_), .B1(new_n416_), .B2(new_n300_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n407_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n418_));
  XNOR2_X1  g217(.A(G8gat), .B(G36gat), .ZN(new_n419_));
  XNOR2_X1  g218(.A(new_n419_), .B(KEYINPUT18), .ZN(new_n420_));
  XNOR2_X1  g219(.A(new_n420_), .B(G64gat), .ZN(new_n421_));
  INV_X1    g220(.A(G92gat), .ZN(new_n422_));
  XNOR2_X1  g221(.A(new_n421_), .B(new_n422_), .ZN(new_n423_));
  INV_X1    g222(.A(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n418_), .A2(new_n424_), .ZN(new_n425_));
  OAI211_X1 g224(.A(new_n407_), .B(new_n423_), .C1(new_n412_), .C2(new_n417_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT27), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n409_), .A2(new_n408_), .A3(new_n411_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n388_), .A2(new_n336_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n371_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(new_n431_), .ZN(new_n432_));
  AOI22_X1  g231(.A1(new_n352_), .A2(new_n361_), .B1(new_n432_), .B2(new_n365_), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n410_), .A2(new_n433_), .A3(new_n316_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(KEYINPUT20), .ZN(new_n435_));
  AOI21_X1  g234(.A(new_n435_), .B1(new_n402_), .B2(new_n405_), .ZN(new_n436_));
  OAI21_X1  g235(.A(new_n429_), .B1(new_n436_), .B2(new_n408_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n428_), .B1(new_n437_), .B2(new_n424_), .ZN(new_n438_));
  AOI22_X1  g237(.A1(new_n427_), .A2(new_n428_), .B1(new_n426_), .B2(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(KEYINPUT95), .B(KEYINPUT0), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT96), .ZN(new_n441_));
  XNOR2_X1  g240(.A(new_n440_), .B(new_n441_), .ZN(new_n442_));
  XNOR2_X1  g241(.A(G1gat), .B(G29gat), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n440_), .B(KEYINPUT96), .ZN(new_n445_));
  INV_X1    g244(.A(new_n443_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(new_n445_), .A2(new_n446_), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n444_), .A2(new_n447_), .ZN(new_n448_));
  XNOR2_X1  g247(.A(G57gat), .B(G85gat), .ZN(new_n449_));
  INV_X1    g248(.A(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n448_), .A2(new_n450_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n444_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n451_), .A2(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(G225gat), .A2(G233gat), .ZN(new_n454_));
  XNOR2_X1  g253(.A(new_n454_), .B(KEYINPUT93), .ZN(new_n455_));
  INV_X1    g254(.A(new_n455_), .ZN(new_n456_));
  INV_X1    g255(.A(G134gat), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(G127gat), .ZN(new_n458_));
  INV_X1    g257(.A(G127gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(G134gat), .ZN(new_n460_));
  INV_X1    g259(.A(G120gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(new_n461_), .A2(G113gat), .ZN(new_n462_));
  INV_X1    g261(.A(G113gat), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n463_), .A2(G120gat), .ZN(new_n464_));
  NAND4_X1  g263(.A1(new_n458_), .A2(new_n460_), .A3(new_n462_), .A4(new_n464_), .ZN(new_n465_));
  NAND2_X1  g264(.A1(new_n458_), .A2(new_n460_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n462_), .A2(new_n464_), .ZN(new_n467_));
  NAND2_X1  g266(.A1(new_n466_), .A2(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(G155gat), .B(G162gat), .ZN(new_n469_));
  INV_X1    g268(.A(G141gat), .ZN(new_n470_));
  INV_X1    g269(.A(G148gat), .ZN(new_n471_));
  NAND3_X1  g270(.A1(new_n470_), .A2(new_n471_), .A3(KEYINPUT3), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT3), .ZN(new_n473_));
  OAI21_X1  g272(.A(new_n473_), .B1(G141gat), .B2(G148gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  AND3_X1   g274(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n476_));
  AOI21_X1  g275(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n477_));
  NOR2_X1   g276(.A1(new_n476_), .A2(new_n477_), .ZN(new_n478_));
  AOI21_X1  g277(.A(new_n469_), .B1(new_n475_), .B2(new_n478_), .ZN(new_n479_));
  AND2_X1   g278(.A1(G155gat), .A2(G162gat), .ZN(new_n480_));
  NOR2_X1   g279(.A1(G155gat), .A2(G162gat), .ZN(new_n481_));
  NOR3_X1   g280(.A1(new_n480_), .A2(new_n481_), .A3(KEYINPUT1), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n470_), .A2(new_n471_), .ZN(new_n483_));
  NAND2_X1  g282(.A1(G141gat), .A2(G148gat), .ZN(new_n484_));
  NAND3_X1  g283(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n485_));
  NAND3_X1  g284(.A1(new_n483_), .A2(new_n484_), .A3(new_n485_), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n482_), .A2(new_n486_), .ZN(new_n487_));
  OAI211_X1 g286(.A(new_n465_), .B(new_n468_), .C1(new_n479_), .C2(new_n487_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(KEYINPUT94), .B(KEYINPUT4), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  INV_X1    g289(.A(new_n469_), .ZN(new_n491_));
  AND2_X1   g290(.A1(new_n472_), .A2(new_n474_), .ZN(new_n492_));
  INV_X1    g291(.A(new_n477_), .ZN(new_n493_));
  NAND3_X1  g292(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n494_));
  NAND2_X1  g293(.A1(new_n493_), .A2(new_n494_), .ZN(new_n495_));
  OAI21_X1  g294(.A(new_n491_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  AND2_X1   g295(.A1(new_n483_), .A2(new_n484_), .ZN(new_n497_));
  OAI211_X1 g296(.A(new_n497_), .B(new_n485_), .C1(KEYINPUT1), .C2(new_n469_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n468_), .A2(new_n465_), .ZN(new_n499_));
  NAND3_X1  g298(.A1(new_n496_), .A2(new_n498_), .A3(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(new_n488_), .A2(new_n500_), .A3(KEYINPUT4), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT92), .ZN(new_n502_));
  NAND2_X1  g301(.A1(new_n501_), .A2(new_n502_), .ZN(new_n503_));
  NAND4_X1  g302(.A1(new_n488_), .A2(new_n500_), .A3(KEYINPUT92), .A4(KEYINPUT4), .ZN(new_n504_));
  AOI211_X1 g303(.A(new_n456_), .B(new_n490_), .C1(new_n503_), .C2(new_n504_), .ZN(new_n505_));
  AND2_X1   g304(.A1(new_n488_), .A2(new_n500_), .ZN(new_n506_));
  AND2_X1   g305(.A1(new_n506_), .A2(new_n454_), .ZN(new_n507_));
  OAI21_X1  g306(.A(new_n453_), .B1(new_n505_), .B2(new_n507_), .ZN(new_n508_));
  AOI21_X1  g307(.A(new_n490_), .B1(new_n503_), .B2(new_n504_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n509_), .A2(new_n455_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n453_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n507_), .ZN(new_n512_));
  NAND3_X1  g311(.A1(new_n510_), .A2(new_n511_), .A3(new_n512_), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n508_), .A2(new_n513_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(G71gat), .B(G99gat), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G227gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n515_), .B(new_n516_), .ZN(new_n517_));
  AND3_X1   g316(.A1(new_n391_), .A2(KEYINPUT30), .A3(new_n394_), .ZN(new_n518_));
  AOI21_X1  g317(.A(KEYINPUT30), .B1(new_n391_), .B2(new_n394_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n517_), .B1(new_n518_), .B2(new_n519_), .ZN(new_n520_));
  INV_X1    g319(.A(KEYINPUT30), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n404_), .A2(new_n521_), .ZN(new_n522_));
  NAND3_X1  g321(.A1(new_n391_), .A2(KEYINPUT30), .A3(new_n394_), .ZN(new_n523_));
  INV_X1    g322(.A(new_n517_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n522_), .A2(new_n523_), .A3(new_n524_), .ZN(new_n525_));
  XNOR2_X1  g324(.A(G15gat), .B(G43gat), .ZN(new_n526_));
  AND3_X1   g325(.A1(new_n520_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n527_));
  AOI21_X1  g326(.A(new_n526_), .B1(new_n520_), .B2(new_n525_), .ZN(new_n528_));
  XOR2_X1   g327(.A(new_n499_), .B(KEYINPUT31), .Z(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NOR3_X1   g329(.A1(new_n527_), .A2(new_n528_), .A3(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n526_), .ZN(new_n532_));
  NOR3_X1   g331(.A1(new_n518_), .A2(new_n519_), .A3(new_n517_), .ZN(new_n533_));
  AOI21_X1  g332(.A(new_n524_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n534_));
  OAI21_X1  g333(.A(new_n532_), .B1(new_n533_), .B2(new_n534_), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n520_), .A2(new_n525_), .A3(new_n526_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n529_), .B1(new_n535_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(G233gat), .ZN(new_n538_));
  INV_X1    g337(.A(KEYINPUT82), .ZN(new_n539_));
  NOR2_X1   g338(.A1(new_n539_), .A2(G228gat), .ZN(new_n540_));
  INV_X1    g339(.A(new_n540_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n539_), .A2(G228gat), .ZN(new_n542_));
  AOI21_X1  g341(.A(new_n538_), .B1(new_n541_), .B2(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  NOR2_X1   g343(.A1(new_n479_), .A2(new_n487_), .ZN(new_n545_));
  INV_X1    g344(.A(KEYINPUT29), .ZN(new_n546_));
  NOR2_X1   g345(.A1(new_n545_), .A2(new_n546_), .ZN(new_n547_));
  INV_X1    g346(.A(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n333_), .A2(new_n544_), .A3(new_n548_), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n543_), .B1(new_n401_), .B2(new_n547_), .ZN(new_n550_));
  XNOR2_X1  g349(.A(G78gat), .B(G106gat), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n549_), .A2(new_n550_), .A3(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(new_n552_), .B1(new_n549_), .B2(new_n550_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n545_), .A2(new_n546_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G22gat), .B(G50gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT28), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n556_), .B(new_n558_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  NOR3_X1   g359(.A1(new_n554_), .A2(new_n555_), .A3(new_n560_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n549_), .A2(new_n550_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(new_n551_), .ZN(new_n563_));
  AOI21_X1  g362(.A(new_n559_), .B1(new_n563_), .B2(new_n553_), .ZN(new_n564_));
  OAI22_X1  g363(.A1(new_n531_), .A2(new_n537_), .B1(new_n561_), .B2(new_n564_), .ZN(new_n565_));
  OAI21_X1  g364(.A(new_n530_), .B1(new_n527_), .B2(new_n528_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n560_), .B1(new_n554_), .B2(new_n555_), .ZN(new_n567_));
  NAND3_X1  g366(.A1(new_n535_), .A2(new_n536_), .A3(new_n529_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n563_), .A2(new_n559_), .A3(new_n553_), .ZN(new_n569_));
  NAND4_X1  g368(.A1(new_n566_), .A2(new_n567_), .A3(new_n568_), .A4(new_n569_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n514_), .B1(new_n565_), .B2(new_n570_), .ZN(new_n571_));
  INV_X1    g370(.A(KEYINPUT33), .ZN(new_n572_));
  AOI211_X1 g371(.A(new_n453_), .B(new_n507_), .C1(new_n509_), .C2(new_n455_), .ZN(new_n573_));
  OAI21_X1  g372(.A(new_n572_), .B1(new_n573_), .B2(KEYINPUT97), .ZN(new_n574_));
  INV_X1    g373(.A(KEYINPUT97), .ZN(new_n575_));
  NAND3_X1  g374(.A1(new_n513_), .A2(new_n575_), .A3(KEYINPUT33), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n574_), .A2(new_n576_), .ZN(new_n577_));
  NAND2_X1  g376(.A1(new_n509_), .A2(new_n454_), .ZN(new_n578_));
  NAND2_X1  g377(.A1(new_n506_), .A2(new_n455_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n578_), .A2(new_n453_), .A3(new_n579_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n425_), .A2(new_n577_), .A3(new_n426_), .A4(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n402_), .A2(new_n405_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n377_), .ZN(new_n583_));
  AOI22_X1  g382(.A1(new_n582_), .A2(new_n583_), .B1(KEYINPUT32), .B2(new_n423_), .ZN(new_n584_));
  OAI21_X1  g383(.A(new_n584_), .B1(new_n412_), .B2(new_n417_), .ZN(new_n585_));
  INV_X1    g384(.A(KEYINPUT98), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n585_), .A2(new_n586_), .ZN(new_n587_));
  AND2_X1   g386(.A1(new_n423_), .A2(KEYINPUT32), .ZN(new_n588_));
  AOI22_X1  g387(.A1(new_n437_), .A2(new_n588_), .B1(new_n513_), .B2(new_n508_), .ZN(new_n589_));
  AND3_X1   g388(.A1(new_n362_), .A2(new_n373_), .A3(new_n375_), .ZN(new_n590_));
  OAI21_X1  g389(.A(KEYINPUT20), .B1(new_n590_), .B2(new_n401_), .ZN(new_n591_));
  NOR2_X1   g390(.A1(new_n333_), .A2(new_n404_), .ZN(new_n592_));
  OAI21_X1  g391(.A(new_n300_), .B1(new_n591_), .B2(new_n592_), .ZN(new_n593_));
  NAND2_X1  g392(.A1(new_n593_), .A2(KEYINPUT90), .ZN(new_n594_));
  NAND3_X1  g393(.A1(new_n416_), .A2(new_n413_), .A3(new_n300_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(new_n594_), .A2(new_n595_), .ZN(new_n596_));
  NAND3_X1  g395(.A1(new_n596_), .A2(KEYINPUT98), .A3(new_n584_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n587_), .A2(new_n589_), .A3(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n581_), .A2(new_n598_), .ZN(new_n599_));
  NOR2_X1   g398(.A1(new_n531_), .A2(new_n537_), .ZN(new_n600_));
  NAND2_X1  g399(.A1(new_n567_), .A2(new_n569_), .ZN(new_n601_));
  NOR2_X1   g400(.A1(new_n600_), .A2(new_n601_), .ZN(new_n602_));
  AOI22_X1  g401(.A1(new_n439_), .A2(new_n571_), .B1(new_n599_), .B2(new_n602_), .ZN(new_n603_));
  NOR2_X1   g402(.A1(new_n264_), .A2(new_n265_), .ZN(new_n604_));
  NAND2_X1  g403(.A1(G1gat), .A2(G8gat), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n605_), .A2(KEYINPUT14), .ZN(new_n606_));
  NOR2_X1   g405(.A1(G15gat), .A2(G22gat), .ZN(new_n607_));
  AND2_X1   g406(.A1(G15gat), .A2(G22gat), .ZN(new_n608_));
  OAI21_X1  g407(.A(new_n606_), .B1(new_n607_), .B2(new_n608_), .ZN(new_n609_));
  OR2_X1    g408(.A1(new_n609_), .A2(KEYINPUT75), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n609_), .A2(KEYINPUT75), .ZN(new_n611_));
  NAND2_X1  g410(.A1(new_n610_), .A2(new_n611_), .ZN(new_n612_));
  XOR2_X1   g411(.A(G1gat), .B(G8gat), .Z(new_n613_));
  INV_X1    g412(.A(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n612_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n610_), .A2(new_n613_), .A3(new_n611_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n604_), .A2(new_n617_), .ZN(new_n618_));
  NOR2_X1   g417(.A1(new_n604_), .A2(new_n617_), .ZN(new_n619_));
  INV_X1    g418(.A(G231gat), .ZN(new_n620_));
  NOR2_X1   g419(.A1(new_n620_), .A2(new_n538_), .ZN(new_n621_));
  OR3_X1    g420(.A1(new_n618_), .A2(new_n619_), .A3(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(KEYINPUT76), .B(KEYINPUT16), .ZN(new_n623_));
  XNOR2_X1  g422(.A(G127gat), .B(G155gat), .ZN(new_n624_));
  XNOR2_X1  g423(.A(new_n623_), .B(new_n624_), .ZN(new_n625_));
  XNOR2_X1  g424(.A(G183gat), .B(G211gat), .ZN(new_n626_));
  XNOR2_X1  g425(.A(new_n625_), .B(new_n626_), .ZN(new_n627_));
  OAI21_X1  g426(.A(new_n621_), .B1(new_n618_), .B2(new_n619_), .ZN(new_n628_));
  AND4_X1   g427(.A1(KEYINPUT17), .A2(new_n622_), .A3(new_n627_), .A4(new_n628_), .ZN(new_n629_));
  XNOR2_X1  g428(.A(new_n627_), .B(KEYINPUT17), .ZN(new_n630_));
  AOI21_X1  g429(.A(new_n630_), .B1(new_n622_), .B2(new_n628_), .ZN(new_n631_));
  NOR2_X1   g430(.A1(new_n629_), .A2(new_n631_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT77), .ZN(new_n633_));
  XOR2_X1   g432(.A(G29gat), .B(G36gat), .Z(new_n634_));
  XOR2_X1   g433(.A(G43gat), .B(G50gat), .Z(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n617_), .A2(new_n636_), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n634_), .B(new_n635_), .Z(new_n638_));
  NAND2_X1  g437(.A1(new_n638_), .A2(KEYINPUT15), .ZN(new_n639_));
  INV_X1    g438(.A(KEYINPUT15), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n636_), .A2(new_n640_), .ZN(new_n641_));
  NAND4_X1  g440(.A1(new_n639_), .A2(new_n616_), .A3(new_n615_), .A4(new_n641_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n637_), .A2(new_n642_), .ZN(new_n643_));
  NAND2_X1  g442(.A1(G229gat), .A2(G233gat), .ZN(new_n644_));
  INV_X1    g443(.A(new_n644_), .ZN(new_n645_));
  OAI21_X1  g444(.A(new_n633_), .B1(new_n643_), .B2(new_n645_), .ZN(new_n646_));
  NAND4_X1  g445(.A1(new_n637_), .A2(new_n642_), .A3(KEYINPUT77), .A4(new_n644_), .ZN(new_n647_));
  INV_X1    g446(.A(new_n637_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n617_), .A2(new_n636_), .ZN(new_n649_));
  OAI21_X1  g448(.A(new_n645_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n650_));
  NAND3_X1  g449(.A1(new_n646_), .A2(new_n647_), .A3(new_n650_), .ZN(new_n651_));
  XNOR2_X1  g450(.A(G113gat), .B(G141gat), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(G169gat), .ZN(new_n653_));
  XNOR2_X1  g452(.A(new_n653_), .B(new_n306_), .ZN(new_n654_));
  INV_X1    g453(.A(new_n654_), .ZN(new_n655_));
  NAND2_X1  g454(.A1(new_n651_), .A2(new_n655_), .ZN(new_n656_));
  NAND4_X1  g455(.A1(new_n646_), .A2(new_n650_), .A3(new_n647_), .A4(new_n654_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n632_), .A2(new_n658_), .ZN(new_n659_));
  XOR2_X1   g458(.A(G190gat), .B(G218gat), .Z(new_n660_));
  XNOR2_X1  g459(.A(G134gat), .B(G162gat), .ZN(new_n661_));
  XNOR2_X1  g460(.A(new_n660_), .B(new_n661_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT36), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n256_), .A2(new_n636_), .ZN(new_n664_));
  INV_X1    g463(.A(KEYINPUT72), .ZN(new_n665_));
  NAND2_X1  g464(.A1(G232gat), .A2(G233gat), .ZN(new_n666_));
  XOR2_X1   g465(.A(new_n666_), .B(KEYINPUT70), .Z(new_n667_));
  XNOR2_X1  g466(.A(new_n667_), .B(KEYINPUT34), .ZN(new_n668_));
  INV_X1    g467(.A(KEYINPUT35), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n665_), .B1(new_n668_), .B2(new_n669_), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n639_), .A2(new_n641_), .ZN(new_n671_));
  OAI211_X1 g470(.A(new_n664_), .B(new_n670_), .C1(new_n671_), .C2(new_n256_), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n668_), .A2(new_n669_), .ZN(new_n673_));
  AND2_X1   g472(.A1(new_n672_), .A2(new_n673_), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n672_), .A2(new_n673_), .ZN(new_n675_));
  OAI21_X1  g474(.A(new_n663_), .B1(new_n674_), .B2(new_n675_), .ZN(new_n676_));
  OR2_X1    g475(.A1(new_n672_), .A2(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n672_), .A2(new_n673_), .ZN(new_n678_));
  INV_X1    g477(.A(KEYINPUT36), .ZN(new_n679_));
  NAND2_X1  g478(.A1(new_n662_), .A2(new_n679_), .ZN(new_n680_));
  XNOR2_X1  g479(.A(new_n680_), .B(KEYINPUT71), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n677_), .A2(new_n678_), .A3(new_n681_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT37), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n676_), .A2(new_n682_), .A3(new_n683_), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT74), .ZN(new_n685_));
  XNOR2_X1  g484(.A(new_n684_), .B(new_n685_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n682_), .A2(KEYINPUT73), .ZN(new_n687_));
  NAND2_X1  g486(.A1(new_n687_), .A2(new_n676_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n682_), .A2(KEYINPUT73), .ZN(new_n689_));
  OAI21_X1  g488(.A(KEYINPUT37), .B1(new_n688_), .B2(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n686_), .A2(new_n690_), .ZN(new_n691_));
  INV_X1    g490(.A(new_n691_), .ZN(new_n692_));
  OR4_X1    g491(.A1(new_n298_), .A2(new_n603_), .A3(new_n659_), .A4(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT99), .ZN(new_n694_));
  INV_X1    g493(.A(G1gat), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n694_), .A2(new_n695_), .A3(new_n514_), .ZN(new_n696_));
  INV_X1    g495(.A(KEYINPUT38), .ZN(new_n697_));
  OR2_X1    g496(.A1(new_n696_), .A2(new_n697_), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n599_), .A2(new_n602_), .ZN(new_n699_));
  AOI21_X1  g498(.A(new_n423_), .B1(new_n596_), .B2(new_n407_), .ZN(new_n700_));
  AOI211_X1 g499(.A(new_n424_), .B(new_n406_), .C1(new_n594_), .C2(new_n595_), .ZN(new_n701_));
  OAI21_X1  g500(.A(new_n428_), .B1(new_n700_), .B2(new_n701_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n565_), .A2(new_n570_), .ZN(new_n703_));
  INV_X1    g502(.A(new_n514_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n438_), .A2(new_n426_), .ZN(new_n705_));
  NAND4_X1  g504(.A1(new_n702_), .A2(new_n703_), .A3(new_n704_), .A4(new_n705_), .ZN(new_n706_));
  NAND2_X1  g505(.A1(new_n699_), .A2(new_n706_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n676_), .A2(new_n682_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n707_), .A2(new_n708_), .ZN(new_n709_));
  XNOR2_X1  g508(.A(new_n709_), .B(KEYINPUT100), .ZN(new_n710_));
  INV_X1    g509(.A(new_n294_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(new_n711_), .A2(new_n659_), .ZN(new_n712_));
  NAND2_X1  g511(.A1(new_n710_), .A2(new_n712_), .ZN(new_n713_));
  OAI21_X1  g512(.A(G1gat), .B1(new_n713_), .B2(new_n704_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n696_), .A2(new_n697_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n698_), .A2(new_n714_), .A3(new_n715_), .ZN(G1324gat));
  INV_X1    g515(.A(G8gat), .ZN(new_n717_));
  INV_X1    g516(.A(new_n439_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n694_), .A2(new_n717_), .A3(new_n718_), .ZN(new_n719_));
  OAI21_X1  g518(.A(G8gat), .B1(new_n713_), .B2(new_n439_), .ZN(new_n720_));
  AND2_X1   g519(.A1(new_n720_), .A2(KEYINPUT39), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n720_), .A2(KEYINPUT39), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n719_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  XOR2_X1   g522(.A(new_n723_), .B(KEYINPUT40), .Z(G1325gat));
  INV_X1    g523(.A(new_n600_), .ZN(new_n725_));
  OAI21_X1  g524(.A(G15gat), .B1(new_n713_), .B2(new_n725_), .ZN(new_n726_));
  XOR2_X1   g525(.A(new_n726_), .B(KEYINPUT41), .Z(new_n727_));
  OR2_X1    g526(.A1(new_n725_), .A2(G15gat), .ZN(new_n728_));
  OAI21_X1  g527(.A(new_n727_), .B1(new_n693_), .B2(new_n728_), .ZN(G1326gat));
  INV_X1    g528(.A(new_n601_), .ZN(new_n730_));
  OR3_X1    g529(.A1(new_n693_), .A2(G22gat), .A3(new_n730_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G22gat), .B1(new_n713_), .B2(new_n730_), .ZN(new_n732_));
  AND2_X1   g531(.A1(new_n732_), .A2(KEYINPUT42), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(KEYINPUT42), .ZN(new_n734_));
  OAI21_X1  g533(.A(new_n731_), .B1(new_n733_), .B2(new_n734_), .ZN(new_n735_));
  XOR2_X1   g534(.A(new_n735_), .B(KEYINPUT101), .Z(G1327gat));
  NOR2_X1   g535(.A1(new_n603_), .A2(new_n708_), .ZN(new_n737_));
  OAI21_X1  g536(.A(new_n658_), .B1(new_n629_), .B2(new_n631_), .ZN(new_n738_));
  NOR2_X1   g537(.A1(new_n711_), .A2(new_n738_), .ZN(new_n739_));
  AND2_X1   g538(.A1(new_n737_), .A2(new_n739_), .ZN(new_n740_));
  INV_X1    g539(.A(new_n740_), .ZN(new_n741_));
  OR3_X1    g540(.A1(new_n741_), .A2(G29gat), .A3(new_n704_), .ZN(new_n742_));
  INV_X1    g541(.A(new_n738_), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT102), .B1(new_n294_), .B2(new_n743_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  NAND3_X1  g544(.A1(new_n294_), .A2(KEYINPUT102), .A3(new_n743_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n745_), .A2(new_n746_), .ZN(new_n747_));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n748_));
  AOI21_X1  g547(.A(new_n748_), .B1(new_n707_), .B2(new_n692_), .ZN(new_n749_));
  AOI211_X1 g548(.A(KEYINPUT43), .B(new_n691_), .C1(new_n699_), .C2(new_n706_), .ZN(new_n750_));
  OAI21_X1  g549(.A(new_n747_), .B1(new_n749_), .B2(new_n750_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT105), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT44), .ZN(new_n753_));
  NOR3_X1   g552(.A1(new_n751_), .A2(new_n752_), .A3(new_n753_), .ZN(new_n754_));
  INV_X1    g553(.A(KEYINPUT102), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n276_), .B1(new_n283_), .B2(new_n286_), .ZN(new_n756_));
  INV_X1    g555(.A(new_n293_), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  AOI211_X1 g557(.A(new_n755_), .B(new_n738_), .C1(new_n758_), .C2(new_n287_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(new_n744_), .ZN(new_n760_));
  OAI21_X1  g559(.A(KEYINPUT43), .B1(new_n603_), .B2(new_n691_), .ZN(new_n761_));
  NAND3_X1  g560(.A1(new_n707_), .A2(new_n748_), .A3(new_n692_), .ZN(new_n762_));
  AOI21_X1  g561(.A(new_n760_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n763_));
  AOI21_X1  g562(.A(KEYINPUT105), .B1(new_n763_), .B2(KEYINPUT44), .ZN(new_n764_));
  OAI21_X1  g563(.A(new_n514_), .B1(new_n754_), .B2(new_n764_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n753_), .B1(new_n763_), .B2(KEYINPUT103), .ZN(new_n766_));
  INV_X1    g565(.A(KEYINPUT103), .ZN(new_n767_));
  AOI211_X1 g566(.A(new_n767_), .B(new_n760_), .C1(new_n761_), .C2(new_n762_), .ZN(new_n768_));
  OAI21_X1  g567(.A(KEYINPUT104), .B1(new_n766_), .B2(new_n768_), .ZN(new_n769_));
  AOI21_X1  g568(.A(KEYINPUT44), .B1(new_n751_), .B2(new_n767_), .ZN(new_n770_));
  INV_X1    g569(.A(KEYINPUT104), .ZN(new_n771_));
  NAND2_X1  g570(.A1(new_n763_), .A2(KEYINPUT103), .ZN(new_n772_));
  NAND3_X1  g571(.A1(new_n770_), .A2(new_n771_), .A3(new_n772_), .ZN(new_n773_));
  AOI21_X1  g572(.A(new_n765_), .B1(new_n769_), .B2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT106), .ZN(new_n775_));
  OAI21_X1  g574(.A(G29gat), .B1(new_n774_), .B2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n769_), .A2(new_n773_), .ZN(new_n777_));
  OAI21_X1  g576(.A(new_n752_), .B1(new_n751_), .B2(new_n753_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n763_), .A2(KEYINPUT105), .A3(KEYINPUT44), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n777_), .A2(new_n775_), .A3(new_n780_), .A4(new_n514_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n781_), .ZN(new_n782_));
  OAI21_X1  g581(.A(new_n742_), .B1(new_n776_), .B2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  OAI211_X1 g584(.A(KEYINPUT107), .B(new_n742_), .C1(new_n776_), .C2(new_n782_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n785_), .A2(new_n786_), .ZN(G1328gat));
  INV_X1    g586(.A(KEYINPUT46), .ZN(new_n788_));
  INV_X1    g587(.A(G36gat), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n740_), .A2(new_n789_), .A3(new_n718_), .ZN(new_n790_));
  XOR2_X1   g589(.A(new_n790_), .B(KEYINPUT45), .Z(new_n791_));
  AOI21_X1  g590(.A(new_n439_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n766_), .A2(new_n768_), .A3(KEYINPUT104), .ZN(new_n793_));
  AOI21_X1  g592(.A(new_n771_), .B1(new_n770_), .B2(new_n772_), .ZN(new_n794_));
  OAI21_X1  g593(.A(new_n792_), .B1(new_n793_), .B2(new_n794_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n791_), .B1(new_n795_), .B2(G36gat), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT108), .ZN(new_n797_));
  OAI211_X1 g596(.A(KEYINPUT109), .B(new_n788_), .C1(new_n796_), .C2(new_n797_), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT109), .ZN(new_n799_));
  INV_X1    g598(.A(new_n791_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n718_), .B1(new_n754_), .B2(new_n764_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n801_), .B1(new_n769_), .B2(new_n773_), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n800_), .B1(new_n802_), .B2(new_n789_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n799_), .B1(new_n803_), .B2(KEYINPUT108), .ZN(new_n804_));
  OAI21_X1  g603(.A(KEYINPUT46), .B1(new_n796_), .B2(KEYINPUT109), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n798_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  INV_X1    g605(.A(new_n806_), .ZN(G1329gat));
  INV_X1    g606(.A(G43gat), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n808_), .B1(new_n741_), .B2(new_n725_), .ZN(new_n809_));
  AOI211_X1 g608(.A(new_n808_), .B(new_n725_), .C1(new_n778_), .C2(new_n779_), .ZN(new_n810_));
  NAND3_X1  g609(.A1(new_n777_), .A2(new_n810_), .A3(KEYINPUT110), .ZN(new_n811_));
  INV_X1    g610(.A(new_n811_), .ZN(new_n812_));
  AOI21_X1  g611(.A(KEYINPUT110), .B1(new_n777_), .B2(new_n810_), .ZN(new_n813_));
  OAI21_X1  g612(.A(new_n809_), .B1(new_n812_), .B2(new_n813_), .ZN(new_n814_));
  XNOR2_X1  g613(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n814_), .B(new_n816_), .ZN(G1330gat));
  AND3_X1   g616(.A1(new_n777_), .A2(new_n601_), .A3(new_n780_), .ZN(new_n818_));
  INV_X1    g617(.A(G50gat), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n601_), .A2(new_n819_), .ZN(new_n820_));
  XOR2_X1   g619(.A(new_n820_), .B(KEYINPUT112), .Z(new_n821_));
  OAI22_X1  g620(.A1(new_n818_), .A2(new_n819_), .B1(new_n741_), .B2(new_n821_), .ZN(G1331gat));
  INV_X1    g621(.A(new_n658_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n298_), .A2(new_n823_), .ZN(new_n824_));
  INV_X1    g623(.A(new_n632_), .ZN(new_n825_));
  NOR2_X1   g624(.A1(new_n824_), .A2(new_n825_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n710_), .ZN(new_n827_));
  INV_X1    g626(.A(new_n827_), .ZN(new_n828_));
  OAI21_X1  g627(.A(KEYINPUT113), .B1(new_n704_), .B2(new_n204_), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  NAND4_X1  g629(.A1(new_n711_), .A2(new_n823_), .A3(new_n632_), .A4(new_n691_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n831_), .A2(new_n603_), .ZN(new_n832_));
  NAND3_X1  g631(.A1(new_n830_), .A2(new_n514_), .A3(new_n832_), .ZN(new_n833_));
  INV_X1    g632(.A(new_n830_), .ZN(new_n834_));
  AOI22_X1  g633(.A1(new_n833_), .A2(new_n204_), .B1(new_n834_), .B2(KEYINPUT113), .ZN(G1332gat));
  NAND3_X1  g634(.A1(new_n832_), .A2(new_n206_), .A3(new_n718_), .ZN(new_n836_));
  OAI21_X1  g635(.A(G64gat), .B1(new_n827_), .B2(new_n439_), .ZN(new_n837_));
  OR2_X1    g636(.A1(new_n837_), .A2(KEYINPUT114), .ZN(new_n838_));
  NAND2_X1  g637(.A1(new_n837_), .A2(KEYINPUT114), .ZN(new_n839_));
  AND3_X1   g638(.A1(new_n838_), .A2(KEYINPUT48), .A3(new_n839_), .ZN(new_n840_));
  AOI21_X1  g639(.A(KEYINPUT48), .B1(new_n838_), .B2(new_n839_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n836_), .B1(new_n840_), .B2(new_n841_), .ZN(G1333gat));
  INV_X1    g641(.A(new_n832_), .ZN(new_n843_));
  OR3_X1    g642(.A1(new_n843_), .A2(G71gat), .A3(new_n725_), .ZN(new_n844_));
  OAI21_X1  g643(.A(G71gat), .B1(new_n827_), .B2(new_n725_), .ZN(new_n845_));
  OR2_X1    g644(.A1(new_n845_), .A2(KEYINPUT115), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(KEYINPUT115), .ZN(new_n847_));
  AND3_X1   g646(.A1(new_n846_), .A2(KEYINPUT49), .A3(new_n847_), .ZN(new_n848_));
  AOI21_X1  g647(.A(KEYINPUT49), .B1(new_n846_), .B2(new_n847_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n844_), .B1(new_n848_), .B2(new_n849_), .ZN(G1334gat));
  OAI21_X1  g649(.A(G78gat), .B1(new_n827_), .B2(new_n730_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(new_n851_), .B(KEYINPUT50), .ZN(new_n852_));
  OR2_X1    g651(.A1(new_n730_), .A2(G78gat), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n843_), .B2(new_n853_), .ZN(G1335gat));
  NAND3_X1  g653(.A1(new_n711_), .A2(new_n823_), .A3(new_n825_), .ZN(new_n855_));
  AOI21_X1  g654(.A(new_n855_), .B1(new_n761_), .B2(new_n762_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n249_), .B1(new_n856_), .B2(new_n514_), .ZN(new_n857_));
  NOR4_X1   g656(.A1(new_n824_), .A2(new_n603_), .A3(new_n632_), .A4(new_n708_), .ZN(new_n858_));
  NOR2_X1   g657(.A1(new_n704_), .A2(G85gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(new_n857_), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  XOR2_X1   g659(.A(new_n860_), .B(KEYINPUT116), .Z(G1336gat));
  AOI21_X1  g660(.A(G92gat), .B1(new_n858_), .B2(new_n718_), .ZN(new_n862_));
  AOI21_X1  g661(.A(new_n439_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n863_));
  AOI21_X1  g662(.A(new_n862_), .B1(new_n856_), .B2(new_n863_), .ZN(G1337gat));
  AOI21_X1  g663(.A(new_n231_), .B1(new_n856_), .B2(new_n600_), .ZN(new_n865_));
  XOR2_X1   g664(.A(new_n865_), .B(KEYINPUT117), .Z(new_n866_));
  AND2_X1   g665(.A1(new_n600_), .A2(new_n246_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT118), .ZN(new_n868_));
  AOI22_X1  g667(.A1(new_n858_), .A2(new_n867_), .B1(new_n868_), .B2(KEYINPUT51), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n866_), .A2(new_n869_), .ZN(new_n870_));
  NOR2_X1   g669(.A1(new_n868_), .A2(KEYINPUT51), .ZN(new_n871_));
  XOR2_X1   g670(.A(new_n870_), .B(new_n871_), .Z(G1338gat));
  AOI21_X1  g671(.A(new_n232_), .B1(new_n856_), .B2(new_n601_), .ZN(new_n873_));
  XOR2_X1   g672(.A(new_n873_), .B(KEYINPUT52), .Z(new_n874_));
  NAND3_X1  g673(.A1(new_n858_), .A2(new_n232_), .A3(new_n601_), .ZN(new_n875_));
  NAND2_X1  g674(.A1(new_n874_), .A2(new_n875_), .ZN(new_n876_));
  XNOR2_X1  g675(.A(new_n876_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g676(.A1(new_n730_), .A2(new_n600_), .A3(new_n514_), .ZN(new_n878_));
  NOR2_X1   g677(.A1(new_n718_), .A2(new_n878_), .ZN(new_n879_));
  INV_X1    g678(.A(new_n879_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n643_), .A2(KEYINPUT121), .ZN(new_n881_));
  NOR2_X1   g680(.A1(new_n643_), .A2(KEYINPUT121), .ZN(new_n882_));
  NOR3_X1   g681(.A1(new_n881_), .A2(new_n882_), .A3(new_n644_), .ZN(new_n883_));
  OAI21_X1  g682(.A(new_n644_), .B1(new_n648_), .B2(new_n649_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n655_), .ZN(new_n885_));
  OAI21_X1  g684(.A(new_n657_), .B1(new_n883_), .B2(new_n885_), .ZN(new_n886_));
  NOR2_X1   g685(.A1(new_n291_), .A2(new_n886_), .ZN(new_n887_));
  OAI21_X1  g686(.A(KEYINPUT55), .B1(new_n281_), .B2(new_n202_), .ZN(new_n888_));
  AND2_X1   g687(.A1(new_n888_), .A2(new_n285_), .ZN(new_n889_));
  NOR2_X1   g688(.A1(new_n888_), .A2(new_n285_), .ZN(new_n890_));
  NOR3_X1   g689(.A1(new_n889_), .A2(new_n890_), .A3(new_n274_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n891_), .A2(KEYINPUT56), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n892_), .A2(KEYINPUT120), .ZN(new_n893_));
  NAND2_X1  g692(.A1(new_n892_), .A2(KEYINPUT120), .ZN(new_n894_));
  OR2_X1    g693(.A1(new_n891_), .A2(KEYINPUT56), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n893_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  NOR2_X1   g695(.A1(new_n283_), .A2(new_n286_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n823_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n887_), .B1(new_n896_), .B2(new_n898_), .ZN(new_n899_));
  INV_X1    g698(.A(new_n708_), .ZN(new_n900_));
  NOR2_X1   g699(.A1(new_n899_), .A2(new_n900_), .ZN(new_n901_));
  NAND2_X1  g700(.A1(new_n895_), .A2(new_n892_), .ZN(new_n902_));
  NOR2_X1   g701(.A1(new_n897_), .A2(new_n886_), .ZN(new_n903_));
  NAND3_X1  g702(.A1(new_n902_), .A2(KEYINPUT58), .A3(new_n903_), .ZN(new_n904_));
  AOI21_X1  g703(.A(KEYINPUT58), .B1(new_n902_), .B2(new_n903_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n691_), .ZN(new_n906_));
  AOI22_X1  g705(.A1(new_n901_), .A2(KEYINPUT57), .B1(new_n904_), .B2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(KEYINPUT57), .ZN(new_n908_));
  OAI21_X1  g707(.A(new_n908_), .B1(new_n899_), .B2(new_n900_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n909_), .A2(KEYINPUT122), .ZN(new_n910_));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911_));
  OAI211_X1 g710(.A(new_n911_), .B(new_n908_), .C1(new_n899_), .C2(new_n900_), .ZN(new_n912_));
  NAND3_X1  g711(.A1(new_n907_), .A2(new_n910_), .A3(new_n912_), .ZN(new_n913_));
  NAND2_X1  g712(.A1(new_n913_), .A2(new_n825_), .ZN(new_n914_));
  OR3_X1    g713(.A1(new_n825_), .A2(KEYINPUT119), .A3(new_n658_), .ZN(new_n915_));
  OAI21_X1  g714(.A(KEYINPUT119), .B1(new_n825_), .B2(new_n658_), .ZN(new_n916_));
  NAND4_X1  g715(.A1(new_n915_), .A2(new_n294_), .A3(new_n691_), .A4(new_n916_), .ZN(new_n917_));
  XOR2_X1   g716(.A(new_n917_), .B(KEYINPUT54), .Z(new_n918_));
  INV_X1    g717(.A(new_n918_), .ZN(new_n919_));
  AOI21_X1  g718(.A(new_n880_), .B1(new_n914_), .B2(new_n919_), .ZN(new_n920_));
  AOI21_X1  g719(.A(G113gat), .B1(new_n920_), .B2(new_n658_), .ZN(new_n921_));
  NAND2_X1  g720(.A1(new_n914_), .A2(new_n919_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n922_), .A2(new_n879_), .ZN(new_n923_));
  AND2_X1   g722(.A1(new_n907_), .A2(new_n909_), .ZN(new_n924_));
  OAI21_X1  g723(.A(new_n919_), .B1(new_n924_), .B2(new_n632_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n880_), .A2(KEYINPUT59), .ZN(new_n926_));
  AOI22_X1  g725(.A1(new_n923_), .A2(KEYINPUT59), .B1(new_n925_), .B2(new_n926_), .ZN(new_n927_));
  NAND2_X1  g726(.A1(new_n658_), .A2(G113gat), .ZN(new_n928_));
  XOR2_X1   g727(.A(new_n928_), .B(KEYINPUT123), .Z(new_n929_));
  AOI21_X1  g728(.A(new_n921_), .B1(new_n927_), .B2(new_n929_), .ZN(G1340gat));
  NAND2_X1  g729(.A1(new_n925_), .A2(new_n926_), .ZN(new_n931_));
  INV_X1    g730(.A(KEYINPUT59), .ZN(new_n932_));
  OAI21_X1  g731(.A(new_n931_), .B1(new_n920_), .B2(new_n932_), .ZN(new_n933_));
  OAI21_X1  g732(.A(G120gat), .B1(new_n933_), .B2(new_n297_), .ZN(new_n934_));
  NOR2_X1   g733(.A1(new_n461_), .A2(KEYINPUT60), .ZN(new_n935_));
  OAI21_X1  g734(.A(new_n461_), .B1(new_n294_), .B2(KEYINPUT60), .ZN(new_n936_));
  INV_X1    g735(.A(KEYINPUT124), .ZN(new_n937_));
  AOI21_X1  g736(.A(new_n935_), .B1(new_n936_), .B2(new_n937_), .ZN(new_n938_));
  OAI211_X1 g737(.A(new_n920_), .B(new_n938_), .C1(new_n937_), .C2(new_n936_), .ZN(new_n939_));
  NAND2_X1  g738(.A1(new_n934_), .A2(new_n939_), .ZN(G1341gat));
  AOI21_X1  g739(.A(G127gat), .B1(new_n920_), .B2(new_n632_), .ZN(new_n941_));
  AOI21_X1  g740(.A(new_n459_), .B1(new_n632_), .B2(KEYINPUT125), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n942_), .B1(KEYINPUT125), .B2(new_n459_), .ZN(new_n943_));
  AOI21_X1  g742(.A(new_n941_), .B1(new_n927_), .B2(new_n943_), .ZN(G1342gat));
  AOI211_X1 g743(.A(new_n708_), .B(new_n880_), .C1(new_n914_), .C2(new_n919_), .ZN(new_n945_));
  OAI21_X1  g744(.A(KEYINPUT126), .B1(new_n945_), .B2(G134gat), .ZN(new_n946_));
  INV_X1    g745(.A(KEYINPUT126), .ZN(new_n947_));
  OAI211_X1 g746(.A(new_n947_), .B(new_n457_), .C1(new_n923_), .C2(new_n708_), .ZN(new_n948_));
  NOR2_X1   g747(.A1(new_n691_), .A2(new_n457_), .ZN(new_n949_));
  AOI22_X1  g748(.A1(new_n946_), .A2(new_n948_), .B1(new_n927_), .B2(new_n949_), .ZN(G1343gat));
  NOR3_X1   g749(.A1(new_n718_), .A2(new_n704_), .A3(new_n565_), .ZN(new_n951_));
  NAND2_X1  g750(.A1(new_n922_), .A2(new_n951_), .ZN(new_n952_));
  INV_X1    g751(.A(new_n952_), .ZN(new_n953_));
  NAND3_X1  g752(.A1(new_n953_), .A2(new_n470_), .A3(new_n658_), .ZN(new_n954_));
  OAI21_X1  g753(.A(G141gat), .B1(new_n952_), .B2(new_n823_), .ZN(new_n955_));
  NAND2_X1  g754(.A1(new_n954_), .A2(new_n955_), .ZN(G1344gat));
  NAND3_X1  g755(.A1(new_n953_), .A2(new_n471_), .A3(new_n298_), .ZN(new_n957_));
  OAI21_X1  g756(.A(G148gat), .B1(new_n952_), .B2(new_n297_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n957_), .A2(new_n958_), .ZN(G1345gat));
  XNOR2_X1  g758(.A(KEYINPUT61), .B(G155gat), .ZN(new_n960_));
  OR3_X1    g759(.A1(new_n952_), .A2(new_n825_), .A3(new_n960_), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n960_), .B1(new_n952_), .B2(new_n825_), .ZN(new_n962_));
  NAND2_X1  g761(.A1(new_n961_), .A2(new_n962_), .ZN(G1346gat));
  OR3_X1    g762(.A1(new_n952_), .A2(G162gat), .A3(new_n708_), .ZN(new_n964_));
  OAI21_X1  g763(.A(G162gat), .B1(new_n952_), .B2(new_n691_), .ZN(new_n965_));
  NAND2_X1  g764(.A1(new_n964_), .A2(new_n965_), .ZN(G1347gat));
  NOR2_X1   g765(.A1(new_n439_), .A2(new_n514_), .ZN(new_n967_));
  NAND2_X1  g766(.A1(new_n967_), .A2(new_n600_), .ZN(new_n968_));
  NOR2_X1   g767(.A1(new_n968_), .A2(new_n601_), .ZN(new_n969_));
  NAND2_X1  g768(.A1(new_n925_), .A2(new_n969_), .ZN(new_n970_));
  OAI21_X1  g769(.A(G169gat), .B1(new_n970_), .B2(new_n823_), .ZN(new_n971_));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n972_));
  NAND2_X1  g771(.A1(new_n971_), .A2(new_n972_), .ZN(new_n973_));
  OAI211_X1 g772(.A(KEYINPUT62), .B(G169gat), .C1(new_n970_), .C2(new_n823_), .ZN(new_n974_));
  AND2_X1   g773(.A1(new_n925_), .A2(new_n969_), .ZN(new_n975_));
  NAND3_X1  g774(.A1(new_n975_), .A2(new_n364_), .A3(new_n658_), .ZN(new_n976_));
  NAND3_X1  g775(.A1(new_n973_), .A2(new_n974_), .A3(new_n976_), .ZN(G1348gat));
  AOI21_X1  g776(.A(G176gat), .B1(new_n975_), .B2(new_n711_), .ZN(new_n978_));
  AOI21_X1  g777(.A(new_n601_), .B1(new_n914_), .B2(new_n919_), .ZN(new_n979_));
  NOR3_X1   g778(.A1(new_n297_), .A2(new_n341_), .A3(new_n968_), .ZN(new_n980_));
  NAND2_X1  g779(.A1(new_n979_), .A2(new_n980_), .ZN(new_n981_));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n982_));
  NAND2_X1  g781(.A1(new_n981_), .A2(new_n982_), .ZN(new_n983_));
  NAND3_X1  g782(.A1(new_n979_), .A2(KEYINPUT127), .A3(new_n980_), .ZN(new_n984_));
  AOI21_X1  g783(.A(new_n978_), .B1(new_n983_), .B2(new_n984_), .ZN(G1349gat));
  NOR3_X1   g784(.A1(new_n970_), .A2(new_n356_), .A3(new_n825_), .ZN(new_n986_));
  NAND4_X1  g785(.A1(new_n979_), .A2(new_n600_), .A3(new_n632_), .A4(new_n967_), .ZN(new_n987_));
  AOI21_X1  g786(.A(new_n986_), .B1(new_n987_), .B2(new_n334_), .ZN(G1350gat));
  OAI21_X1  g787(.A(G190gat), .B1(new_n970_), .B2(new_n691_), .ZN(new_n989_));
  OAI21_X1  g788(.A(new_n900_), .B1(new_n359_), .B2(new_n360_), .ZN(new_n990_));
  OAI21_X1  g789(.A(new_n989_), .B1(new_n970_), .B2(new_n990_), .ZN(G1351gat));
  NAND3_X1  g790(.A1(new_n967_), .A2(new_n725_), .A3(new_n601_), .ZN(new_n992_));
  AOI21_X1  g791(.A(new_n992_), .B1(new_n914_), .B2(new_n919_), .ZN(new_n993_));
  NAND2_X1  g792(.A1(new_n993_), .A2(new_n658_), .ZN(new_n994_));
  XNOR2_X1  g793(.A(new_n994_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g794(.A1(new_n993_), .A2(new_n298_), .ZN(new_n996_));
  NOR2_X1   g795(.A1(new_n996_), .A2(new_n312_), .ZN(new_n997_));
  AOI21_X1  g796(.A(new_n997_), .B1(new_n271_), .B2(new_n996_), .ZN(G1353gat));
  NAND2_X1  g797(.A1(new_n993_), .A2(new_n632_), .ZN(new_n999_));
  XNOR2_X1  g798(.A(KEYINPUT63), .B(G211gat), .ZN(new_n1000_));
  NOR2_X1   g799(.A1(new_n999_), .A2(new_n1000_), .ZN(new_n1001_));
  NOR2_X1   g800(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n1002_));
  AOI21_X1  g801(.A(new_n1001_), .B1(new_n999_), .B2(new_n1002_), .ZN(G1354gat));
  INV_X1    g802(.A(G218gat), .ZN(new_n1004_));
  NAND3_X1  g803(.A1(new_n993_), .A2(new_n1004_), .A3(new_n900_), .ZN(new_n1005_));
  AND2_X1   g804(.A1(new_n993_), .A2(new_n692_), .ZN(new_n1006_));
  OAI21_X1  g805(.A(new_n1005_), .B1(new_n1006_), .B2(new_n1004_), .ZN(G1355gat));
endmodule


