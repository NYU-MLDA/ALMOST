//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1 1 0 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:31:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n585_, new_n586_, new_n587_,
    new_n588_, new_n590_, new_n591_, new_n592_, new_n593_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n644_, new_n645_, new_n646_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n657_, new_n658_, new_n659_, new_n660_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n684_, new_n685_, new_n686_, new_n687_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n806_, new_n807_,
    new_n809_, new_n810_, new_n812_, new_n813_, new_n814_, new_n815_,
    new_n816_, new_n818_, new_n820_, new_n821_, new_n822_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n845_, new_n846_, new_n847_, new_n849_, new_n851_, new_n852_,
    new_n853_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n862_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_;
  INV_X1    g000(.A(G1gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G127gat), .B(G134gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(G113gat), .ZN(new_n204_));
  INV_X1    g003(.A(G120gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  NOR2_X1   g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  NAND2_X1  g007(.A1(G141gat), .A2(G148gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(G155gat), .A2(G162gat), .ZN(new_n210_));
  XNOR2_X1  g009(.A(new_n210_), .B(KEYINPUT84), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212_));
  XNOR2_X1  g011(.A(new_n212_), .B(KEYINPUT1), .ZN(new_n213_));
  OAI211_X1 g012(.A(new_n208_), .B(new_n209_), .C1(new_n211_), .C2(new_n213_), .ZN(new_n214_));
  XOR2_X1   g013(.A(new_n207_), .B(KEYINPUT3), .Z(new_n215_));
  XOR2_X1   g014(.A(new_n209_), .B(KEYINPUT2), .Z(new_n216_));
  OAI21_X1  g015(.A(new_n212_), .B1(new_n215_), .B2(new_n216_), .ZN(new_n217_));
  OAI21_X1  g016(.A(new_n214_), .B1(new_n217_), .B2(new_n211_), .ZN(new_n218_));
  XOR2_X1   g017(.A(new_n206_), .B(new_n218_), .Z(new_n219_));
  NAND2_X1  g018(.A1(new_n219_), .A2(KEYINPUT4), .ZN(new_n220_));
  NAND2_X1  g019(.A1(new_n206_), .A2(new_n218_), .ZN(new_n221_));
  OAI21_X1  g020(.A(new_n220_), .B1(KEYINPUT4), .B2(new_n221_), .ZN(new_n222_));
  NAND2_X1  g021(.A1(G225gat), .A2(G233gat), .ZN(new_n223_));
  OR2_X1    g022(.A1(new_n222_), .A2(new_n223_), .ZN(new_n224_));
  NAND2_X1  g023(.A1(new_n219_), .A2(new_n223_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n224_), .A2(new_n225_), .ZN(new_n226_));
  XNOR2_X1  g025(.A(KEYINPUT0), .B(G57gat), .ZN(new_n227_));
  XNOR2_X1  g026(.A(new_n227_), .B(G85gat), .ZN(new_n228_));
  XOR2_X1   g027(.A(G1gat), .B(G29gat), .Z(new_n229_));
  XOR2_X1   g028(.A(new_n228_), .B(new_n229_), .Z(new_n230_));
  NAND2_X1  g029(.A1(new_n226_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(new_n230_), .ZN(new_n232_));
  NAND3_X1  g031(.A1(new_n224_), .A2(new_n225_), .A3(new_n232_), .ZN(new_n233_));
  NAND2_X1  g032(.A1(new_n231_), .A2(new_n233_), .ZN(new_n234_));
  INV_X1    g033(.A(KEYINPUT94), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n234_), .A2(new_n235_), .ZN(new_n236_));
  NAND3_X1  g035(.A1(new_n231_), .A2(KEYINPUT94), .A3(new_n233_), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(new_n238_), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT12), .ZN(new_n240_));
  XOR2_X1   g039(.A(KEYINPUT10), .B(G99gat), .Z(new_n241_));
  INV_X1    g040(.A(G106gat), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  XOR2_X1   g042(.A(G85gat), .B(G92gat), .Z(new_n244_));
  NAND2_X1  g043(.A1(new_n244_), .A2(KEYINPUT9), .ZN(new_n245_));
  INV_X1    g044(.A(KEYINPUT9), .ZN(new_n246_));
  NAND3_X1  g045(.A1(new_n246_), .A2(G85gat), .A3(G92gat), .ZN(new_n247_));
  NAND2_X1  g046(.A1(G99gat), .A2(G106gat), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT6), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(new_n252_), .ZN(new_n253_));
  NAND4_X1  g052(.A1(new_n243_), .A2(new_n245_), .A3(new_n247_), .A4(new_n253_), .ZN(new_n254_));
  INV_X1    g053(.A(new_n254_), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT65), .ZN(new_n256_));
  AND3_X1   g055(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n257_));
  AOI21_X1  g056(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n256_), .B1(new_n257_), .B2(new_n258_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n250_), .A2(KEYINPUT65), .A3(new_n251_), .ZN(new_n260_));
  AND2_X1   g059(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n261_));
  NOR2_X1   g060(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n262_));
  OAI22_X1  g061(.A1(new_n261_), .A2(new_n262_), .B1(G99gat), .B2(G106gat), .ZN(new_n263_));
  NAND2_X1  g062(.A1(KEYINPUT64), .A2(KEYINPUT7), .ZN(new_n264_));
  INV_X1    g063(.A(G99gat), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n264_), .A2(new_n265_), .A3(new_n242_), .ZN(new_n266_));
  NAND4_X1  g065(.A1(new_n259_), .A2(new_n260_), .A3(new_n263_), .A4(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n267_), .A2(new_n244_), .ZN(new_n268_));
  AOI21_X1  g067(.A(KEYINPUT66), .B1(new_n268_), .B2(KEYINPUT8), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT66), .ZN(new_n270_));
  INV_X1    g069(.A(KEYINPUT8), .ZN(new_n271_));
  AOI211_X1 g070(.A(new_n270_), .B(new_n271_), .C1(new_n267_), .C2(new_n244_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n269_), .A2(new_n272_), .ZN(new_n273_));
  NAND3_X1  g072(.A1(new_n253_), .A2(new_n263_), .A3(new_n266_), .ZN(new_n274_));
  NAND3_X1  g073(.A1(new_n274_), .A2(new_n271_), .A3(new_n244_), .ZN(new_n275_));
  AOI21_X1  g074(.A(new_n255_), .B1(new_n273_), .B2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(KEYINPUT67), .B(G78gat), .ZN(new_n277_));
  OR2_X1    g076(.A1(new_n277_), .A2(G71gat), .ZN(new_n278_));
  XOR2_X1   g077(.A(G57gat), .B(G64gat), .Z(new_n279_));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n280_));
  NAND2_X1  g079(.A1(new_n279_), .A2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n277_), .A2(G71gat), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n278_), .A2(new_n281_), .A3(new_n282_), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n283_), .A2(KEYINPUT68), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n285_));
  NAND4_X1  g084(.A1(new_n281_), .A2(new_n278_), .A3(new_n285_), .A4(new_n282_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n279_), .A2(new_n280_), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n284_), .A2(new_n286_), .A3(new_n287_), .ZN(new_n288_));
  INV_X1    g087(.A(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n287_), .B1(new_n284_), .B2(new_n286_), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n289_), .A2(new_n290_), .ZN(new_n291_));
  OAI21_X1  g090(.A(new_n240_), .B1(new_n276_), .B2(new_n291_), .ZN(new_n292_));
  AND2_X1   g091(.A1(G230gat), .A2(G233gat), .ZN(new_n293_));
  AOI21_X1  g092(.A(new_n293_), .B1(new_n276_), .B2(new_n291_), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n268_), .A2(KEYINPUT8), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n295_), .A2(new_n270_), .ZN(new_n296_));
  NAND3_X1  g095(.A1(new_n268_), .A2(KEYINPUT66), .A3(KEYINPUT8), .ZN(new_n297_));
  NAND3_X1  g096(.A1(new_n296_), .A2(new_n297_), .A3(new_n275_), .ZN(new_n298_));
  NAND2_X1  g097(.A1(new_n298_), .A2(new_n254_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n290_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n288_), .ZN(new_n301_));
  NAND3_X1  g100(.A1(new_n299_), .A2(new_n301_), .A3(KEYINPUT12), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n292_), .A2(new_n294_), .A3(new_n302_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n304_));
  NAND2_X1  g103(.A1(new_n303_), .A2(new_n304_), .ZN(new_n305_));
  NAND4_X1  g104(.A1(new_n292_), .A2(new_n294_), .A3(KEYINPUT69), .A4(new_n302_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n276_), .A2(new_n291_), .ZN(new_n308_));
  INV_X1    g107(.A(new_n308_), .ZN(new_n309_));
  NOR2_X1   g108(.A1(new_n276_), .A2(new_n291_), .ZN(new_n310_));
  OAI21_X1  g109(.A(new_n293_), .B1(new_n309_), .B2(new_n310_), .ZN(new_n311_));
  AND2_X1   g110(.A1(new_n307_), .A2(new_n311_), .ZN(new_n312_));
  XOR2_X1   g111(.A(G120gat), .B(G148gat), .Z(new_n313_));
  XNOR2_X1  g112(.A(new_n313_), .B(G204gat), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT5), .ZN(new_n315_));
  INV_X1    g114(.A(G176gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(new_n315_), .B(new_n316_), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n312_), .A2(new_n317_), .ZN(new_n318_));
  XNOR2_X1  g117(.A(new_n317_), .B(KEYINPUT70), .ZN(new_n319_));
  OAI21_X1  g118(.A(new_n318_), .B1(new_n312_), .B2(new_n319_), .ZN(new_n320_));
  INV_X1    g119(.A(KEYINPUT13), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n320_), .A2(new_n321_), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n320_), .A2(new_n321_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  XNOR2_X1  g123(.A(G29gat), .B(G36gat), .ZN(new_n325_));
  XNOR2_X1  g124(.A(G43gat), .B(G50gat), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n325_), .B(new_n326_), .ZN(new_n327_));
  XNOR2_X1  g126(.A(KEYINPUT72), .B(KEYINPUT73), .ZN(new_n328_));
  INV_X1    g127(.A(new_n328_), .ZN(new_n329_));
  OR2_X1    g128(.A1(new_n327_), .A2(new_n329_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n327_), .A2(new_n329_), .ZN(new_n331_));
  NAND2_X1  g130(.A1(new_n330_), .A2(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(new_n332_), .ZN(new_n333_));
  NAND2_X1  g132(.A1(new_n333_), .A2(KEYINPUT15), .ZN(new_n334_));
  INV_X1    g133(.A(KEYINPUT15), .ZN(new_n335_));
  NAND2_X1  g134(.A1(new_n332_), .A2(new_n335_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n334_), .A2(new_n336_), .ZN(new_n337_));
  INV_X1    g136(.A(new_n337_), .ZN(new_n338_));
  XOR2_X1   g137(.A(G15gat), .B(G22gat), .Z(new_n339_));
  NAND2_X1  g138(.A1(G1gat), .A2(G8gat), .ZN(new_n340_));
  AOI21_X1  g139(.A(new_n339_), .B1(KEYINPUT14), .B2(new_n340_), .ZN(new_n341_));
  XNOR2_X1  g140(.A(new_n341_), .B(KEYINPUT76), .ZN(new_n342_));
  XOR2_X1   g141(.A(G1gat), .B(G8gat), .Z(new_n343_));
  NAND2_X1  g142(.A1(new_n342_), .A2(new_n343_), .ZN(new_n344_));
  INV_X1    g143(.A(KEYINPUT76), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n341_), .B(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n343_), .ZN(new_n347_));
  NAND2_X1  g146(.A1(new_n346_), .A2(new_n347_), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n344_), .A2(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n338_), .A2(new_n350_), .ZN(new_n351_));
  AOI21_X1  g150(.A(new_n333_), .B1(new_n344_), .B2(new_n348_), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n354_));
  NAND2_X1  g153(.A1(G229gat), .A2(G233gat), .ZN(new_n355_));
  NAND4_X1  g154(.A1(new_n351_), .A2(new_n353_), .A3(new_n354_), .A4(new_n355_), .ZN(new_n356_));
  NOR2_X1   g155(.A1(new_n349_), .A2(new_n332_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n357_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n358_), .A2(new_n353_), .A3(KEYINPUT77), .ZN(new_n359_));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n360_));
  OAI21_X1  g159(.A(new_n360_), .B1(new_n357_), .B2(new_n352_), .ZN(new_n361_));
  INV_X1    g160(.A(new_n355_), .ZN(new_n362_));
  NAND3_X1  g161(.A1(new_n359_), .A2(new_n361_), .A3(new_n362_), .ZN(new_n363_));
  OAI211_X1 g162(.A(new_n353_), .B(new_n355_), .C1(new_n349_), .C2(new_n337_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n364_), .A2(KEYINPUT78), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n356_), .A2(new_n363_), .A3(new_n365_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(G113gat), .B(G141gat), .ZN(new_n367_));
  INV_X1    g166(.A(G169gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(new_n367_), .B(new_n368_), .ZN(new_n369_));
  INV_X1    g168(.A(G197gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  NAND2_X1  g170(.A1(new_n366_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(new_n371_), .ZN(new_n373_));
  NAND4_X1  g172(.A1(new_n356_), .A2(new_n363_), .A3(new_n365_), .A4(new_n373_), .ZN(new_n374_));
  NAND2_X1  g173(.A1(new_n372_), .A2(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NOR2_X1   g175(.A1(new_n324_), .A2(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  NAND2_X1  g177(.A1(G183gat), .A2(G190gat), .ZN(new_n379_));
  XNOR2_X1  g178(.A(new_n379_), .B(KEYINPUT23), .ZN(new_n380_));
  OAI21_X1  g179(.A(new_n380_), .B1(G183gat), .B2(G190gat), .ZN(new_n381_));
  NAND2_X1  g180(.A1(G169gat), .A2(G176gat), .ZN(new_n382_));
  AND2_X1   g181(.A1(new_n381_), .A2(new_n382_), .ZN(new_n383_));
  NAND2_X1  g182(.A1(new_n368_), .A2(KEYINPUT22), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n384_), .A2(KEYINPUT81), .ZN(new_n385_));
  OR2_X1    g184(.A1(new_n368_), .A2(KEYINPUT22), .ZN(new_n386_));
  NAND2_X1  g185(.A1(new_n384_), .A2(KEYINPUT81), .ZN(new_n387_));
  NAND4_X1  g186(.A1(new_n385_), .A2(new_n316_), .A3(new_n386_), .A4(new_n387_), .ZN(new_n388_));
  NAND2_X1  g187(.A1(new_n383_), .A2(new_n388_), .ZN(new_n389_));
  NOR2_X1   g188(.A1(G169gat), .A2(G176gat), .ZN(new_n390_));
  INV_X1    g189(.A(new_n390_), .ZN(new_n391_));
  AND3_X1   g190(.A1(new_n391_), .A2(KEYINPUT24), .A3(new_n382_), .ZN(new_n392_));
  INV_X1    g191(.A(new_n392_), .ZN(new_n393_));
  XNOR2_X1  g192(.A(KEYINPUT79), .B(KEYINPUT26), .ZN(new_n394_));
  INV_X1    g193(.A(KEYINPUT80), .ZN(new_n395_));
  AND2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  OR2_X1    g195(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n397_));
  INV_X1    g196(.A(G190gat), .ZN(new_n398_));
  OAI21_X1  g197(.A(new_n397_), .B1(new_n394_), .B2(new_n398_), .ZN(new_n399_));
  AOI22_X1  g198(.A1(G190gat), .A2(new_n396_), .B1(new_n399_), .B2(KEYINPUT80), .ZN(new_n400_));
  XNOR2_X1  g199(.A(KEYINPUT25), .B(G183gat), .ZN(new_n401_));
  INV_X1    g200(.A(new_n401_), .ZN(new_n402_));
  OAI21_X1  g201(.A(new_n393_), .B1(new_n400_), .B2(new_n402_), .ZN(new_n403_));
  OR2_X1    g202(.A1(new_n391_), .A2(KEYINPUT24), .ZN(new_n404_));
  NAND2_X1  g203(.A1(new_n404_), .A2(new_n380_), .ZN(new_n405_));
  OAI21_X1  g204(.A(new_n389_), .B1(new_n403_), .B2(new_n405_), .ZN(new_n406_));
  XNOR2_X1  g205(.A(G211gat), .B(G218gat), .ZN(new_n407_));
  XOR2_X1   g206(.A(G197gat), .B(G204gat), .Z(new_n408_));
  OAI21_X1  g207(.A(new_n407_), .B1(new_n408_), .B2(KEYINPUT21), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n408_), .A2(KEYINPUT21), .ZN(new_n410_));
  XNOR2_X1  g209(.A(new_n409_), .B(new_n410_), .ZN(new_n411_));
  INV_X1    g210(.A(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n406_), .A2(new_n412_), .ZN(new_n413_));
  NAND3_X1  g212(.A1(new_n386_), .A2(new_n384_), .A3(new_n316_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n383_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(KEYINPUT88), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n405_), .A2(new_n416_), .ZN(new_n417_));
  XNOR2_X1  g216(.A(KEYINPUT26), .B(G190gat), .ZN(new_n418_));
  AOI21_X1  g217(.A(new_n392_), .B1(new_n401_), .B2(new_n418_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n380_), .A2(KEYINPUT88), .A3(new_n404_), .ZN(new_n420_));
  NAND3_X1  g219(.A1(new_n417_), .A2(new_n419_), .A3(new_n420_), .ZN(new_n421_));
  NAND3_X1  g220(.A1(new_n415_), .A2(new_n411_), .A3(new_n421_), .ZN(new_n422_));
  AND3_X1   g221(.A1(new_n413_), .A2(KEYINPUT20), .A3(new_n422_), .ZN(new_n423_));
  NAND2_X1  g222(.A1(G226gat), .A2(G233gat), .ZN(new_n424_));
  XOR2_X1   g223(.A(new_n424_), .B(KEYINPUT19), .Z(new_n425_));
  NAND2_X1  g224(.A1(new_n423_), .A2(new_n425_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n415_), .A2(new_n421_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n427_), .A2(new_n412_), .ZN(new_n428_));
  OAI211_X1 g227(.A(new_n428_), .B(KEYINPUT20), .C1(new_n406_), .C2(new_n412_), .ZN(new_n429_));
  XNOR2_X1  g228(.A(new_n425_), .B(KEYINPUT87), .ZN(new_n430_));
  NAND2_X1  g229(.A1(new_n429_), .A2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n426_), .A2(new_n431_), .ZN(new_n432_));
  XOR2_X1   g231(.A(G8gat), .B(G36gat), .Z(new_n433_));
  XNOR2_X1  g232(.A(G64gat), .B(G92gat), .ZN(new_n434_));
  XNOR2_X1  g233(.A(new_n433_), .B(new_n434_), .ZN(new_n435_));
  XNOR2_X1  g234(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n436_));
  XOR2_X1   g235(.A(new_n435_), .B(new_n436_), .Z(new_n437_));
  NAND2_X1  g236(.A1(new_n432_), .A2(new_n437_), .ZN(new_n438_));
  INV_X1    g237(.A(new_n437_), .ZN(new_n439_));
  NAND3_X1  g238(.A1(new_n426_), .A2(new_n431_), .A3(new_n439_), .ZN(new_n440_));
  NAND3_X1  g239(.A1(new_n438_), .A2(KEYINPUT90), .A3(new_n440_), .ZN(new_n441_));
  INV_X1    g240(.A(new_n441_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n432_), .ZN(new_n443_));
  NOR3_X1   g242(.A1(new_n443_), .A2(KEYINPUT90), .A3(new_n439_), .ZN(new_n444_));
  OR3_X1    g243(.A1(new_n442_), .A2(KEYINPUT27), .A3(new_n444_), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n423_), .A2(new_n425_), .ZN(new_n446_));
  NOR2_X1   g245(.A1(new_n429_), .A2(new_n430_), .ZN(new_n447_));
  NOR2_X1   g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  OAI211_X1 g247(.A(KEYINPUT27), .B(new_n440_), .C1(new_n448_), .C2(new_n439_), .ZN(new_n449_));
  AOI21_X1  g248(.A(new_n411_), .B1(new_n218_), .B2(KEYINPUT29), .ZN(new_n450_));
  XOR2_X1   g249(.A(KEYINPUT85), .B(G233gat), .Z(new_n451_));
  AND2_X1   g250(.A1(new_n451_), .A2(G228gat), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n450_), .A2(KEYINPUT86), .A3(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(new_n452_), .B(KEYINPUT86), .ZN(new_n454_));
  OAI21_X1  g253(.A(new_n453_), .B1(new_n450_), .B2(new_n454_), .ZN(new_n455_));
  XNOR2_X1  g254(.A(G22gat), .B(G50gat), .ZN(new_n456_));
  XNOR2_X1  g255(.A(new_n456_), .B(G78gat), .ZN(new_n457_));
  XNOR2_X1  g256(.A(new_n455_), .B(new_n457_), .ZN(new_n458_));
  NOR2_X1   g257(.A1(new_n218_), .A2(KEYINPUT29), .ZN(new_n459_));
  XNOR2_X1  g258(.A(new_n459_), .B(KEYINPUT28), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n460_), .B(new_n242_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n458_), .A2(new_n461_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n458_), .A2(new_n461_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(G15gat), .B(G43gat), .ZN(new_n465_));
  NAND2_X1  g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n465_), .B(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n206_), .B(new_n467_), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(new_n406_), .ZN(new_n469_));
  XNOR2_X1  g268(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n470_));
  XNOR2_X1  g269(.A(KEYINPUT82), .B(KEYINPUT30), .ZN(new_n471_));
  XNOR2_X1  g270(.A(new_n470_), .B(new_n471_), .ZN(new_n472_));
  XNOR2_X1  g271(.A(G71gat), .B(G99gat), .ZN(new_n473_));
  XNOR2_X1  g272(.A(new_n472_), .B(new_n473_), .ZN(new_n474_));
  XOR2_X1   g273(.A(new_n469_), .B(new_n474_), .Z(new_n475_));
  NOR2_X1   g274(.A1(new_n464_), .A2(new_n475_), .ZN(new_n476_));
  NAND4_X1  g275(.A1(new_n238_), .A2(new_n445_), .A3(new_n449_), .A4(new_n476_), .ZN(new_n477_));
  XNOR2_X1  g276(.A(new_n477_), .B(KEYINPUT95), .ZN(new_n478_));
  INV_X1    g277(.A(KEYINPUT91), .ZN(new_n479_));
  OAI21_X1  g278(.A(new_n479_), .B1(new_n442_), .B2(new_n444_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n444_), .ZN(new_n481_));
  NAND3_X1  g280(.A1(new_n481_), .A2(KEYINPUT91), .A3(new_n441_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n480_), .A2(new_n482_), .ZN(new_n483_));
  NOR2_X1   g282(.A1(KEYINPUT92), .A2(KEYINPUT33), .ZN(new_n484_));
  OR2_X1    g283(.A1(new_n233_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n223_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n230_), .B1(new_n222_), .B2(new_n486_), .ZN(new_n487_));
  AOI21_X1  g286(.A(new_n487_), .B1(new_n486_), .B2(new_n219_), .ZN(new_n488_));
  XNOR2_X1  g287(.A(new_n488_), .B(KEYINPUT93), .ZN(new_n489_));
  AND2_X1   g288(.A1(KEYINPUT92), .A2(KEYINPUT33), .ZN(new_n490_));
  OAI21_X1  g289(.A(new_n233_), .B1(new_n484_), .B2(new_n490_), .ZN(new_n491_));
  NAND4_X1  g290(.A1(new_n483_), .A2(new_n485_), .A3(new_n489_), .A4(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n439_), .A2(KEYINPUT32), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n443_), .A2(new_n493_), .ZN(new_n494_));
  OAI211_X1 g293(.A(new_n234_), .B(new_n494_), .C1(new_n493_), .C2(new_n448_), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n464_), .B1(new_n492_), .B2(new_n495_), .ZN(new_n496_));
  AND4_X1   g295(.A1(new_n238_), .A2(new_n445_), .A3(new_n464_), .A4(new_n449_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n475_), .B1(new_n496_), .B2(new_n497_), .ZN(new_n498_));
  AOI21_X1  g297(.A(new_n378_), .B1(new_n478_), .B2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(G231gat), .A2(G233gat), .ZN(new_n500_));
  XNOR2_X1  g299(.A(new_n301_), .B(new_n500_), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(new_n350_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(KEYINPUT16), .B(G183gat), .ZN(new_n503_));
  INV_X1    g302(.A(G211gat), .ZN(new_n504_));
  XNOR2_X1  g303(.A(new_n503_), .B(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G127gat), .B(G155gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(new_n505_), .B(new_n506_), .ZN(new_n507_));
  INV_X1    g306(.A(KEYINPUT17), .ZN(new_n508_));
  NOR2_X1   g307(.A1(new_n507_), .A2(new_n508_), .ZN(new_n509_));
  AND2_X1   g308(.A1(new_n507_), .A2(new_n508_), .ZN(new_n510_));
  NOR3_X1   g309(.A1(new_n502_), .A2(new_n509_), .A3(new_n510_), .ZN(new_n511_));
  AOI21_X1  g310(.A(new_n511_), .B1(new_n509_), .B2(new_n502_), .ZN(new_n512_));
  INV_X1    g311(.A(new_n512_), .ZN(new_n513_));
  NOR2_X1   g312(.A1(new_n299_), .A2(new_n333_), .ZN(new_n514_));
  XNOR2_X1  g313(.A(new_n514_), .B(KEYINPUT74), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G232gat), .A2(G233gat), .ZN(new_n516_));
  XNOR2_X1  g315(.A(new_n516_), .B(KEYINPUT34), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n517_), .A2(KEYINPUT35), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n518_), .B1(new_n338_), .B2(new_n299_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n515_), .A2(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n517_), .A2(KEYINPUT35), .ZN(new_n521_));
  XOR2_X1   g320(.A(new_n521_), .B(KEYINPUT71), .Z(new_n522_));
  NAND2_X1  g321(.A1(new_n520_), .A2(new_n522_), .ZN(new_n523_));
  INV_X1    g322(.A(KEYINPUT36), .ZN(new_n524_));
  XNOR2_X1  g323(.A(G190gat), .B(G218gat), .ZN(new_n525_));
  XNOR2_X1  g324(.A(new_n525_), .B(G134gat), .ZN(new_n526_));
  INV_X1    g325(.A(G162gat), .ZN(new_n527_));
  XNOR2_X1  g326(.A(new_n526_), .B(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n522_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n515_), .A2(new_n529_), .A3(new_n519_), .ZN(new_n530_));
  NAND4_X1  g329(.A1(new_n523_), .A2(new_n524_), .A3(new_n528_), .A4(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(new_n531_), .ZN(new_n532_));
  XNOR2_X1  g331(.A(new_n528_), .B(KEYINPUT36), .ZN(new_n533_));
  INV_X1    g332(.A(new_n533_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n534_), .B1(new_n523_), .B2(new_n530_), .ZN(new_n535_));
  NOR2_X1   g334(.A1(new_n532_), .A2(new_n535_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT75), .ZN(new_n537_));
  NAND2_X1  g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(KEYINPUT75), .B1(new_n532_), .B2(new_n535_), .ZN(new_n539_));
  NAND3_X1  g338(.A1(new_n538_), .A2(KEYINPUT37), .A3(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT37), .ZN(new_n541_));
  NOR3_X1   g340(.A1(new_n532_), .A2(KEYINPUT75), .A3(new_n535_), .ZN(new_n542_));
  INV_X1    g341(.A(new_n535_), .ZN(new_n543_));
  AOI21_X1  g342(.A(new_n537_), .B1(new_n543_), .B2(new_n531_), .ZN(new_n544_));
  OAI21_X1  g343(.A(new_n541_), .B1(new_n542_), .B2(new_n544_), .ZN(new_n545_));
  AOI21_X1  g344(.A(new_n513_), .B1(new_n540_), .B2(new_n545_), .ZN(new_n546_));
  AND3_X1   g345(.A1(new_n499_), .A2(KEYINPUT96), .A3(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(KEYINPUT96), .B1(new_n499_), .B2(new_n546_), .ZN(new_n548_));
  OAI211_X1 g347(.A(new_n202_), .B(new_n239_), .C1(new_n547_), .C2(new_n548_), .ZN(new_n549_));
  INV_X1    g348(.A(KEYINPUT38), .ZN(new_n550_));
  OR2_X1    g349(.A1(new_n549_), .A2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(new_n478_), .A2(new_n498_), .ZN(new_n552_));
  INV_X1    g351(.A(new_n536_), .ZN(new_n553_));
  NAND4_X1  g352(.A1(new_n552_), .A2(new_n512_), .A3(new_n377_), .A4(new_n553_), .ZN(new_n554_));
  OAI21_X1  g353(.A(G1gat), .B1(new_n554_), .B2(new_n238_), .ZN(new_n555_));
  NAND2_X1  g354(.A1(new_n549_), .A2(new_n550_), .ZN(new_n556_));
  NAND3_X1  g355(.A1(new_n551_), .A2(new_n555_), .A3(new_n556_), .ZN(G1324gat));
  INV_X1    g356(.A(G8gat), .ZN(new_n558_));
  AND2_X1   g357(.A1(new_n445_), .A2(new_n449_), .ZN(new_n559_));
  INV_X1    g358(.A(new_n559_), .ZN(new_n560_));
  OAI211_X1 g359(.A(new_n558_), .B(new_n560_), .C1(new_n547_), .C2(new_n548_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT97), .ZN(new_n562_));
  NAND3_X1  g361(.A1(new_n552_), .A2(new_n377_), .A3(new_n546_), .ZN(new_n563_));
  INV_X1    g362(.A(KEYINPUT96), .ZN(new_n564_));
  NAND2_X1  g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NAND3_X1  g364(.A1(new_n499_), .A2(KEYINPUT96), .A3(new_n546_), .ZN(new_n566_));
  AOI21_X1  g365(.A(G8gat), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(KEYINPUT97), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n567_), .A2(new_n568_), .A3(new_n560_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n562_), .A2(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT98), .ZN(new_n571_));
  OAI21_X1  g370(.A(G8gat), .B1(new_n554_), .B2(new_n559_), .ZN(new_n572_));
  XNOR2_X1  g371(.A(new_n572_), .B(KEYINPUT39), .ZN(new_n573_));
  AND3_X1   g372(.A1(new_n570_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n574_));
  AOI21_X1  g373(.A(new_n571_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT40), .ZN(new_n576_));
  NOR3_X1   g375(.A1(new_n574_), .A2(new_n575_), .A3(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n561_), .A2(KEYINPUT97), .ZN(new_n578_));
  AOI21_X1  g377(.A(new_n568_), .B1(new_n567_), .B2(new_n560_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n573_), .B1(new_n578_), .B2(new_n579_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT98), .ZN(new_n581_));
  NAND3_X1  g380(.A1(new_n570_), .A2(new_n571_), .A3(new_n573_), .ZN(new_n582_));
  AOI21_X1  g381(.A(KEYINPUT40), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n577_), .A2(new_n583_), .ZN(G1325gat));
  OAI21_X1  g383(.A(G15gat), .B1(new_n554_), .B2(new_n475_), .ZN(new_n585_));
  XOR2_X1   g384(.A(new_n585_), .B(KEYINPUT99), .Z(new_n586_));
  XNOR2_X1  g385(.A(new_n586_), .B(KEYINPUT41), .ZN(new_n587_));
  NOR3_X1   g386(.A1(new_n563_), .A2(G15gat), .A3(new_n475_), .ZN(new_n588_));
  OR2_X1    g387(.A1(new_n587_), .A2(new_n588_), .ZN(G1326gat));
  INV_X1    g388(.A(new_n464_), .ZN(new_n590_));
  OAI21_X1  g389(.A(G22gat), .B1(new_n554_), .B2(new_n590_), .ZN(new_n591_));
  XNOR2_X1  g390(.A(new_n591_), .B(KEYINPUT42), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n590_), .A2(G22gat), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n592_), .B1(new_n563_), .B2(new_n593_), .ZN(G1327gat));
  NAND2_X1  g393(.A1(new_n540_), .A2(new_n545_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n552_), .A2(new_n596_), .ZN(new_n597_));
  NAND3_X1  g396(.A1(new_n597_), .A2(KEYINPUT100), .A3(KEYINPUT43), .ZN(new_n598_));
  INV_X1    g397(.A(KEYINPUT43), .ZN(new_n599_));
  AOI21_X1  g398(.A(new_n595_), .B1(new_n478_), .B2(new_n498_), .ZN(new_n600_));
  INV_X1    g399(.A(KEYINPUT100), .ZN(new_n601_));
  OAI21_X1  g400(.A(new_n599_), .B1(new_n600_), .B2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n598_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(new_n513_), .A3(new_n377_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT44), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  AOI21_X1  g406(.A(new_n512_), .B1(new_n598_), .B2(new_n602_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n608_), .A2(KEYINPUT44), .A3(new_n377_), .ZN(new_n609_));
  NAND2_X1  g408(.A1(new_n609_), .A2(new_n239_), .ZN(new_n610_));
  OAI21_X1  g409(.A(G29gat), .B1(new_n607_), .B2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n553_), .A2(new_n512_), .ZN(new_n612_));
  AND2_X1   g411(.A1(new_n499_), .A2(new_n612_), .ZN(new_n613_));
  NOR2_X1   g412(.A1(new_n238_), .A2(G29gat), .ZN(new_n614_));
  XNOR2_X1  g413(.A(new_n614_), .B(KEYINPUT101), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n613_), .A2(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n611_), .A2(new_n616_), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT102), .ZN(new_n618_));
  NAND2_X1  g417(.A1(new_n617_), .A2(new_n618_), .ZN(new_n619_));
  NAND3_X1  g418(.A1(new_n611_), .A2(KEYINPUT102), .A3(new_n616_), .ZN(new_n620_));
  NAND2_X1  g419(.A1(new_n619_), .A2(new_n620_), .ZN(G1328gat));
  NAND3_X1  g420(.A1(new_n606_), .A2(new_n560_), .A3(new_n609_), .ZN(new_n622_));
  NAND2_X1  g421(.A1(new_n622_), .A2(G36gat), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT103), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT46), .ZN(new_n625_));
  INV_X1    g424(.A(G36gat), .ZN(new_n626_));
  NAND3_X1  g425(.A1(new_n613_), .A2(new_n626_), .A3(new_n560_), .ZN(new_n627_));
  XNOR2_X1  g426(.A(new_n627_), .B(KEYINPUT45), .ZN(new_n628_));
  NAND4_X1  g427(.A1(new_n623_), .A2(new_n624_), .A3(new_n625_), .A4(new_n628_), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n624_), .A2(new_n625_), .ZN(new_n630_));
  NAND2_X1  g429(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n631_));
  AOI21_X1  g430(.A(new_n559_), .B1(new_n604_), .B2(new_n605_), .ZN(new_n632_));
  AOI21_X1  g431(.A(new_n626_), .B1(new_n632_), .B2(new_n609_), .ZN(new_n633_));
  INV_X1    g432(.A(new_n628_), .ZN(new_n634_));
  OAI211_X1 g433(.A(new_n630_), .B(new_n631_), .C1(new_n633_), .C2(new_n634_), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n629_), .A2(new_n635_), .ZN(G1329gat));
  INV_X1    g435(.A(new_n475_), .ZN(new_n637_));
  AOI21_X1  g436(.A(G43gat), .B1(new_n613_), .B2(new_n637_), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n638_), .B(KEYINPUT104), .Z(new_n639_));
  NAND2_X1  g438(.A1(new_n606_), .A2(new_n637_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n609_), .A2(G43gat), .ZN(new_n641_));
  OAI21_X1  g440(.A(new_n639_), .B1(new_n640_), .B2(new_n641_), .ZN(new_n642_));
  XNOR2_X1  g441(.A(new_n642_), .B(KEYINPUT47), .ZN(G1330gat));
  AOI21_X1  g442(.A(G50gat), .B1(new_n613_), .B2(new_n464_), .ZN(new_n644_));
  NOR2_X1   g443(.A1(new_n607_), .A2(new_n590_), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n609_), .A2(G50gat), .ZN(new_n646_));
  AOI21_X1  g445(.A(new_n644_), .B1(new_n645_), .B2(new_n646_), .ZN(G1331gat));
  INV_X1    g446(.A(new_n324_), .ZN(new_n648_));
  NOR2_X1   g447(.A1(new_n648_), .A2(new_n375_), .ZN(new_n649_));
  AND2_X1   g448(.A1(new_n552_), .A2(new_n649_), .ZN(new_n650_));
  AND2_X1   g449(.A1(new_n650_), .A2(new_n546_), .ZN(new_n651_));
  AOI21_X1  g450(.A(G57gat), .B1(new_n651_), .B2(new_n239_), .ZN(new_n652_));
  NAND3_X1  g451(.A1(new_n650_), .A2(new_n512_), .A3(new_n553_), .ZN(new_n653_));
  INV_X1    g452(.A(G57gat), .ZN(new_n654_));
  NOR3_X1   g453(.A1(new_n653_), .A2(new_n654_), .A3(new_n238_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n652_), .A2(new_n655_), .ZN(G1332gat));
  OAI21_X1  g455(.A(G64gat), .B1(new_n653_), .B2(new_n559_), .ZN(new_n657_));
  XNOR2_X1  g456(.A(new_n657_), .B(KEYINPUT48), .ZN(new_n658_));
  INV_X1    g457(.A(G64gat), .ZN(new_n659_));
  NAND3_X1  g458(.A1(new_n651_), .A2(new_n659_), .A3(new_n560_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n658_), .A2(new_n660_), .ZN(G1333gat));
  OAI21_X1  g460(.A(G71gat), .B1(new_n653_), .B2(new_n475_), .ZN(new_n662_));
  XNOR2_X1  g461(.A(new_n662_), .B(KEYINPUT49), .ZN(new_n663_));
  INV_X1    g462(.A(G71gat), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n651_), .A2(new_n664_), .A3(new_n637_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n663_), .A2(new_n665_), .ZN(G1334gat));
  NAND4_X1  g465(.A1(new_n650_), .A2(new_n512_), .A3(new_n464_), .A4(new_n553_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G78gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G78gat), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT50), .ZN(new_n671_));
  OR3_X1    g470(.A1(new_n669_), .A2(new_n670_), .A3(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(new_n671_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n673_));
  INV_X1    g472(.A(G78gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n651_), .A2(new_n674_), .A3(new_n464_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n672_), .A2(new_n673_), .A3(new_n675_), .ZN(new_n676_));
  XNOR2_X1  g475(.A(new_n676_), .B(KEYINPUT106), .ZN(G1335gat));
  NAND2_X1  g476(.A1(new_n650_), .A2(new_n612_), .ZN(new_n678_));
  INV_X1    g477(.A(new_n678_), .ZN(new_n679_));
  AOI21_X1  g478(.A(G85gat), .B1(new_n679_), .B2(new_n239_), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n608_), .A2(new_n649_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n239_), .A2(G85gat), .ZN(new_n682_));
  AOI21_X1  g481(.A(new_n680_), .B1(new_n681_), .B2(new_n682_), .ZN(G1336gat));
  NOR3_X1   g482(.A1(new_n678_), .A2(G92gat), .A3(new_n559_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n681_), .A2(new_n560_), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n684_), .B1(new_n685_), .B2(G92gat), .ZN(new_n686_));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1337gat));
  NAND2_X1  g487(.A1(new_n681_), .A2(new_n637_), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n689_), .A2(G99gat), .ZN(new_n690_));
  NAND3_X1  g489(.A1(new_n679_), .A2(new_n241_), .A3(new_n637_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n690_), .A2(new_n691_), .ZN(new_n692_));
  XNOR2_X1  g491(.A(new_n692_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g492(.A1(new_n679_), .A2(new_n242_), .A3(new_n464_), .ZN(new_n694_));
  NAND3_X1  g493(.A1(new_n608_), .A2(new_n464_), .A3(new_n649_), .ZN(new_n695_));
  INV_X1    g494(.A(KEYINPUT52), .ZN(new_n696_));
  AND3_X1   g495(.A1(new_n695_), .A2(new_n696_), .A3(G106gat), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n695_), .B2(G106gat), .ZN(new_n698_));
  OAI21_X1  g497(.A(new_n694_), .B1(new_n697_), .B2(new_n698_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(new_n699_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g499(.A(KEYINPUT116), .ZN(new_n701_));
  INV_X1    g500(.A(KEYINPUT110), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT55), .ZN(new_n703_));
  AOI21_X1  g502(.A(new_n702_), .B1(new_n307_), .B2(new_n703_), .ZN(new_n704_));
  AOI211_X1 g503(.A(KEYINPUT110), .B(KEYINPUT55), .C1(new_n305_), .C2(new_n306_), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  NAND3_X1  g505(.A1(new_n292_), .A2(new_n308_), .A3(new_n302_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n707_), .A2(new_n293_), .ZN(new_n708_));
  NAND2_X1  g507(.A1(new_n708_), .A2(KEYINPUT111), .ZN(new_n709_));
  INV_X1    g508(.A(KEYINPUT111), .ZN(new_n710_));
  NAND3_X1  g509(.A1(new_n707_), .A2(new_n710_), .A3(new_n293_), .ZN(new_n711_));
  AND2_X1   g510(.A1(new_n292_), .A2(new_n302_), .ZN(new_n712_));
  NAND4_X1  g511(.A1(new_n712_), .A2(KEYINPUT112), .A3(KEYINPUT55), .A4(new_n294_), .ZN(new_n713_));
  INV_X1    g512(.A(KEYINPUT112), .ZN(new_n714_));
  OAI21_X1  g513(.A(new_n714_), .B1(new_n303_), .B2(new_n703_), .ZN(new_n715_));
  AOI22_X1  g514(.A1(new_n709_), .A2(new_n711_), .B1(new_n713_), .B2(new_n715_), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n319_), .B1(new_n706_), .B2(new_n716_), .ZN(new_n717_));
  OAI21_X1  g516(.A(new_n701_), .B1(new_n717_), .B2(KEYINPUT56), .ZN(new_n718_));
  NAND2_X1  g517(.A1(new_n307_), .A2(new_n703_), .ZN(new_n719_));
  NAND2_X1  g518(.A1(new_n719_), .A2(KEYINPUT110), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n307_), .A2(new_n702_), .A3(new_n703_), .ZN(new_n721_));
  NAND3_X1  g520(.A1(new_n720_), .A2(new_n721_), .A3(new_n716_), .ZN(new_n722_));
  INV_X1    g521(.A(new_n319_), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n722_), .A2(KEYINPUT56), .A3(new_n723_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n724_), .A2(KEYINPUT115), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT115), .ZN(new_n726_));
  NAND4_X1  g525(.A1(new_n722_), .A2(new_n726_), .A3(KEYINPUT56), .A4(new_n723_), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT56), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n709_), .A2(new_n711_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n713_), .A2(new_n715_), .ZN(new_n730_));
  NAND2_X1  g529(.A1(new_n729_), .A2(new_n730_), .ZN(new_n731_));
  NOR3_X1   g530(.A1(new_n731_), .A2(new_n704_), .A3(new_n705_), .ZN(new_n732_));
  OAI211_X1 g531(.A(KEYINPUT116), .B(new_n728_), .C1(new_n732_), .C2(new_n319_), .ZN(new_n733_));
  NAND4_X1  g532(.A1(new_n718_), .A2(new_n725_), .A3(new_n727_), .A4(new_n733_), .ZN(new_n734_));
  NOR2_X1   g533(.A1(KEYINPUT117), .A2(KEYINPUT58), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n359_), .A2(new_n361_), .A3(new_n355_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n351_), .A2(new_n362_), .A3(new_n353_), .ZN(new_n737_));
  NAND3_X1  g536(.A1(new_n736_), .A2(new_n737_), .A3(new_n371_), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n374_), .A2(new_n738_), .ZN(new_n739_));
  XNOR2_X1  g538(.A(new_n739_), .B(KEYINPUT113), .ZN(new_n740_));
  AND2_X1   g539(.A1(new_n740_), .A2(new_n318_), .ZN(new_n741_));
  AND3_X1   g540(.A1(new_n734_), .A2(new_n735_), .A3(new_n741_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n735_), .B1(new_n734_), .B2(new_n741_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n596_), .B1(new_n742_), .B2(new_n743_), .ZN(new_n744_));
  XNOR2_X1  g543(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n318_), .A2(new_n375_), .ZN(new_n746_));
  INV_X1    g545(.A(KEYINPUT109), .ZN(new_n747_));
  XNOR2_X1  g546(.A(new_n746_), .B(new_n747_), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n728_), .B1(new_n732_), .B2(new_n319_), .ZN(new_n749_));
  NAND2_X1  g548(.A1(new_n749_), .A2(new_n724_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n748_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n740_), .A2(new_n320_), .ZN(new_n752_));
  AND2_X1   g551(.A1(new_n751_), .A2(new_n752_), .ZN(new_n753_));
  OAI21_X1  g552(.A(new_n745_), .B1(new_n753_), .B2(new_n536_), .ZN(new_n754_));
  NAND2_X1  g553(.A1(new_n744_), .A2(new_n754_), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n536_), .B1(new_n751_), .B2(new_n752_), .ZN(new_n756_));
  NAND2_X1  g555(.A1(new_n756_), .A2(KEYINPUT57), .ZN(new_n757_));
  INV_X1    g556(.A(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n513_), .B1(new_n755_), .B2(new_n758_), .ZN(new_n759_));
  INV_X1    g558(.A(KEYINPUT54), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n761_));
  NOR2_X1   g560(.A1(new_n324_), .A2(new_n375_), .ZN(new_n762_));
  NAND3_X1  g561(.A1(new_n546_), .A2(new_n761_), .A3(new_n762_), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  AOI21_X1  g563(.A(new_n761_), .B1(new_n546_), .B2(new_n762_), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n760_), .B1(new_n764_), .B2(new_n765_), .ZN(new_n766_));
  INV_X1    g565(.A(new_n765_), .ZN(new_n767_));
  NAND3_X1  g566(.A1(new_n767_), .A2(KEYINPUT54), .A3(new_n763_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n766_), .A2(new_n768_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n759_), .A2(new_n769_), .ZN(new_n770_));
  NAND2_X1  g569(.A1(new_n239_), .A2(new_n559_), .ZN(new_n771_));
  INV_X1    g570(.A(new_n476_), .ZN(new_n772_));
  NOR2_X1   g571(.A1(new_n771_), .A2(new_n772_), .ZN(new_n773_));
  NAND2_X1  g572(.A1(new_n770_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(new_n774_), .ZN(new_n775_));
  AOI21_X1  g574(.A(G113gat), .B1(new_n775_), .B2(new_n375_), .ZN(new_n776_));
  INV_X1    g575(.A(KEYINPUT59), .ZN(new_n777_));
  AOI21_X1  g576(.A(new_n758_), .B1(new_n755_), .B2(KEYINPUT118), .ZN(new_n778_));
  INV_X1    g577(.A(KEYINPUT118), .ZN(new_n779_));
  NAND3_X1  g578(.A1(new_n744_), .A2(new_n779_), .A3(new_n754_), .ZN(new_n780_));
  AOI21_X1  g579(.A(new_n512_), .B1(new_n778_), .B2(new_n780_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n769_), .ZN(new_n782_));
  OAI211_X1 g581(.A(new_n777_), .B(new_n773_), .C1(new_n781_), .C2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT119), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n774_), .A2(KEYINPUT59), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n734_), .A2(new_n741_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n735_), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND3_X1  g588(.A1(new_n734_), .A2(new_n735_), .A3(new_n741_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n595_), .B1(new_n789_), .B2(new_n790_), .ZN(new_n791_));
  INV_X1    g590(.A(new_n745_), .ZN(new_n792_));
  NOR2_X1   g591(.A1(new_n756_), .A2(new_n792_), .ZN(new_n793_));
  OAI21_X1  g592(.A(KEYINPUT118), .B1(new_n791_), .B2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(new_n757_), .A3(new_n780_), .ZN(new_n795_));
  NAND2_X1  g594(.A1(new_n795_), .A2(new_n513_), .ZN(new_n796_));
  NAND2_X1  g595(.A1(new_n796_), .A2(new_n769_), .ZN(new_n797_));
  NAND4_X1  g596(.A1(new_n797_), .A2(KEYINPUT119), .A3(new_n777_), .A4(new_n773_), .ZN(new_n798_));
  AND4_X1   g597(.A1(new_n375_), .A2(new_n785_), .A3(new_n786_), .A4(new_n798_), .ZN(new_n799_));
  AOI21_X1  g598(.A(new_n776_), .B1(new_n799_), .B2(G113gat), .ZN(G1340gat));
  NAND4_X1  g599(.A1(new_n785_), .A2(new_n324_), .A3(new_n798_), .A4(new_n786_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(G120gat), .ZN(new_n802_));
  OAI21_X1  g601(.A(new_n205_), .B1(new_n648_), .B2(KEYINPUT60), .ZN(new_n803_));
  OAI211_X1 g602(.A(new_n775_), .B(new_n803_), .C1(KEYINPUT60), .C2(new_n205_), .ZN(new_n804_));
  NAND2_X1  g603(.A1(new_n802_), .A2(new_n804_), .ZN(G1341gat));
  AOI21_X1  g604(.A(G127gat), .B1(new_n775_), .B2(new_n512_), .ZN(new_n806_));
  AND4_X1   g605(.A1(G127gat), .A2(new_n785_), .A3(new_n786_), .A4(new_n798_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n806_), .B1(new_n807_), .B2(new_n512_), .ZN(G1342gat));
  AOI21_X1  g607(.A(G134gat), .B1(new_n775_), .B2(new_n536_), .ZN(new_n809_));
  AND4_X1   g608(.A1(G134gat), .A2(new_n785_), .A3(new_n786_), .A4(new_n798_), .ZN(new_n810_));
  AOI21_X1  g609(.A(new_n809_), .B1(new_n810_), .B2(new_n596_), .ZN(G1343gat));
  AOI21_X1  g610(.A(new_n637_), .B1(new_n759_), .B2(new_n769_), .ZN(new_n812_));
  NOR2_X1   g611(.A1(new_n771_), .A2(new_n590_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n812_), .A2(new_n813_), .ZN(new_n814_));
  NAND2_X1  g613(.A1(new_n814_), .A2(new_n375_), .ZN(new_n815_));
  XNOR2_X1  g614(.A(KEYINPUT120), .B(G141gat), .ZN(new_n816_));
  XNOR2_X1  g615(.A(new_n815_), .B(new_n816_), .ZN(G1344gat));
  NAND2_X1  g616(.A1(new_n814_), .A2(new_n324_), .ZN(new_n818_));
  XNOR2_X1  g617(.A(new_n818_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g618(.A1(new_n814_), .A2(new_n512_), .ZN(new_n820_));
  XOR2_X1   g619(.A(KEYINPUT61), .B(G155gat), .Z(new_n821_));
  XNOR2_X1  g620(.A(new_n821_), .B(KEYINPUT121), .ZN(new_n822_));
  XNOR2_X1  g621(.A(new_n820_), .B(new_n822_), .ZN(G1346gat));
  NAND3_X1  g622(.A1(new_n814_), .A2(G162gat), .A3(new_n596_), .ZN(new_n824_));
  NAND4_X1  g623(.A1(new_n770_), .A2(new_n475_), .A3(new_n536_), .A4(new_n813_), .ZN(new_n825_));
  AND3_X1   g624(.A1(new_n825_), .A2(KEYINPUT122), .A3(new_n527_), .ZN(new_n826_));
  AOI21_X1  g625(.A(KEYINPUT122), .B1(new_n825_), .B2(new_n527_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n824_), .B1(new_n826_), .B2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(KEYINPUT123), .ZN(new_n829_));
  NAND2_X1  g628(.A1(new_n828_), .A2(new_n829_), .ZN(new_n830_));
  OAI211_X1 g629(.A(new_n824_), .B(KEYINPUT123), .C1(new_n826_), .C2(new_n827_), .ZN(new_n831_));
  NAND2_X1  g630(.A1(new_n830_), .A2(new_n831_), .ZN(G1347gat));
  INV_X1    g631(.A(KEYINPUT124), .ZN(new_n833_));
  NOR3_X1   g632(.A1(new_n239_), .A2(new_n559_), .A3(new_n772_), .ZN(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  AOI211_X1 g634(.A(new_n376_), .B(new_n835_), .C1(new_n796_), .C2(new_n769_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n833_), .B1(new_n836_), .B2(new_n368_), .ZN(new_n837_));
  NAND2_X1  g636(.A1(new_n797_), .A2(new_n834_), .ZN(new_n838_));
  OAI211_X1 g637(.A(KEYINPUT124), .B(G169gat), .C1(new_n838_), .C2(new_n376_), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n837_), .A2(new_n839_), .A3(KEYINPUT62), .ZN(new_n840_));
  NAND3_X1  g639(.A1(new_n836_), .A2(new_n386_), .A3(new_n384_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT62), .ZN(new_n842_));
  OAI211_X1 g641(.A(new_n833_), .B(new_n842_), .C1(new_n836_), .C2(new_n368_), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n840_), .A2(new_n841_), .A3(new_n843_), .ZN(G1348gat));
  NAND2_X1  g643(.A1(new_n770_), .A2(new_n834_), .ZN(new_n845_));
  NOR3_X1   g644(.A1(new_n845_), .A2(new_n316_), .A3(new_n648_), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n797_), .A2(new_n324_), .A3(new_n834_), .ZN(new_n847_));
  AOI21_X1  g646(.A(new_n846_), .B1(new_n847_), .B2(new_n316_), .ZN(G1349gat));
  NOR2_X1   g647(.A1(new_n845_), .A2(new_n513_), .ZN(new_n849_));
  MUX2_X1   g648(.A(G183gat), .B(new_n401_), .S(new_n849_), .Z(G1350gat));
  OAI21_X1  g649(.A(G190gat), .B1(new_n838_), .B2(new_n595_), .ZN(new_n851_));
  NAND2_X1  g650(.A1(new_n536_), .A2(new_n418_), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n852_), .B(KEYINPUT125), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n851_), .B1(new_n838_), .B2(new_n853_), .ZN(G1351gat));
  AND2_X1   g653(.A1(new_n812_), .A2(new_n560_), .ZN(new_n855_));
  NOR2_X1   g654(.A1(new_n239_), .A2(new_n590_), .ZN(new_n856_));
  AND2_X1   g655(.A1(new_n855_), .A2(new_n856_), .ZN(new_n857_));
  NAND2_X1  g656(.A1(new_n857_), .A2(new_n375_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(G197gat), .ZN(new_n859_));
  NAND3_X1  g658(.A1(new_n857_), .A2(new_n370_), .A3(new_n375_), .ZN(new_n860_));
  NAND2_X1  g659(.A1(new_n859_), .A2(new_n860_), .ZN(G1352gat));
  NAND3_X1  g660(.A1(new_n855_), .A2(new_n324_), .A3(new_n856_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g662(.A1(new_n812_), .A2(new_n512_), .A3(new_n856_), .A4(new_n560_), .ZN(new_n864_));
  AND2_X1   g663(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n865_));
  NOR2_X1   g664(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n866_));
  NOR3_X1   g665(.A1(new_n864_), .A2(new_n865_), .A3(new_n866_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT126), .ZN(new_n868_));
  AOI21_X1  g667(.A(new_n868_), .B1(new_n864_), .B2(new_n866_), .ZN(new_n869_));
  NOR2_X1   g668(.A1(new_n867_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n870_), .B1(KEYINPUT126), .B2(new_n867_), .ZN(G1354gat));
  NAND4_X1  g670(.A1(new_n812_), .A2(new_n856_), .A3(new_n560_), .A4(new_n536_), .ZN(new_n872_));
  OR2_X1    g671(.A1(new_n872_), .A2(KEYINPUT127), .ZN(new_n873_));
  INV_X1    g672(.A(G218gat), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n872_), .A2(KEYINPUT127), .ZN(new_n875_));
  NAND3_X1  g674(.A1(new_n873_), .A2(new_n874_), .A3(new_n875_), .ZN(new_n876_));
  NAND3_X1  g675(.A1(new_n857_), .A2(G218gat), .A3(new_n596_), .ZN(new_n877_));
  AND2_X1   g676(.A1(new_n876_), .A2(new_n877_), .ZN(G1355gat));
endmodule


