//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:30:50 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n640_, new_n641_,
    new_n642_, new_n644_, new_n645_, new_n646_, new_n647_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n721_, new_n722_,
    new_n723_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n741_, new_n742_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n748_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n838_, new_n839_, new_n840_, new_n842_, new_n843_, new_n844_,
    new_n846_, new_n847_, new_n848_, new_n849_, new_n851_, new_n852_,
    new_n854_, new_n855_, new_n857_, new_n858_, new_n859_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n871_, new_n872_, new_n873_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n881_, new_n882_,
    new_n883_, new_n884_, new_n885_, new_n886_, new_n888_, new_n889_,
    new_n891_, new_n893_, new_n894_, new_n895_, new_n896_, new_n898_,
    new_n899_, new_n900_;
  NOR2_X1   g000(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n202_));
  INV_X1    g001(.A(new_n202_), .ZN(new_n203_));
  NAND2_X1  g002(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n204_));
  NAND3_X1  g003(.A1(new_n203_), .A2(KEYINPUT64), .A3(new_n204_), .ZN(new_n205_));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n206_));
  AND2_X1   g005(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n207_));
  OAI21_X1  g006(.A(new_n206_), .B1(new_n207_), .B2(new_n202_), .ZN(new_n208_));
  AOI21_X1  g007(.A(G106gat), .B1(new_n205_), .B2(new_n208_), .ZN(new_n209_));
  NAND2_X1  g008(.A1(G99gat), .A2(G106gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n211_));
  INV_X1    g010(.A(KEYINPUT6), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n212_), .A2(G99gat), .A3(G106gat), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n211_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(G85gat), .ZN(new_n215_));
  INV_X1    g014(.A(G92gat), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(G85gat), .A2(G92gat), .ZN(new_n218_));
  NAND3_X1  g017(.A1(new_n217_), .A2(KEYINPUT9), .A3(new_n218_), .ZN(new_n219_));
  OR2_X1    g018(.A1(new_n218_), .A2(KEYINPUT9), .ZN(new_n220_));
  NAND3_X1  g019(.A1(new_n214_), .A2(new_n219_), .A3(new_n220_), .ZN(new_n221_));
  OR2_X1    g020(.A1(new_n209_), .A2(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT7), .ZN(new_n225_));
  INV_X1    g024(.A(G99gat), .ZN(new_n226_));
  INV_X1    g025(.A(G106gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n225_), .A2(new_n226_), .A3(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n212_), .B1(G99gat), .B2(G106gat), .ZN(new_n229_));
  NOR2_X1   g028(.A1(new_n210_), .A2(KEYINPUT6), .ZN(new_n230_));
  OAI211_X1 g029(.A(new_n224_), .B(new_n228_), .C1(new_n229_), .C2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n232_));
  AND2_X1   g031(.A1(G85gat), .A2(G92gat), .ZN(new_n233_));
  NOR2_X1   g032(.A1(G85gat), .A2(G92gat), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n232_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  NAND3_X1  g034(.A1(new_n217_), .A2(KEYINPUT65), .A3(new_n218_), .ZN(new_n236_));
  AND4_X1   g035(.A1(new_n223_), .A2(new_n231_), .A3(new_n235_), .A4(new_n236_), .ZN(new_n237_));
  AND2_X1   g036(.A1(new_n235_), .A2(new_n236_), .ZN(new_n238_));
  AOI21_X1  g037(.A(new_n223_), .B1(new_n238_), .B2(new_n231_), .ZN(new_n239_));
  OAI21_X1  g038(.A(new_n222_), .B1(new_n237_), .B2(new_n239_), .ZN(new_n240_));
  NAND2_X1  g039(.A1(new_n240_), .A2(KEYINPUT69), .ZN(new_n241_));
  XNOR2_X1  g040(.A(G29gat), .B(G36gat), .ZN(new_n242_));
  XNOR2_X1  g041(.A(G43gat), .B(G50gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n244_), .B(KEYINPUT15), .ZN(new_n245_));
  AND2_X1   g044(.A1(new_n211_), .A2(new_n213_), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n228_), .A2(new_n224_), .ZN(new_n247_));
  NOR2_X1   g046(.A1(new_n246_), .A2(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(new_n235_), .A2(new_n236_), .ZN(new_n249_));
  OAI21_X1  g048(.A(KEYINPUT8), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n238_), .A2(new_n223_), .A3(new_n231_), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n250_), .A2(new_n251_), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n252_), .A2(new_n253_), .A3(new_n222_), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n241_), .A2(new_n245_), .A3(new_n254_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n240_), .A2(KEYINPUT66), .ZN(new_n256_));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n257_));
  NAND3_X1  g056(.A1(new_n252_), .A2(new_n257_), .A3(new_n222_), .ZN(new_n258_));
  NAND3_X1  g057(.A1(new_n256_), .A2(new_n244_), .A3(new_n258_), .ZN(new_n259_));
  NAND2_X1  g058(.A1(G232gat), .A2(G233gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n260_), .B(KEYINPUT34), .ZN(new_n261_));
  XOR2_X1   g060(.A(new_n261_), .B(KEYINPUT35), .Z(new_n262_));
  NAND4_X1  g061(.A1(new_n255_), .A2(new_n259_), .A3(KEYINPUT75), .A4(new_n262_), .ZN(new_n263_));
  NAND3_X1  g062(.A1(new_n255_), .A2(new_n259_), .A3(new_n262_), .ZN(new_n264_));
  INV_X1    g063(.A(KEYINPUT75), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n264_), .A2(new_n265_), .ZN(new_n266_));
  NAND2_X1  g065(.A1(new_n261_), .A2(KEYINPUT35), .ZN(new_n267_));
  AOI21_X1  g066(.A(new_n267_), .B1(new_n255_), .B2(new_n259_), .ZN(new_n268_));
  OAI21_X1  g067(.A(new_n263_), .B1(new_n266_), .B2(new_n268_), .ZN(new_n269_));
  XOR2_X1   g068(.A(G190gat), .B(G218gat), .Z(new_n270_));
  XNOR2_X1  g069(.A(G134gat), .B(G162gat), .ZN(new_n271_));
  OR2_X1    g070(.A1(new_n270_), .A2(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n270_), .A2(new_n271_), .ZN(new_n273_));
  AOI21_X1  g072(.A(KEYINPUT36), .B1(new_n272_), .B2(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT74), .ZN(new_n275_));
  NAND3_X1  g074(.A1(new_n269_), .A2(KEYINPUT76), .A3(new_n275_), .ZN(new_n276_));
  AND3_X1   g075(.A1(new_n272_), .A2(KEYINPUT36), .A3(new_n273_), .ZN(new_n277_));
  NOR2_X1   g076(.A1(new_n277_), .A2(new_n274_), .ZN(new_n278_));
  OAI211_X1 g077(.A(new_n263_), .B(new_n278_), .C1(new_n266_), .C2(new_n268_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n276_), .A2(new_n279_), .ZN(new_n280_));
  AOI21_X1  g079(.A(KEYINPUT76), .B1(new_n269_), .B2(new_n275_), .ZN(new_n281_));
  OAI21_X1  g080(.A(KEYINPUT37), .B1(new_n280_), .B2(new_n281_), .ZN(new_n282_));
  INV_X1    g081(.A(KEYINPUT78), .ZN(new_n283_));
  NAND2_X1  g082(.A1(new_n269_), .A2(KEYINPUT77), .ZN(new_n284_));
  INV_X1    g083(.A(KEYINPUT77), .ZN(new_n285_));
  OAI211_X1 g084(.A(new_n285_), .B(new_n263_), .C1(new_n266_), .C2(new_n268_), .ZN(new_n286_));
  NAND3_X1  g085(.A1(new_n284_), .A2(new_n278_), .A3(new_n286_), .ZN(new_n287_));
  INV_X1    g086(.A(KEYINPUT37), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n269_), .A2(new_n275_), .ZN(new_n289_));
  NAND3_X1  g088(.A1(new_n287_), .A2(new_n288_), .A3(new_n289_), .ZN(new_n290_));
  AND3_X1   g089(.A1(new_n282_), .A2(new_n283_), .A3(new_n290_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n283_), .B1(new_n282_), .B2(new_n290_), .ZN(new_n292_));
  OR2_X1    g091(.A1(new_n291_), .A2(new_n292_), .ZN(new_n293_));
  XOR2_X1   g092(.A(G127gat), .B(G155gat), .Z(new_n294_));
  XNOR2_X1  g093(.A(new_n294_), .B(KEYINPUT16), .ZN(new_n295_));
  XNOR2_X1  g094(.A(G183gat), .B(G211gat), .ZN(new_n296_));
  XNOR2_X1  g095(.A(new_n295_), .B(new_n296_), .ZN(new_n297_));
  XNOR2_X1  g096(.A(G1gat), .B(G8gat), .ZN(new_n298_));
  INV_X1    g097(.A(KEYINPUT79), .ZN(new_n299_));
  XNOR2_X1  g098(.A(new_n298_), .B(new_n299_), .ZN(new_n300_));
  INV_X1    g099(.A(G15gat), .ZN(new_n301_));
  INV_X1    g100(.A(G22gat), .ZN(new_n302_));
  NAND2_X1  g101(.A1(new_n301_), .A2(new_n302_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G15gat), .A2(G22gat), .ZN(new_n304_));
  NAND2_X1  g103(.A1(G1gat), .A2(G8gat), .ZN(new_n305_));
  AOI22_X1  g104(.A1(new_n303_), .A2(new_n304_), .B1(KEYINPUT14), .B2(new_n305_), .ZN(new_n306_));
  XNOR2_X1  g105(.A(new_n300_), .B(new_n306_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(G231gat), .A2(G233gat), .ZN(new_n308_));
  XOR2_X1   g107(.A(new_n308_), .B(KEYINPUT80), .Z(new_n309_));
  XNOR2_X1  g108(.A(new_n307_), .B(new_n309_), .ZN(new_n310_));
  XNOR2_X1  g109(.A(KEYINPUT67), .B(G71gat), .ZN(new_n311_));
  INV_X1    g110(.A(G78gat), .ZN(new_n312_));
  XNOR2_X1  g111(.A(new_n311_), .B(new_n312_), .ZN(new_n313_));
  XNOR2_X1  g112(.A(G57gat), .B(G64gat), .ZN(new_n314_));
  AND2_X1   g113(.A1(new_n314_), .A2(KEYINPUT11), .ZN(new_n315_));
  OR2_X1    g114(.A1(new_n313_), .A2(new_n315_), .ZN(new_n316_));
  NOR2_X1   g115(.A1(new_n314_), .A2(KEYINPUT11), .ZN(new_n317_));
  OAI21_X1  g116(.A(new_n313_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  AND2_X1   g117(.A1(new_n316_), .A2(new_n318_), .ZN(new_n319_));
  XNOR2_X1  g118(.A(new_n310_), .B(new_n319_), .ZN(new_n320_));
  OAI21_X1  g119(.A(new_n297_), .B1(new_n320_), .B2(KEYINPUT17), .ZN(new_n321_));
  OAI21_X1  g120(.A(new_n321_), .B1(KEYINPUT17), .B2(new_n297_), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n320_), .A2(KEYINPUT81), .ZN(new_n323_));
  XNOR2_X1  g122(.A(new_n322_), .B(new_n323_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n316_), .A2(new_n318_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n209_), .A2(new_n221_), .ZN(new_n326_));
  AOI211_X1 g125(.A(KEYINPUT66), .B(new_n326_), .C1(new_n250_), .C2(new_n251_), .ZN(new_n327_));
  AOI21_X1  g126(.A(new_n257_), .B1(new_n252_), .B2(new_n222_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n325_), .B1(new_n327_), .B2(new_n328_), .ZN(new_n329_));
  XNOR2_X1  g128(.A(KEYINPUT71), .B(KEYINPUT12), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT12), .ZN(new_n333_));
  AOI21_X1  g132(.A(new_n333_), .B1(new_n316_), .B2(new_n318_), .ZN(new_n334_));
  NAND4_X1  g133(.A1(new_n241_), .A2(new_n332_), .A3(new_n254_), .A4(new_n334_), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n241_), .A2(new_n254_), .A3(new_n334_), .ZN(new_n336_));
  NAND2_X1  g135(.A1(new_n336_), .A2(KEYINPUT70), .ZN(new_n337_));
  AND3_X1   g136(.A1(new_n331_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n256_), .A2(new_n258_), .A3(new_n319_), .ZN(new_n339_));
  NAND2_X1  g138(.A1(G230gat), .A2(G233gat), .ZN(new_n340_));
  NAND2_X1  g139(.A1(new_n339_), .A2(new_n340_), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n339_), .A2(KEYINPUT72), .A3(new_n340_), .ZN(new_n344_));
  NAND2_X1  g143(.A1(new_n343_), .A2(new_n344_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n338_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(new_n340_), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT68), .ZN(new_n348_));
  XNOR2_X1  g147(.A(new_n339_), .B(new_n348_), .ZN(new_n349_));
  INV_X1    g148(.A(new_n329_), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n347_), .B1(new_n349_), .B2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(new_n346_), .A2(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G120gat), .B(G148gat), .ZN(new_n353_));
  XNOR2_X1  g152(.A(new_n353_), .B(KEYINPUT5), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G176gat), .B(G204gat), .ZN(new_n355_));
  XOR2_X1   g154(.A(new_n354_), .B(new_n355_), .Z(new_n356_));
  NAND2_X1  g155(.A1(new_n352_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(new_n356_), .ZN(new_n358_));
  NAND3_X1  g157(.A1(new_n346_), .A2(new_n351_), .A3(new_n358_), .ZN(new_n359_));
  NAND2_X1  g158(.A1(new_n357_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT73), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n360_), .B1(new_n361_), .B2(KEYINPUT13), .ZN(new_n362_));
  XOR2_X1   g161(.A(KEYINPUT73), .B(KEYINPUT13), .Z(new_n363_));
  NAND3_X1  g162(.A1(new_n357_), .A2(new_n359_), .A3(new_n363_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n293_), .A2(new_n324_), .A3(new_n365_), .ZN(new_n366_));
  INV_X1    g165(.A(new_n366_), .ZN(new_n367_));
  INV_X1    g166(.A(KEYINPUT99), .ZN(new_n368_));
  INV_X1    g167(.A(KEYINPUT20), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT87), .ZN(new_n370_));
  INV_X1    g169(.A(G169gat), .ZN(new_n371_));
  OAI21_X1  g170(.A(KEYINPUT22), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(G176gat), .ZN(new_n373_));
  NAND2_X1  g172(.A1(new_n372_), .A2(new_n373_), .ZN(new_n374_));
  NOR3_X1   g173(.A1(new_n370_), .A2(new_n371_), .A3(KEYINPUT22), .ZN(new_n375_));
  OAI22_X1  g174(.A1(new_n374_), .A2(new_n375_), .B1(new_n371_), .B2(new_n373_), .ZN(new_n376_));
  AOI21_X1  g175(.A(KEYINPUT23), .B1(G183gat), .B2(G190gat), .ZN(new_n377_));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378_));
  XNOR2_X1  g177(.A(new_n378_), .B(KEYINPUT86), .ZN(new_n379_));
  AOI21_X1  g178(.A(new_n377_), .B1(new_n379_), .B2(KEYINPUT23), .ZN(new_n380_));
  NOR2_X1   g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381_));
  INV_X1    g180(.A(new_n381_), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n376_), .B1(new_n380_), .B2(new_n382_), .ZN(new_n383_));
  XNOR2_X1  g182(.A(KEYINPUT25), .B(G183gat), .ZN(new_n384_));
  XNOR2_X1  g183(.A(KEYINPUT26), .B(G190gat), .ZN(new_n385_));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386_));
  NOR2_X1   g185(.A1(G169gat), .A2(G176gat), .ZN(new_n387_));
  AOI22_X1  g186(.A1(new_n384_), .A2(new_n385_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n371_), .A2(new_n373_), .ZN(new_n389_));
  OR3_X1    g188(.A1(new_n389_), .A2(new_n386_), .A3(new_n387_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n388_), .A2(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n392_), .B1(G183gat), .B2(G190gat), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n393_), .B1(new_n379_), .B2(new_n392_), .ZN(new_n394_));
  NOR2_X1   g193(.A1(new_n391_), .A2(new_n394_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n383_), .A2(new_n395_), .ZN(new_n396_));
  INV_X1    g195(.A(G197gat), .ZN(new_n397_));
  NOR2_X1   g196(.A1(new_n397_), .A2(G204gat), .ZN(new_n398_));
  INV_X1    g197(.A(G204gat), .ZN(new_n399_));
  NOR2_X1   g198(.A1(new_n399_), .A2(G197gat), .ZN(new_n400_));
  OAI21_X1  g199(.A(KEYINPUT21), .B1(new_n398_), .B2(new_n400_), .ZN(new_n401_));
  XNOR2_X1  g200(.A(G211gat), .B(G218gat), .ZN(new_n402_));
  OAI21_X1  g201(.A(KEYINPUT92), .B1(new_n397_), .B2(G204gat), .ZN(new_n403_));
  INV_X1    g202(.A(KEYINPUT92), .ZN(new_n404_));
  NAND3_X1  g203(.A1(new_n404_), .A2(new_n399_), .A3(G197gat), .ZN(new_n405_));
  OAI211_X1 g204(.A(new_n403_), .B(new_n405_), .C1(G197gat), .C2(new_n399_), .ZN(new_n406_));
  OAI211_X1 g205(.A(new_n401_), .B(new_n402_), .C1(new_n406_), .C2(KEYINPUT21), .ZN(new_n407_));
  INV_X1    g206(.A(new_n402_), .ZN(new_n408_));
  NAND3_X1  g207(.A1(new_n406_), .A2(KEYINPUT21), .A3(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n407_), .A2(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n369_), .B1(new_n396_), .B2(new_n411_), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n413_));
  XNOR2_X1  g212(.A(new_n378_), .B(new_n413_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n414_), .A2(KEYINPUT23), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n382_), .B1(new_n415_), .B2(new_n393_), .ZN(new_n416_));
  XNOR2_X1  g215(.A(KEYINPUT22), .B(G169gat), .ZN(new_n417_));
  AOI21_X1  g216(.A(new_n389_), .B1(new_n417_), .B2(new_n373_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n388_), .A2(new_n390_), .ZN(new_n419_));
  AOI22_X1  g218(.A1(new_n416_), .A2(new_n418_), .B1(new_n419_), .B2(new_n380_), .ZN(new_n420_));
  OAI21_X1  g219(.A(KEYINPUT95), .B1(new_n420_), .B2(new_n411_), .ZN(new_n421_));
  XNOR2_X1  g220(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n422_));
  NAND2_X1  g221(.A1(G226gat), .A2(G233gat), .ZN(new_n423_));
  XNOR2_X1  g222(.A(new_n422_), .B(new_n423_), .ZN(new_n424_));
  NAND2_X1  g223(.A1(new_n419_), .A2(new_n380_), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n418_), .B1(new_n394_), .B2(new_n381_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n425_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(KEYINPUT95), .ZN(new_n428_));
  NAND3_X1  g227(.A1(new_n427_), .A2(new_n428_), .A3(new_n410_), .ZN(new_n429_));
  NAND4_X1  g228(.A1(new_n412_), .A2(new_n421_), .A3(new_n424_), .A4(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n411_), .A2(new_n425_), .A3(new_n426_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n410_), .B1(new_n383_), .B2(new_n395_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n431_), .A2(new_n432_), .A3(KEYINPUT20), .ZN(new_n433_));
  INV_X1    g232(.A(new_n424_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n433_), .A2(new_n434_), .ZN(new_n435_));
  NAND2_X1  g234(.A1(new_n430_), .A2(new_n435_), .ZN(new_n436_));
  XOR2_X1   g235(.A(G8gat), .B(G36gat), .Z(new_n437_));
  XNOR2_X1  g236(.A(new_n437_), .B(KEYINPUT18), .ZN(new_n438_));
  XNOR2_X1  g237(.A(G64gat), .B(G92gat), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n438_), .B(new_n439_), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  AOI21_X1  g240(.A(new_n368_), .B1(new_n436_), .B2(new_n441_), .ZN(new_n442_));
  AOI211_X1 g241(.A(KEYINPUT99), .B(new_n440_), .C1(new_n430_), .C2(new_n435_), .ZN(new_n443_));
  OR2_X1    g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(KEYINPUT27), .ZN(new_n445_));
  NOR2_X1   g244(.A1(new_n433_), .A2(new_n434_), .ZN(new_n446_));
  NAND3_X1  g245(.A1(new_n412_), .A2(new_n421_), .A3(new_n429_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n446_), .B1(new_n447_), .B2(new_n434_), .ZN(new_n448_));
  AOI21_X1  g247(.A(new_n445_), .B1(new_n448_), .B2(new_n440_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n434_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n446_), .ZN(new_n451_));
  NAND2_X1  g250(.A1(new_n450_), .A2(new_n451_), .ZN(new_n452_));
  NAND2_X1  g251(.A1(new_n452_), .A2(new_n441_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n448_), .A2(new_n440_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(new_n454_), .ZN(new_n455_));
  AOI22_X1  g254(.A1(new_n444_), .A2(new_n449_), .B1(new_n455_), .B2(new_n445_), .ZN(new_n456_));
  INV_X1    g255(.A(KEYINPUT91), .ZN(new_n457_));
  XNOR2_X1  g256(.A(G155gat), .B(G162gat), .ZN(new_n458_));
  OR2_X1    g257(.A1(G141gat), .A2(G148gat), .ZN(new_n459_));
  NAND2_X1  g258(.A1(new_n459_), .A2(KEYINPUT3), .ZN(new_n460_));
  OR3_X1    g259(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n461_));
  NAND2_X1  g260(.A1(G141gat), .A2(G148gat), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT2), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n462_), .A2(new_n463_), .ZN(new_n464_));
  AND3_X1   g263(.A1(new_n460_), .A2(new_n461_), .A3(new_n464_), .ZN(new_n465_));
  NAND3_X1  g264(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(new_n466_), .B(KEYINPUT90), .ZN(new_n467_));
  AOI21_X1  g266(.A(new_n458_), .B1(new_n465_), .B2(new_n467_), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n458_), .A2(KEYINPUT1), .ZN(new_n469_));
  NAND3_X1  g268(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n470_));
  NAND3_X1  g269(.A1(new_n459_), .A2(new_n470_), .A3(new_n462_), .ZN(new_n471_));
  NOR2_X1   g270(.A1(new_n469_), .A2(new_n471_), .ZN(new_n472_));
  OR2_X1    g271(.A1(new_n468_), .A2(new_n472_), .ZN(new_n473_));
  OAI21_X1  g272(.A(KEYINPUT28), .B1(new_n473_), .B2(KEYINPUT29), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n468_), .A2(new_n472_), .ZN(new_n475_));
  INV_X1    g274(.A(KEYINPUT28), .ZN(new_n476_));
  INV_X1    g275(.A(KEYINPUT29), .ZN(new_n477_));
  NAND3_X1  g276(.A1(new_n475_), .A2(new_n476_), .A3(new_n477_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G22gat), .B(G50gat), .ZN(new_n479_));
  NAND3_X1  g278(.A1(new_n474_), .A2(new_n478_), .A3(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(new_n480_), .ZN(new_n481_));
  AOI21_X1  g280(.A(new_n479_), .B1(new_n474_), .B2(new_n478_), .ZN(new_n482_));
  OAI21_X1  g281(.A(new_n457_), .B1(new_n481_), .B2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n482_), .ZN(new_n484_));
  NAND3_X1  g283(.A1(new_n484_), .A2(KEYINPUT91), .A3(new_n480_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n483_), .A2(new_n485_), .ZN(new_n486_));
  OAI21_X1  g285(.A(new_n410_), .B1(new_n475_), .B2(new_n477_), .ZN(new_n487_));
  INV_X1    g286(.A(G228gat), .ZN(new_n488_));
  INV_X1    g287(.A(G233gat), .ZN(new_n489_));
  NOR2_X1   g288(.A1(new_n488_), .A2(new_n489_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n487_), .A2(new_n490_), .ZN(new_n491_));
  OAI221_X1 g290(.A(new_n410_), .B1(new_n488_), .B2(new_n489_), .C1(new_n475_), .C2(new_n477_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n491_), .A2(new_n492_), .ZN(new_n493_));
  XNOR2_X1  g292(.A(G78gat), .B(G106gat), .ZN(new_n494_));
  XNOR2_X1  g293(.A(new_n493_), .B(new_n494_), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(KEYINPUT93), .ZN(new_n496_));
  NAND3_X1  g295(.A1(new_n491_), .A2(new_n492_), .A3(new_n496_), .ZN(new_n497_));
  AND3_X1   g296(.A1(new_n484_), .A2(new_n497_), .A3(new_n480_), .ZN(new_n498_));
  NAND3_X1  g297(.A1(new_n493_), .A2(KEYINPUT93), .A3(new_n494_), .ZN(new_n499_));
  AOI22_X1  g298(.A1(new_n486_), .A2(new_n495_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(G227gat), .A2(G233gat), .ZN(new_n501_));
  XNOR2_X1  g300(.A(new_n501_), .B(new_n301_), .ZN(new_n502_));
  XNOR2_X1  g301(.A(new_n502_), .B(KEYINPUT30), .ZN(new_n503_));
  XNOR2_X1  g302(.A(new_n503_), .B(KEYINPUT31), .ZN(new_n504_));
  INV_X1    g303(.A(new_n504_), .ZN(new_n505_));
  XOR2_X1   g304(.A(G71gat), .B(G99gat), .Z(new_n506_));
  XOR2_X1   g305(.A(KEYINPUT88), .B(G43gat), .Z(new_n507_));
  XOR2_X1   g306(.A(new_n506_), .B(new_n507_), .Z(new_n508_));
  INV_X1    g307(.A(new_n508_), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n396_), .A2(new_n509_), .ZN(new_n510_));
  XNOR2_X1  g309(.A(G127gat), .B(G134gat), .ZN(new_n511_));
  INV_X1    g310(.A(KEYINPUT89), .ZN(new_n512_));
  XNOR2_X1  g311(.A(new_n511_), .B(new_n512_), .ZN(new_n513_));
  XNOR2_X1  g312(.A(G113gat), .B(G120gat), .ZN(new_n514_));
  NAND2_X1  g313(.A1(new_n513_), .A2(new_n514_), .ZN(new_n515_));
  XNOR2_X1  g314(.A(new_n511_), .B(KEYINPUT89), .ZN(new_n516_));
  INV_X1    g315(.A(new_n514_), .ZN(new_n517_));
  NAND2_X1  g316(.A1(new_n516_), .A2(new_n517_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n515_), .A2(new_n518_), .ZN(new_n519_));
  OAI21_X1  g318(.A(new_n508_), .B1(new_n383_), .B2(new_n395_), .ZN(new_n520_));
  NAND3_X1  g319(.A1(new_n510_), .A2(new_n519_), .A3(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(new_n521_), .ZN(new_n522_));
  AOI21_X1  g321(.A(new_n519_), .B1(new_n510_), .B2(new_n520_), .ZN(new_n523_));
  OAI21_X1  g322(.A(new_n505_), .B1(new_n522_), .B2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n523_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n525_), .A2(new_n504_), .A3(new_n521_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n526_), .ZN(new_n527_));
  INV_X1    g326(.A(new_n527_), .ZN(new_n528_));
  NAND2_X1  g327(.A1(new_n519_), .A2(new_n475_), .ZN(new_n529_));
  OAI211_X1 g328(.A(new_n515_), .B(new_n518_), .C1(new_n468_), .C2(new_n472_), .ZN(new_n530_));
  NAND3_X1  g329(.A1(new_n529_), .A2(KEYINPUT4), .A3(new_n530_), .ZN(new_n531_));
  NAND2_X1  g330(.A1(G225gat), .A2(G233gat), .ZN(new_n532_));
  INV_X1    g331(.A(new_n532_), .ZN(new_n533_));
  INV_X1    g332(.A(new_n519_), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT4), .ZN(new_n535_));
  NAND3_X1  g334(.A1(new_n534_), .A2(new_n535_), .A3(new_n473_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n531_), .A2(new_n533_), .A3(new_n536_), .ZN(new_n537_));
  NAND3_X1  g336(.A1(new_n529_), .A2(new_n530_), .A3(new_n532_), .ZN(new_n538_));
  NAND2_X1  g337(.A1(new_n537_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G1gat), .B(G29gat), .ZN(new_n540_));
  XNOR2_X1  g339(.A(new_n540_), .B(G85gat), .ZN(new_n541_));
  XNOR2_X1  g340(.A(KEYINPUT0), .B(G57gat), .ZN(new_n542_));
  XNOR2_X1  g341(.A(new_n541_), .B(new_n542_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n539_), .A2(new_n543_), .ZN(new_n544_));
  INV_X1    g343(.A(new_n543_), .ZN(new_n545_));
  NAND3_X1  g344(.A1(new_n537_), .A2(new_n538_), .A3(new_n545_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n544_), .A2(new_n546_), .ZN(new_n547_));
  NOR2_X1   g346(.A1(new_n528_), .A2(new_n547_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n456_), .A2(KEYINPUT100), .A3(new_n500_), .A4(new_n548_), .ZN(new_n549_));
  NAND2_X1  g348(.A1(new_n455_), .A2(new_n445_), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n449_), .B1(new_n442_), .B2(new_n443_), .ZN(new_n551_));
  NAND4_X1  g350(.A1(new_n550_), .A2(new_n548_), .A3(new_n551_), .A4(new_n500_), .ZN(new_n552_));
  INV_X1    g351(.A(KEYINPUT100), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(new_n549_), .A2(new_n554_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT98), .ZN(new_n556_));
  INV_X1    g355(.A(KEYINPUT97), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n440_), .A2(KEYINPUT32), .ZN(new_n558_));
  INV_X1    g357(.A(new_n558_), .ZN(new_n559_));
  AOI21_X1  g358(.A(new_n557_), .B1(new_n436_), .B2(new_n559_), .ZN(new_n560_));
  AOI211_X1 g359(.A(KEYINPUT97), .B(new_n558_), .C1(new_n430_), .C2(new_n435_), .ZN(new_n561_));
  NOR2_X1   g360(.A1(new_n560_), .A2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n448_), .A2(new_n558_), .ZN(new_n563_));
  NAND2_X1  g362(.A1(new_n547_), .A2(new_n563_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n556_), .B1(new_n562_), .B2(new_n564_), .ZN(new_n565_));
  AOI22_X1  g364(.A1(new_n544_), .A2(new_n546_), .B1(new_n448_), .B2(new_n558_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n566_), .B(KEYINPUT98), .C1(new_n560_), .C2(new_n561_), .ZN(new_n567_));
  AND3_X1   g366(.A1(new_n531_), .A2(new_n532_), .A3(new_n536_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n529_), .A2(new_n530_), .A3(new_n533_), .ZN(new_n569_));
  AND2_X1   g368(.A1(new_n569_), .A2(new_n543_), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n568_), .B1(KEYINPUT96), .B2(new_n570_), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n570_), .A2(KEYINPUT96), .ZN(new_n572_));
  INV_X1    g371(.A(KEYINPUT33), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n571_), .A2(new_n572_), .B1(new_n573_), .B2(new_n546_), .ZN(new_n574_));
  OR2_X1    g373(.A1(new_n546_), .A2(new_n573_), .ZN(new_n575_));
  NAND4_X1  g374(.A1(new_n574_), .A2(new_n454_), .A3(new_n453_), .A4(new_n575_), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n565_), .A2(new_n567_), .A3(new_n576_), .ZN(new_n577_));
  NOR2_X1   g376(.A1(new_n500_), .A2(new_n547_), .ZN(new_n578_));
  AOI22_X1  g377(.A1(new_n577_), .A2(new_n500_), .B1(new_n578_), .B2(new_n456_), .ZN(new_n579_));
  OAI21_X1  g378(.A(new_n555_), .B1(new_n579_), .B2(new_n527_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n245_), .ZN(new_n581_));
  OR2_X1    g380(.A1(new_n581_), .A2(new_n307_), .ZN(new_n582_));
  NAND2_X1  g381(.A1(G229gat), .A2(G233gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n583_), .B(KEYINPUT84), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT82), .ZN(new_n585_));
  XNOR2_X1  g384(.A(new_n244_), .B(new_n585_), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n586_), .A2(new_n307_), .A3(KEYINPUT83), .ZN(new_n587_));
  INV_X1    g386(.A(new_n587_), .ZN(new_n588_));
  AOI21_X1  g387(.A(KEYINPUT83), .B1(new_n586_), .B2(new_n307_), .ZN(new_n589_));
  OAI211_X1 g388(.A(new_n582_), .B(new_n584_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n590_));
  NOR2_X1   g389(.A1(new_n586_), .A2(new_n307_), .ZN(new_n591_));
  INV_X1    g390(.A(new_n589_), .ZN(new_n592_));
  AOI21_X1  g391(.A(new_n591_), .B1(new_n592_), .B2(new_n587_), .ZN(new_n593_));
  OAI21_X1  g392(.A(new_n590_), .B1(new_n593_), .B2(new_n583_), .ZN(new_n594_));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G169gat), .B(G197gat), .ZN(new_n596_));
  XOR2_X1   g395(.A(new_n595_), .B(new_n596_), .Z(new_n597_));
  INV_X1    g396(.A(new_n597_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n598_), .A2(KEYINPUT85), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n594_), .B(new_n599_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n580_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(new_n367_), .A2(new_n602_), .ZN(new_n603_));
  OR2_X1    g402(.A1(new_n547_), .A2(KEYINPUT101), .ZN(new_n604_));
  NAND2_X1  g403(.A1(new_n547_), .A2(KEYINPUT101), .ZN(new_n605_));
  NAND2_X1  g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  INV_X1    g405(.A(new_n606_), .ZN(new_n607_));
  NOR3_X1   g406(.A1(new_n603_), .A2(G1gat), .A3(new_n607_), .ZN(new_n608_));
  NAND3_X1  g407(.A1(new_n365_), .A2(new_n601_), .A3(new_n324_), .ZN(new_n609_));
  INV_X1    g408(.A(KEYINPUT102), .ZN(new_n610_));
  OR2_X1    g409(.A1(new_n609_), .A2(new_n610_), .ZN(new_n611_));
  AND2_X1   g410(.A1(new_n287_), .A2(new_n289_), .ZN(new_n612_));
  INV_X1    g411(.A(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n580_), .A2(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n609_), .A2(new_n610_), .ZN(new_n615_));
  AND3_X1   g414(.A1(new_n611_), .A2(new_n614_), .A3(new_n615_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(new_n547_), .ZN(new_n617_));
  AOI22_X1  g416(.A1(new_n608_), .A2(KEYINPUT38), .B1(new_n617_), .B2(G1gat), .ZN(new_n618_));
  INV_X1    g417(.A(KEYINPUT103), .ZN(new_n619_));
  OR3_X1    g418(.A1(new_n603_), .A2(G1gat), .A3(new_n607_), .ZN(new_n620_));
  INV_X1    g419(.A(KEYINPUT38), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n619_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  NOR3_X1   g421(.A1(new_n608_), .A2(KEYINPUT103), .A3(KEYINPUT38), .ZN(new_n623_));
  OAI21_X1  g422(.A(new_n618_), .B1(new_n622_), .B2(new_n623_), .ZN(new_n624_));
  INV_X1    g423(.A(KEYINPUT104), .ZN(new_n625_));
  XNOR2_X1  g424(.A(new_n624_), .B(new_n625_), .ZN(G1324gat));
  INV_X1    g425(.A(new_n603_), .ZN(new_n627_));
  INV_X1    g426(.A(G8gat), .ZN(new_n628_));
  INV_X1    g427(.A(new_n456_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n627_), .A2(new_n628_), .A3(new_n629_), .ZN(new_n630_));
  INV_X1    g429(.A(KEYINPUT105), .ZN(new_n631_));
  NAND2_X1  g430(.A1(new_n616_), .A2(new_n629_), .ZN(new_n632_));
  INV_X1    g431(.A(KEYINPUT39), .ZN(new_n633_));
  AND4_X1   g432(.A1(new_n631_), .A2(new_n632_), .A3(new_n633_), .A4(G8gat), .ZN(new_n634_));
  AOI21_X1  g433(.A(new_n628_), .B1(KEYINPUT105), .B2(KEYINPUT39), .ZN(new_n635_));
  AOI22_X1  g434(.A1(new_n632_), .A2(new_n635_), .B1(new_n631_), .B2(new_n633_), .ZN(new_n636_));
  OAI21_X1  g435(.A(new_n630_), .B1(new_n634_), .B2(new_n636_), .ZN(new_n637_));
  XNOR2_X1  g436(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n638_));
  XOR2_X1   g437(.A(new_n637_), .B(new_n638_), .Z(G1325gat));
  AOI21_X1  g438(.A(new_n301_), .B1(new_n616_), .B2(new_n527_), .ZN(new_n640_));
  XNOR2_X1  g439(.A(new_n640_), .B(KEYINPUT41), .ZN(new_n641_));
  NAND3_X1  g440(.A1(new_n627_), .A2(new_n301_), .A3(new_n527_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1326gat));
  INV_X1    g442(.A(new_n500_), .ZN(new_n644_));
  AOI21_X1  g443(.A(new_n302_), .B1(new_n616_), .B2(new_n644_), .ZN(new_n645_));
  XOR2_X1   g444(.A(new_n645_), .B(KEYINPUT42), .Z(new_n646_));
  NAND3_X1  g445(.A1(new_n627_), .A2(new_n302_), .A3(new_n644_), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(new_n647_), .ZN(G1327gat));
  INV_X1    g447(.A(new_n365_), .ZN(new_n649_));
  INV_X1    g448(.A(new_n324_), .ZN(new_n650_));
  NAND2_X1  g449(.A1(new_n650_), .A2(new_n612_), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n649_), .A2(new_n651_), .ZN(new_n652_));
  AND2_X1   g451(.A1(new_n602_), .A2(new_n652_), .ZN(new_n653_));
  AOI21_X1  g452(.A(G29gat), .B1(new_n653_), .B2(new_n547_), .ZN(new_n654_));
  INV_X1    g453(.A(KEYINPUT44), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n365_), .A2(new_n601_), .A3(new_n650_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n291_), .A2(new_n292_), .ZN(new_n657_));
  NAND2_X1  g456(.A1(new_n580_), .A2(new_n657_), .ZN(new_n658_));
  NAND2_X1  g457(.A1(new_n658_), .A2(KEYINPUT43), .ZN(new_n659_));
  INV_X1    g458(.A(KEYINPUT43), .ZN(new_n660_));
  NAND3_X1  g459(.A1(new_n580_), .A2(new_n657_), .A3(new_n660_), .ZN(new_n661_));
  AOI21_X1  g460(.A(new_n656_), .B1(new_n659_), .B2(new_n661_), .ZN(new_n662_));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n655_), .B1(new_n662_), .B2(new_n663_), .ZN(new_n664_));
  AOI211_X1 g463(.A(KEYINPUT107), .B(new_n656_), .C1(new_n659_), .C2(new_n661_), .ZN(new_n665_));
  NOR2_X1   g464(.A1(new_n664_), .A2(new_n665_), .ZN(new_n666_));
  AOI21_X1  g465(.A(new_n666_), .B1(KEYINPUT44), .B2(new_n662_), .ZN(new_n667_));
  AND2_X1   g466(.A1(new_n606_), .A2(G29gat), .ZN(new_n668_));
  AOI21_X1  g467(.A(new_n654_), .B1(new_n667_), .B2(new_n668_), .ZN(G1328gat));
  OR2_X1    g468(.A1(new_n456_), .A2(KEYINPUT108), .ZN(new_n670_));
  NAND2_X1  g469(.A1(new_n456_), .A2(KEYINPUT108), .ZN(new_n671_));
  NAND2_X1  g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  INV_X1    g471(.A(new_n672_), .ZN(new_n673_));
  NOR2_X1   g472(.A1(new_n673_), .A2(G36gat), .ZN(new_n674_));
  NAND3_X1  g473(.A1(new_n602_), .A2(new_n652_), .A3(new_n674_), .ZN(new_n675_));
  XNOR2_X1  g474(.A(new_n675_), .B(KEYINPUT45), .ZN(new_n676_));
  INV_X1    g475(.A(KEYINPUT109), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n676_), .B1(new_n677_), .B2(KEYINPUT46), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n662_), .A2(KEYINPUT44), .ZN(new_n679_));
  OAI211_X1 g478(.A(new_n629_), .B(new_n679_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n680_));
  AOI21_X1  g479(.A(new_n678_), .B1(G36gat), .B2(new_n680_), .ZN(new_n681_));
  AND2_X1   g480(.A1(new_n677_), .A2(KEYINPUT46), .ZN(new_n682_));
  XNOR2_X1  g481(.A(new_n681_), .B(new_n682_), .ZN(G1329gat));
  AOI21_X1  g482(.A(G43gat), .B1(new_n653_), .B2(new_n527_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n527_), .A2(G43gat), .ZN(new_n685_));
  AOI21_X1  g484(.A(new_n685_), .B1(new_n662_), .B2(KEYINPUT44), .ZN(new_n686_));
  OAI21_X1  g485(.A(new_n686_), .B1(new_n664_), .B2(new_n665_), .ZN(new_n687_));
  INV_X1    g486(.A(KEYINPUT110), .ZN(new_n688_));
  NAND2_X1  g487(.A1(new_n687_), .A2(new_n688_), .ZN(new_n689_));
  OAI211_X1 g488(.A(KEYINPUT110), .B(new_n686_), .C1(new_n664_), .C2(new_n665_), .ZN(new_n690_));
  AOI21_X1  g489(.A(new_n684_), .B1(new_n689_), .B2(new_n690_), .ZN(new_n691_));
  XNOR2_X1  g490(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n691_), .B(new_n693_), .ZN(G1330gat));
  NAND2_X1  g493(.A1(new_n667_), .A2(new_n644_), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n695_), .A2(G50gat), .ZN(new_n696_));
  NOR2_X1   g495(.A1(new_n500_), .A2(G50gat), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT112), .ZN(new_n698_));
  NAND2_X1  g497(.A1(new_n653_), .A2(new_n698_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n696_), .A2(new_n699_), .ZN(G1331gat));
  NAND4_X1  g499(.A1(new_n614_), .A2(new_n600_), .A3(new_n324_), .A4(new_n649_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n701_), .B(KEYINPUT114), .ZN(new_n702_));
  INV_X1    g501(.A(new_n547_), .ZN(new_n703_));
  OAI21_X1  g502(.A(G57gat), .B1(new_n702_), .B2(new_n703_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n580_), .A2(new_n600_), .ZN(new_n705_));
  XOR2_X1   g504(.A(new_n705_), .B(KEYINPUT113), .Z(new_n706_));
  NOR3_X1   g505(.A1(new_n657_), .A2(new_n650_), .A3(new_n365_), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OR2_X1    g507(.A1(new_n607_), .A2(G57gat), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n704_), .B1(new_n708_), .B2(new_n709_), .ZN(G1332gat));
  OAI21_X1  g509(.A(G64gat), .B1(new_n702_), .B2(new_n673_), .ZN(new_n711_));
  XOR2_X1   g510(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n712_));
  XNOR2_X1  g511(.A(new_n711_), .B(new_n712_), .ZN(new_n713_));
  OR3_X1    g512(.A1(new_n708_), .A2(G64gat), .A3(new_n673_), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n713_), .A2(new_n714_), .ZN(G1333gat));
  OR3_X1    g514(.A1(new_n708_), .A2(G71gat), .A3(new_n528_), .ZN(new_n716_));
  OAI21_X1  g515(.A(G71gat), .B1(new_n702_), .B2(new_n528_), .ZN(new_n717_));
  AND2_X1   g516(.A1(new_n717_), .A2(KEYINPUT49), .ZN(new_n718_));
  NOR2_X1   g517(.A1(new_n717_), .A2(KEYINPUT49), .ZN(new_n719_));
  OAI21_X1  g518(.A(new_n716_), .B1(new_n718_), .B2(new_n719_), .ZN(G1334gat));
  OAI21_X1  g519(.A(G78gat), .B1(new_n702_), .B2(new_n500_), .ZN(new_n721_));
  XNOR2_X1  g520(.A(new_n721_), .B(KEYINPUT50), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n644_), .A2(new_n312_), .ZN(new_n723_));
  OAI21_X1  g522(.A(new_n722_), .B1(new_n708_), .B2(new_n723_), .ZN(G1335gat));
  NOR2_X1   g523(.A1(new_n651_), .A2(new_n365_), .ZN(new_n725_));
  NAND2_X1  g524(.A1(new_n706_), .A2(new_n725_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n726_), .A2(KEYINPUT116), .ZN(new_n727_));
  INV_X1    g526(.A(KEYINPUT116), .ZN(new_n728_));
  NAND3_X1  g527(.A1(new_n706_), .A2(new_n728_), .A3(new_n725_), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n727_), .A2(new_n729_), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n730_), .A2(new_n215_), .A3(new_n606_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n659_), .A2(new_n661_), .ZN(new_n732_));
  NAND4_X1  g531(.A1(new_n650_), .A2(new_n362_), .A3(new_n600_), .A4(new_n364_), .ZN(new_n733_));
  XNOR2_X1  g532(.A(new_n733_), .B(KEYINPUT117), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(new_n735_));
  AND2_X1   g534(.A1(new_n735_), .A2(KEYINPUT118), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n735_), .A2(KEYINPUT118), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  OAI21_X1  g537(.A(G85gat), .B1(new_n738_), .B2(new_n703_), .ZN(new_n739_));
  NAND2_X1  g538(.A1(new_n731_), .A2(new_n739_), .ZN(G1336gat));
  NAND3_X1  g539(.A1(new_n730_), .A2(new_n216_), .A3(new_n629_), .ZN(new_n741_));
  OAI21_X1  g540(.A(G92gat), .B1(new_n738_), .B2(new_n673_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n741_), .A2(new_n742_), .ZN(G1337gat));
  OAI21_X1  g542(.A(G99gat), .B1(new_n738_), .B2(new_n528_), .ZN(new_n744_));
  AND2_X1   g543(.A1(new_n205_), .A2(new_n208_), .ZN(new_n745_));
  NOR2_X1   g544(.A1(new_n528_), .A2(new_n745_), .ZN(new_n746_));
  NAND2_X1  g545(.A1(new_n730_), .A2(new_n746_), .ZN(new_n747_));
  NAND4_X1  g546(.A1(new_n744_), .A2(new_n747_), .A3(KEYINPUT119), .A4(KEYINPUT51), .ZN(new_n748_));
  OR2_X1    g547(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n749_));
  NAND2_X1  g548(.A1(KEYINPUT119), .A2(KEYINPUT51), .ZN(new_n750_));
  XNOR2_X1  g549(.A(new_n735_), .B(KEYINPUT118), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n226_), .B1(new_n751_), .B2(new_n527_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n746_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n753_), .B1(new_n727_), .B2(new_n729_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n749_), .B(new_n750_), .C1(new_n752_), .C2(new_n754_), .ZN(new_n755_));
  AND2_X1   g554(.A1(new_n748_), .A2(new_n755_), .ZN(G1338gat));
  NOR2_X1   g555(.A1(new_n500_), .A2(G106gat), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n730_), .A2(new_n757_), .ZN(new_n758_));
  OAI21_X1  g557(.A(G106gat), .B1(new_n735_), .B2(new_n500_), .ZN(new_n759_));
  NOR2_X1   g558(.A1(new_n759_), .A2(KEYINPUT52), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n759_), .A2(KEYINPUT52), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n758_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  NAND2_X1  g561(.A1(new_n762_), .A2(KEYINPUT53), .ZN(new_n763_));
  INV_X1    g562(.A(KEYINPUT53), .ZN(new_n764_));
  OAI211_X1 g563(.A(new_n758_), .B(new_n764_), .C1(new_n761_), .C2(new_n760_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n763_), .A2(new_n765_), .ZN(G1339gat));
  INV_X1    g565(.A(new_n584_), .ZN(new_n767_));
  OAI211_X1 g566(.A(new_n582_), .B(new_n767_), .C1(new_n588_), .C2(new_n589_), .ZN(new_n768_));
  OAI21_X1  g567(.A(new_n768_), .B1(new_n593_), .B2(new_n767_), .ZN(new_n769_));
  MUX2_X1   g568(.A(new_n769_), .B(new_n594_), .S(new_n597_), .Z(new_n770_));
  INV_X1    g569(.A(KEYINPUT121), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n770_), .A2(new_n359_), .A3(new_n771_), .ZN(new_n772_));
  AOI21_X1  g571(.A(new_n771_), .B1(new_n770_), .B2(new_n359_), .ZN(new_n773_));
  NOR2_X1   g572(.A1(new_n772_), .A2(new_n773_), .ZN(new_n774_));
  INV_X1    g573(.A(KEYINPUT55), .ZN(new_n775_));
  AND3_X1   g574(.A1(new_n339_), .A2(KEYINPUT72), .A3(new_n340_), .ZN(new_n776_));
  AOI21_X1  g575(.A(KEYINPUT72), .B1(new_n339_), .B2(new_n340_), .ZN(new_n777_));
  NOR2_X1   g576(.A1(new_n776_), .A2(new_n777_), .ZN(new_n778_));
  NAND3_X1  g577(.A1(new_n331_), .A2(new_n335_), .A3(new_n337_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n775_), .B1(new_n778_), .B2(new_n779_), .ZN(new_n780_));
  NAND3_X1  g579(.A1(new_n338_), .A2(new_n345_), .A3(KEYINPUT55), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n347_), .B1(new_n349_), .B2(new_n779_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n780_), .A2(new_n781_), .A3(new_n782_), .ZN(new_n783_));
  NAND3_X1  g582(.A1(new_n783_), .A2(KEYINPUT56), .A3(new_n356_), .ZN(new_n784_));
  INV_X1    g583(.A(KEYINPUT122), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n784_), .A2(new_n785_), .ZN(new_n786_));
  NAND2_X1  g585(.A1(new_n783_), .A2(new_n356_), .ZN(new_n787_));
  INV_X1    g586(.A(KEYINPUT56), .ZN(new_n788_));
  NAND2_X1  g587(.A1(new_n787_), .A2(new_n788_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n786_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n787_), .A2(new_n785_), .A3(new_n788_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n774_), .B1(new_n790_), .B2(new_n791_), .ZN(new_n792_));
  OAI21_X1  g591(.A(new_n657_), .B1(new_n792_), .B2(KEYINPUT58), .ZN(new_n793_));
  INV_X1    g592(.A(KEYINPUT58), .ZN(new_n794_));
  AOI211_X1 g593(.A(new_n794_), .B(new_n774_), .C1(new_n790_), .C2(new_n791_), .ZN(new_n795_));
  AND2_X1   g594(.A1(new_n601_), .A2(new_n359_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT56), .B1(new_n783_), .B2(new_n356_), .ZN(new_n797_));
  OAI21_X1  g596(.A(new_n784_), .B1(new_n797_), .B2(KEYINPUT120), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT120), .ZN(new_n799_));
  AOI211_X1 g598(.A(new_n799_), .B(KEYINPUT56), .C1(new_n783_), .C2(new_n356_), .ZN(new_n800_));
  OAI21_X1  g599(.A(new_n796_), .B1(new_n798_), .B2(new_n800_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n360_), .A2(new_n770_), .ZN(new_n802_));
  AOI21_X1  g601(.A(new_n612_), .B1(new_n801_), .B2(new_n802_), .ZN(new_n803_));
  OAI22_X1  g602(.A1(new_n793_), .A2(new_n795_), .B1(new_n803_), .B2(KEYINPUT57), .ZN(new_n804_));
  AND2_X1   g603(.A1(new_n803_), .A2(KEYINPUT57), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  OAI21_X1  g605(.A(KEYINPUT54), .B1(new_n366_), .B2(new_n601_), .ZN(new_n807_));
  OR3_X1    g606(.A1(new_n366_), .A2(KEYINPUT54), .A3(new_n601_), .ZN(new_n808_));
  AOI22_X1  g607(.A1(new_n806_), .A2(new_n650_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  NOR2_X1   g608(.A1(new_n629_), .A2(new_n644_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n607_), .A2(new_n528_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n810_), .A2(new_n811_), .ZN(new_n812_));
  OAI21_X1  g611(.A(KEYINPUT59), .B1(new_n809_), .B2(new_n812_), .ZN(new_n813_));
  INV_X1    g612(.A(KEYINPUT123), .ZN(new_n814_));
  AOI21_X1  g613(.A(new_n805_), .B1(new_n804_), .B2(new_n814_), .ZN(new_n815_));
  OAI221_X1 g614(.A(KEYINPUT123), .B1(new_n803_), .B2(KEYINPUT57), .C1(new_n795_), .C2(new_n793_), .ZN(new_n816_));
  AOI21_X1  g615(.A(new_n324_), .B1(new_n815_), .B2(new_n816_), .ZN(new_n817_));
  AND2_X1   g616(.A1(new_n808_), .A2(new_n807_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OR2_X1    g618(.A1(new_n812_), .A2(KEYINPUT59), .ZN(new_n820_));
  OAI21_X1  g619(.A(new_n813_), .B1(new_n819_), .B2(new_n820_), .ZN(new_n821_));
  OAI21_X1  g620(.A(G113gat), .B1(new_n821_), .B2(new_n600_), .ZN(new_n822_));
  NOR2_X1   g621(.A1(new_n809_), .A2(new_n812_), .ZN(new_n823_));
  INV_X1    g622(.A(G113gat), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n601_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n822_), .A2(new_n825_), .ZN(G1340gat));
  NAND2_X1  g625(.A1(new_n806_), .A2(new_n650_), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n808_), .A2(new_n807_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n827_), .A2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n812_), .ZN(new_n830_));
  NOR2_X1   g629(.A1(new_n365_), .A2(KEYINPUT60), .ZN(new_n831_));
  MUX2_X1   g630(.A(new_n831_), .B(KEYINPUT60), .S(G120gat), .Z(new_n832_));
  NAND3_X1  g631(.A1(new_n829_), .A2(new_n830_), .A3(new_n832_), .ZN(new_n833_));
  XNOR2_X1  g632(.A(new_n833_), .B(KEYINPUT124), .ZN(new_n834_));
  OAI211_X1 g633(.A(new_n813_), .B(new_n649_), .C1(new_n819_), .C2(new_n820_), .ZN(new_n835_));
  NAND2_X1  g634(.A1(new_n835_), .A2(G120gat), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n834_), .A2(new_n836_), .ZN(G1341gat));
  OAI21_X1  g636(.A(G127gat), .B1(new_n821_), .B2(new_n650_), .ZN(new_n838_));
  INV_X1    g637(.A(G127gat), .ZN(new_n839_));
  NAND3_X1  g638(.A1(new_n823_), .A2(new_n839_), .A3(new_n324_), .ZN(new_n840_));
  NAND2_X1  g639(.A1(new_n838_), .A2(new_n840_), .ZN(G1342gat));
  OAI21_X1  g640(.A(G134gat), .B1(new_n821_), .B2(new_n293_), .ZN(new_n842_));
  INV_X1    g641(.A(G134gat), .ZN(new_n843_));
  NAND3_X1  g642(.A1(new_n823_), .A2(new_n843_), .A3(new_n612_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n842_), .A2(new_n844_), .ZN(G1343gat));
  NOR2_X1   g644(.A1(new_n809_), .A2(new_n527_), .ZN(new_n846_));
  NOR3_X1   g645(.A1(new_n672_), .A2(new_n500_), .A3(new_n607_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n846_), .A2(new_n601_), .A3(new_n847_), .ZN(new_n848_));
  XNOR2_X1  g647(.A(KEYINPUT125), .B(G141gat), .ZN(new_n849_));
  XNOR2_X1  g648(.A(new_n848_), .B(new_n849_), .ZN(G1344gat));
  NAND3_X1  g649(.A1(new_n846_), .A2(new_n649_), .A3(new_n847_), .ZN(new_n851_));
  XNOR2_X1  g650(.A(KEYINPUT126), .B(G148gat), .ZN(new_n852_));
  XNOR2_X1  g651(.A(new_n851_), .B(new_n852_), .ZN(G1345gat));
  NAND3_X1  g652(.A1(new_n846_), .A2(new_n324_), .A3(new_n847_), .ZN(new_n854_));
  XNOR2_X1  g653(.A(KEYINPUT61), .B(G155gat), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n854_), .B(new_n855_), .ZN(G1346gat));
  NAND2_X1  g655(.A1(new_n846_), .A2(new_n847_), .ZN(new_n857_));
  OAI21_X1  g656(.A(G162gat), .B1(new_n857_), .B2(new_n293_), .ZN(new_n858_));
  OR2_X1    g657(.A1(new_n613_), .A2(G162gat), .ZN(new_n859_));
  OAI21_X1  g658(.A(new_n858_), .B1(new_n857_), .B2(new_n859_), .ZN(G1347gat));
  NAND3_X1  g659(.A1(new_n672_), .A2(new_n527_), .A3(new_n607_), .ZN(new_n861_));
  NOR3_X1   g660(.A1(new_n819_), .A2(new_n644_), .A3(new_n861_), .ZN(new_n862_));
  NAND3_X1  g661(.A1(new_n862_), .A2(new_n601_), .A3(new_n417_), .ZN(new_n863_));
  NOR2_X1   g662(.A1(new_n861_), .A2(new_n644_), .ZN(new_n864_));
  OAI211_X1 g663(.A(new_n601_), .B(new_n864_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(G169gat), .ZN(new_n866_));
  INV_X1    g665(.A(KEYINPUT62), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n865_), .A2(KEYINPUT62), .A3(G169gat), .ZN(new_n869_));
  NAND3_X1  g668(.A1(new_n863_), .A2(new_n868_), .A3(new_n869_), .ZN(G1348gat));
  NAND2_X1  g669(.A1(new_n862_), .A2(new_n649_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n809_), .A2(new_n644_), .ZN(new_n872_));
  NOR3_X1   g671(.A1(new_n861_), .A2(new_n373_), .A3(new_n365_), .ZN(new_n873_));
  AOI22_X1  g672(.A1(new_n871_), .A2(new_n373_), .B1(new_n872_), .B2(new_n873_), .ZN(G1349gat));
  NOR2_X1   g673(.A1(new_n861_), .A2(new_n650_), .ZN(new_n875_));
  AOI21_X1  g674(.A(G183gat), .B1(new_n872_), .B2(new_n875_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n650_), .A2(new_n384_), .ZN(new_n877_));
  AOI21_X1  g676(.A(new_n876_), .B1(new_n862_), .B2(new_n877_), .ZN(G1350gat));
  OAI211_X1 g677(.A(new_n657_), .B(new_n864_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(G190gat), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n612_), .A2(new_n385_), .ZN(new_n881_));
  OAI211_X1 g680(.A(new_n864_), .B(new_n881_), .C1(new_n817_), .C2(new_n818_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n880_), .A2(new_n882_), .ZN(new_n883_));
  INV_X1    g682(.A(KEYINPUT127), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n883_), .A2(new_n884_), .ZN(new_n885_));
  NAND3_X1  g684(.A1(new_n880_), .A2(KEYINPUT127), .A3(new_n882_), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n885_), .A2(new_n886_), .ZN(G1351gat));
  AND2_X1   g686(.A1(new_n672_), .A2(new_n578_), .ZN(new_n888_));
  NAND3_X1  g687(.A1(new_n846_), .A2(new_n601_), .A3(new_n888_), .ZN(new_n889_));
  XNOR2_X1  g688(.A(new_n889_), .B(G197gat), .ZN(G1352gat));
  NAND3_X1  g689(.A1(new_n846_), .A2(new_n649_), .A3(new_n888_), .ZN(new_n891_));
  XNOR2_X1  g690(.A(new_n891_), .B(G204gat), .ZN(G1353gat));
  NAND4_X1  g691(.A1(new_n829_), .A2(new_n528_), .A3(new_n324_), .A4(new_n888_), .ZN(new_n893_));
  NOR2_X1   g692(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n894_));
  AND2_X1   g693(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n895_));
  NOR3_X1   g694(.A1(new_n893_), .A2(new_n894_), .A3(new_n895_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n896_), .B1(new_n893_), .B2(new_n894_), .ZN(G1354gat));
  NAND2_X1  g696(.A1(new_n846_), .A2(new_n888_), .ZN(new_n898_));
  OAI21_X1  g697(.A(G218gat), .B1(new_n898_), .B2(new_n293_), .ZN(new_n899_));
  OR2_X1    g698(.A1(new_n613_), .A2(G218gat), .ZN(new_n900_));
  OAI21_X1  g699(.A(new_n899_), .B1(new_n898_), .B2(new_n900_), .ZN(G1355gat));
endmodule


