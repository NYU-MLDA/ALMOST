//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 0 1 1 1 0 0 1 1 1 0 1 0 0 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:28:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n643_, new_n644_, new_n645_, new_n646_, new_n647_, new_n648_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n723_, new_n724_, new_n725_, new_n726_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n760_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n847_, new_n848_, new_n849_,
    new_n851_, new_n852_, new_n853_, new_n855_, new_n856_, new_n857_,
    new_n858_, new_n859_, new_n860_, new_n862_, new_n864_, new_n865_,
    new_n867_, new_n868_, new_n869_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n884_, new_n885_, new_n887_, new_n888_,
    new_n889_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n907_, new_n908_, new_n909_,
    new_n911_, new_n912_, new_n913_;
  INV_X1    g000(.A(KEYINPUT101), .ZN(new_n202_));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n203_), .B(KEYINPUT18), .ZN(new_n204_));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205_));
  XNOR2_X1  g004(.A(new_n204_), .B(new_n205_), .ZN(new_n206_));
  INV_X1    g005(.A(new_n206_), .ZN(new_n207_));
  AND2_X1   g006(.A1(new_n207_), .A2(KEYINPUT32), .ZN(new_n208_));
  AND2_X1   g007(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n209_));
  NOR2_X1   g008(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n210_));
  OAI21_X1  g009(.A(G197gat), .B1(new_n209_), .B2(new_n210_), .ZN(new_n211_));
  OAI21_X1  g010(.A(new_n211_), .B1(G197gat), .B2(G204gat), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT21), .ZN(new_n213_));
  XNOR2_X1  g012(.A(G211gat), .B(G218gat), .ZN(new_n214_));
  NOR3_X1   g013(.A1(new_n212_), .A2(new_n213_), .A3(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(new_n214_), .ZN(new_n217_));
  AOI21_X1  g016(.A(new_n217_), .B1(new_n212_), .B2(new_n213_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT91), .ZN(new_n219_));
  NOR3_X1   g018(.A1(new_n209_), .A2(new_n210_), .A3(G197gat), .ZN(new_n220_));
  INV_X1    g019(.A(G197gat), .ZN(new_n221_));
  INV_X1    g020(.A(G204gat), .ZN(new_n222_));
  OAI21_X1  g021(.A(KEYINPUT21), .B1(new_n221_), .B2(new_n222_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n219_), .B1(new_n220_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(KEYINPUT90), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n225_), .A2(new_n222_), .ZN(new_n226_));
  NAND2_X1  g025(.A1(KEYINPUT90), .A2(G204gat), .ZN(new_n227_));
  NAND3_X1  g026(.A1(new_n226_), .A2(new_n221_), .A3(new_n227_), .ZN(new_n228_));
  AOI21_X1  g027(.A(new_n213_), .B1(G197gat), .B2(G204gat), .ZN(new_n229_));
  NAND3_X1  g028(.A1(new_n228_), .A2(KEYINPUT91), .A3(new_n229_), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n224_), .A2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT92), .ZN(new_n232_));
  AND3_X1   g031(.A1(new_n218_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n233_));
  AOI21_X1  g032(.A(new_n232_), .B1(new_n218_), .B2(new_n231_), .ZN(new_n234_));
  OAI21_X1  g033(.A(new_n216_), .B1(new_n233_), .B2(new_n234_), .ZN(new_n235_));
  INV_X1    g034(.A(G169gat), .ZN(new_n236_));
  NAND2_X1  g035(.A1(new_n236_), .A2(KEYINPUT22), .ZN(new_n237_));
  INV_X1    g036(.A(KEYINPUT84), .ZN(new_n238_));
  AOI21_X1  g037(.A(G176gat), .B1(new_n237_), .B2(new_n238_), .ZN(new_n239_));
  XNOR2_X1  g038(.A(KEYINPUT22), .B(G169gat), .ZN(new_n240_));
  OAI21_X1  g039(.A(new_n239_), .B1(new_n238_), .B2(new_n240_), .ZN(new_n241_));
  NAND2_X1  g040(.A1(new_n241_), .A2(KEYINPUT85), .ZN(new_n242_));
  INV_X1    g041(.A(KEYINPUT85), .ZN(new_n243_));
  OAI211_X1 g042(.A(new_n239_), .B(new_n243_), .C1(new_n238_), .C2(new_n240_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n242_), .A2(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(G169gat), .A2(G176gat), .ZN(new_n246_));
  NAND2_X1  g045(.A1(new_n246_), .A2(KEYINPUT81), .ZN(new_n247_));
  INV_X1    g046(.A(KEYINPUT81), .ZN(new_n248_));
  NAND3_X1  g047(.A1(new_n248_), .A2(G169gat), .A3(G176gat), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n247_), .A2(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(G183gat), .A2(G190gat), .ZN(new_n251_));
  NAND2_X1  g050(.A1(new_n251_), .A2(KEYINPUT23), .ZN(new_n252_));
  INV_X1    g051(.A(KEYINPUT23), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n253_), .A2(G183gat), .A3(G190gat), .ZN(new_n254_));
  NAND3_X1  g053(.A1(new_n252_), .A2(new_n254_), .A3(KEYINPUT86), .ZN(new_n255_));
  INV_X1    g054(.A(KEYINPUT86), .ZN(new_n256_));
  NAND4_X1  g055(.A1(new_n256_), .A2(new_n253_), .A3(G183gat), .A4(G190gat), .ZN(new_n257_));
  AND2_X1   g056(.A1(new_n255_), .A2(new_n257_), .ZN(new_n258_));
  INV_X1    g057(.A(G183gat), .ZN(new_n259_));
  INV_X1    g058(.A(G190gat), .ZN(new_n260_));
  NAND2_X1  g059(.A1(new_n259_), .A2(new_n260_), .ZN(new_n261_));
  AOI21_X1  g060(.A(new_n250_), .B1(new_n258_), .B2(new_n261_), .ZN(new_n262_));
  XOR2_X1   g061(.A(new_n252_), .B(KEYINPUT82), .Z(new_n263_));
  XOR2_X1   g062(.A(new_n254_), .B(KEYINPUT83), .Z(new_n264_));
  NAND2_X1  g063(.A1(new_n263_), .A2(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(KEYINPUT25), .B(G183gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(KEYINPUT26), .B(G190gat), .ZN(new_n267_));
  INV_X1    g066(.A(KEYINPUT24), .ZN(new_n268_));
  NOR2_X1   g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269_));
  AOI22_X1  g068(.A1(new_n266_), .A2(new_n267_), .B1(new_n268_), .B2(new_n269_), .ZN(new_n270_));
  INV_X1    g069(.A(new_n269_), .ZN(new_n271_));
  NAND4_X1  g070(.A1(new_n271_), .A2(new_n247_), .A3(new_n249_), .A4(KEYINPUT24), .ZN(new_n272_));
  AND2_X1   g071(.A1(new_n270_), .A2(new_n272_), .ZN(new_n273_));
  AOI22_X1  g072(.A1(new_n245_), .A2(new_n262_), .B1(new_n265_), .B2(new_n273_), .ZN(new_n274_));
  INV_X1    g073(.A(new_n274_), .ZN(new_n275_));
  OAI211_X1 g074(.A(KEYINPUT95), .B(KEYINPUT20), .C1(new_n235_), .C2(new_n275_), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n252_), .B(KEYINPUT82), .ZN(new_n277_));
  XNOR2_X1  g076(.A(new_n254_), .B(KEYINPUT83), .ZN(new_n278_));
  OAI21_X1  g077(.A(new_n261_), .B1(new_n277_), .B2(new_n278_), .ZN(new_n279_));
  INV_X1    g078(.A(G176gat), .ZN(new_n280_));
  AOI21_X1  g079(.A(new_n250_), .B1(new_n280_), .B2(new_n240_), .ZN(new_n281_));
  NAND3_X1  g080(.A1(new_n271_), .A2(KEYINPUT24), .A3(new_n246_), .ZN(new_n282_));
  AND2_X1   g081(.A1(new_n270_), .A2(new_n282_), .ZN(new_n283_));
  AOI22_X1  g082(.A1(new_n279_), .A2(new_n281_), .B1(new_n283_), .B2(new_n258_), .ZN(new_n284_));
  AND3_X1   g083(.A1(new_n228_), .A2(KEYINPUT91), .A3(new_n229_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT91), .B1(new_n228_), .B2(new_n229_), .ZN(new_n286_));
  NOR2_X1   g085(.A1(new_n285_), .A2(new_n286_), .ZN(new_n287_));
  NOR2_X1   g086(.A1(G197gat), .A2(G204gat), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n226_), .A2(new_n227_), .ZN(new_n289_));
  AOI21_X1  g088(.A(new_n288_), .B1(new_n289_), .B2(G197gat), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n214_), .B1(new_n290_), .B2(KEYINPUT21), .ZN(new_n291_));
  OAI21_X1  g090(.A(KEYINPUT92), .B1(new_n287_), .B2(new_n291_), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n218_), .A2(new_n231_), .A3(new_n232_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n292_), .A2(new_n293_), .ZN(new_n294_));
  AOI21_X1  g093(.A(new_n284_), .B1(new_n294_), .B2(new_n216_), .ZN(new_n295_));
  INV_X1    g094(.A(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n276_), .A2(new_n296_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(G226gat), .A2(G233gat), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n298_), .B(KEYINPUT19), .ZN(new_n299_));
  NAND3_X1  g098(.A1(new_n294_), .A2(new_n274_), .A3(new_n216_), .ZN(new_n300_));
  AOI21_X1  g099(.A(KEYINPUT95), .B1(new_n300_), .B2(KEYINPUT20), .ZN(new_n301_));
  NOR3_X1   g100(.A1(new_n297_), .A2(new_n299_), .A3(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n299_), .ZN(new_n303_));
  INV_X1    g102(.A(KEYINPUT20), .ZN(new_n304_));
  AOI21_X1  g103(.A(new_n215_), .B1(new_n292_), .B2(new_n293_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n304_), .B1(new_n305_), .B2(new_n284_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n235_), .A2(new_n275_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n303_), .B1(new_n306_), .B2(new_n307_), .ZN(new_n308_));
  OAI21_X1  g107(.A(new_n208_), .B1(new_n302_), .B2(new_n308_), .ZN(new_n309_));
  OAI21_X1  g108(.A(new_n299_), .B1(new_n297_), .B2(new_n301_), .ZN(new_n310_));
  XOR2_X1   g109(.A(new_n208_), .B(KEYINPUT100), .Z(new_n311_));
  NAND2_X1  g110(.A1(new_n305_), .A2(new_n284_), .ZN(new_n312_));
  AND4_X1   g111(.A1(KEYINPUT20), .A2(new_n307_), .A3(new_n303_), .A4(new_n312_), .ZN(new_n313_));
  INV_X1    g112(.A(new_n313_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n310_), .A2(new_n311_), .A3(new_n314_), .ZN(new_n315_));
  XNOR2_X1  g114(.A(G127gat), .B(G134gat), .ZN(new_n316_));
  XNOR2_X1  g115(.A(G113gat), .B(G120gat), .ZN(new_n317_));
  XNOR2_X1  g116(.A(new_n316_), .B(new_n317_), .ZN(new_n318_));
  NOR2_X1   g117(.A1(G155gat), .A2(G162gat), .ZN(new_n319_));
  NAND2_X1  g118(.A1(G155gat), .A2(G162gat), .ZN(new_n320_));
  AOI21_X1  g119(.A(new_n319_), .B1(KEYINPUT1), .B2(new_n320_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n320_), .A2(KEYINPUT1), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(new_n322_), .ZN(new_n323_));
  NAND2_X1  g122(.A1(G141gat), .A2(G148gat), .ZN(new_n324_));
  INV_X1    g123(.A(new_n324_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(G141gat), .A2(G148gat), .ZN(new_n326_));
  NOR2_X1   g125(.A1(new_n325_), .A2(new_n326_), .ZN(new_n327_));
  NAND2_X1  g126(.A1(new_n323_), .A2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n329_));
  INV_X1    g128(.A(KEYINPUT89), .ZN(new_n330_));
  XNOR2_X1  g129(.A(new_n329_), .B(new_n330_), .ZN(new_n331_));
  NOR3_X1   g130(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n332_));
  AND3_X1   g131(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n333_));
  AOI21_X1  g132(.A(KEYINPUT2), .B1(G141gat), .B2(G148gat), .ZN(new_n334_));
  NOR3_X1   g133(.A1(new_n332_), .A2(new_n333_), .A3(new_n334_), .ZN(new_n335_));
  AND2_X1   g134(.A1(new_n331_), .A2(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n319_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n337_), .A2(new_n320_), .ZN(new_n338_));
  OAI211_X1 g137(.A(new_n318_), .B(new_n328_), .C1(new_n336_), .C2(new_n338_), .ZN(new_n339_));
  XOR2_X1   g138(.A(new_n316_), .B(new_n317_), .Z(new_n340_));
  AOI21_X1  g139(.A(new_n338_), .B1(new_n331_), .B2(new_n335_), .ZN(new_n341_));
  AND2_X1   g140(.A1(new_n323_), .A2(new_n327_), .ZN(new_n342_));
  OAI21_X1  g141(.A(new_n340_), .B1(new_n341_), .B2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(new_n339_), .A2(new_n343_), .A3(KEYINPUT97), .ZN(new_n344_));
  NOR2_X1   g143(.A1(new_n341_), .A2(new_n342_), .ZN(new_n345_));
  INV_X1    g144(.A(KEYINPUT97), .ZN(new_n346_));
  NAND3_X1  g145(.A1(new_n345_), .A2(new_n346_), .A3(new_n318_), .ZN(new_n347_));
  NAND3_X1  g146(.A1(new_n344_), .A2(KEYINPUT4), .A3(new_n347_), .ZN(new_n348_));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n343_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(new_n350_), .ZN(new_n351_));
  NAND2_X1  g150(.A1(G225gat), .A2(G233gat), .ZN(new_n352_));
  INV_X1    g151(.A(new_n352_), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n351_), .A2(new_n353_), .ZN(new_n354_));
  XNOR2_X1  g153(.A(G1gat), .B(G29gat), .ZN(new_n355_));
  XNOR2_X1  g154(.A(new_n355_), .B(G85gat), .ZN(new_n356_));
  XNOR2_X1  g155(.A(KEYINPUT0), .B(G57gat), .ZN(new_n357_));
  XNOR2_X1  g156(.A(new_n356_), .B(new_n357_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n353_), .B1(new_n344_), .B2(new_n347_), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n354_), .A2(new_n359_), .A3(new_n361_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n352_), .B1(new_n348_), .B2(new_n350_), .ZN(new_n363_));
  OAI21_X1  g162(.A(new_n358_), .B1(new_n363_), .B2(new_n360_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n362_), .A2(new_n364_), .ZN(new_n365_));
  AND3_X1   g164(.A1(new_n309_), .A2(new_n315_), .A3(new_n365_), .ZN(new_n366_));
  AOI21_X1  g165(.A(new_n304_), .B1(new_n305_), .B2(new_n274_), .ZN(new_n367_));
  AOI21_X1  g166(.A(new_n295_), .B1(new_n367_), .B2(KEYINPUT95), .ZN(new_n368_));
  NAND2_X1  g167(.A1(new_n300_), .A2(KEYINPUT20), .ZN(new_n369_));
  INV_X1    g168(.A(KEYINPUT95), .ZN(new_n370_));
  NAND2_X1  g169(.A1(new_n369_), .A2(new_n370_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n303_), .B1(new_n368_), .B2(new_n371_), .ZN(new_n372_));
  OAI21_X1  g171(.A(new_n206_), .B1(new_n372_), .B2(new_n313_), .ZN(new_n373_));
  NAND3_X1  g172(.A1(new_n310_), .A2(new_n207_), .A3(new_n314_), .ZN(new_n374_));
  NAND3_X1  g173(.A1(new_n373_), .A2(KEYINPUT96), .A3(new_n374_), .ZN(new_n375_));
  INV_X1    g174(.A(KEYINPUT96), .ZN(new_n376_));
  OAI211_X1 g175(.A(new_n376_), .B(new_n206_), .C1(new_n372_), .C2(new_n313_), .ZN(new_n377_));
  NAND2_X1  g176(.A1(new_n375_), .A2(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n359_), .B1(new_n351_), .B2(new_n352_), .ZN(new_n379_));
  AND3_X1   g178(.A1(new_n344_), .A2(KEYINPUT99), .A3(new_n347_), .ZN(new_n380_));
  AOI21_X1  g179(.A(KEYINPUT99), .B1(new_n344_), .B2(new_n347_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n353_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  NAND2_X1  g181(.A1(new_n379_), .A2(new_n382_), .ZN(new_n383_));
  INV_X1    g182(.A(KEYINPUT33), .ZN(new_n384_));
  OAI21_X1  g183(.A(new_n383_), .B1(new_n362_), .B2(new_n384_), .ZN(new_n385_));
  AOI21_X1  g184(.A(KEYINPUT98), .B1(new_n362_), .B2(new_n384_), .ZN(new_n386_));
  INV_X1    g185(.A(new_n386_), .ZN(new_n387_));
  NAND3_X1  g186(.A1(new_n362_), .A2(KEYINPUT98), .A3(new_n384_), .ZN(new_n388_));
  AOI21_X1  g187(.A(new_n385_), .B1(new_n387_), .B2(new_n388_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n366_), .B1(new_n378_), .B2(new_n389_), .ZN(new_n390_));
  INV_X1    g189(.A(KEYINPUT29), .ZN(new_n391_));
  OAI21_X1  g190(.A(new_n235_), .B1(new_n391_), .B2(new_n345_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n392_), .B(G78gat), .ZN(new_n393_));
  INV_X1    g192(.A(new_n393_), .ZN(new_n394_));
  NAND2_X1  g193(.A1(new_n345_), .A2(new_n391_), .ZN(new_n395_));
  NAND2_X1  g194(.A1(new_n395_), .A2(KEYINPUT28), .ZN(new_n396_));
  INV_X1    g195(.A(KEYINPUT28), .ZN(new_n397_));
  NAND3_X1  g196(.A1(new_n345_), .A2(new_n397_), .A3(new_n391_), .ZN(new_n398_));
  NAND2_X1  g197(.A1(new_n396_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G22gat), .B(G50gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n399_), .A2(new_n400_), .ZN(new_n401_));
  INV_X1    g200(.A(new_n400_), .ZN(new_n402_));
  NAND3_X1  g201(.A1(new_n396_), .A2(new_n398_), .A3(new_n402_), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n401_), .A2(new_n403_), .ZN(new_n404_));
  OAI211_X1 g203(.A(G228gat), .B(G233gat), .C1(new_n305_), .C2(KEYINPUT93), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(new_n405_), .ZN(new_n406_));
  INV_X1    g205(.A(new_n406_), .ZN(new_n407_));
  NOR2_X1   g206(.A1(new_n404_), .A2(new_n405_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n394_), .B1(new_n407_), .B2(new_n408_), .ZN(new_n409_));
  OR2_X1    g208(.A1(new_n404_), .A2(new_n405_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n410_), .A2(new_n406_), .A3(new_n393_), .ZN(new_n411_));
  NAND2_X1  g210(.A1(new_n409_), .A2(new_n411_), .ZN(new_n412_));
  XNOR2_X1  g211(.A(KEYINPUT94), .B(G106gat), .ZN(new_n413_));
  INV_X1    g212(.A(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n412_), .A2(new_n414_), .ZN(new_n415_));
  NAND3_X1  g214(.A1(new_n409_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  OAI21_X1  g216(.A(new_n202_), .B1(new_n390_), .B2(new_n417_), .ZN(new_n418_));
  AND3_X1   g217(.A1(new_n409_), .A2(new_n411_), .A3(new_n413_), .ZN(new_n419_));
  AOI21_X1  g218(.A(new_n413_), .B1(new_n409_), .B2(new_n411_), .ZN(new_n420_));
  NOR2_X1   g219(.A1(new_n419_), .A2(new_n420_), .ZN(new_n421_));
  NOR3_X1   g220(.A1(new_n363_), .A2(new_n358_), .A3(new_n360_), .ZN(new_n422_));
  AOI22_X1  g221(.A1(new_n422_), .A2(KEYINPUT33), .B1(new_n382_), .B2(new_n379_), .ZN(new_n423_));
  INV_X1    g222(.A(KEYINPUT98), .ZN(new_n424_));
  NOR3_X1   g223(.A1(new_n422_), .A2(new_n424_), .A3(KEYINPUT33), .ZN(new_n425_));
  OAI21_X1  g224(.A(new_n423_), .B1(new_n425_), .B2(new_n386_), .ZN(new_n426_));
  AOI21_X1  g225(.A(new_n426_), .B1(new_n377_), .B2(new_n375_), .ZN(new_n427_));
  OAI211_X1 g226(.A(new_n421_), .B(KEYINPUT101), .C1(new_n427_), .C2(new_n366_), .ZN(new_n428_));
  INV_X1    g227(.A(new_n365_), .ZN(new_n429_));
  INV_X1    g228(.A(KEYINPUT27), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n375_), .A2(new_n430_), .A3(new_n377_), .ZN(new_n431_));
  OAI21_X1  g230(.A(new_n206_), .B1(new_n302_), .B2(new_n308_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n432_), .A2(KEYINPUT27), .A3(new_n374_), .ZN(new_n433_));
  NAND4_X1  g232(.A1(new_n417_), .A2(new_n429_), .A3(new_n431_), .A4(new_n433_), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n418_), .A2(new_n428_), .A3(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(KEYINPUT102), .ZN(new_n436_));
  XNOR2_X1  g235(.A(G71gat), .B(G99gat), .ZN(new_n437_));
  XNOR2_X1  g236(.A(KEYINPUT87), .B(G43gat), .ZN(new_n438_));
  XNOR2_X1  g237(.A(new_n437_), .B(new_n438_), .ZN(new_n439_));
  XNOR2_X1  g238(.A(new_n274_), .B(new_n439_), .ZN(new_n440_));
  XOR2_X1   g239(.A(KEYINPUT88), .B(KEYINPUT31), .Z(new_n441_));
  XOR2_X1   g240(.A(new_n440_), .B(new_n441_), .Z(new_n442_));
  NAND2_X1  g241(.A1(G227gat), .A2(G233gat), .ZN(new_n443_));
  XNOR2_X1  g242(.A(new_n443_), .B(G15gat), .ZN(new_n444_));
  XNOR2_X1  g243(.A(new_n444_), .B(KEYINPUT30), .ZN(new_n445_));
  XNOR2_X1  g244(.A(new_n445_), .B(new_n318_), .ZN(new_n446_));
  XOR2_X1   g245(.A(new_n442_), .B(new_n446_), .Z(new_n447_));
  INV_X1    g246(.A(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(new_n435_), .A2(new_n436_), .A3(new_n448_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n431_), .A2(new_n433_), .ZN(new_n450_));
  INV_X1    g249(.A(new_n450_), .ZN(new_n451_));
  NOR2_X1   g250(.A1(new_n448_), .A2(new_n365_), .ZN(new_n452_));
  NAND3_X1  g251(.A1(new_n451_), .A2(new_n421_), .A3(new_n452_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n449_), .A2(new_n453_), .ZN(new_n454_));
  AOI21_X1  g253(.A(new_n436_), .B1(new_n435_), .B2(new_n448_), .ZN(new_n455_));
  NOR2_X1   g254(.A1(new_n454_), .A2(new_n455_), .ZN(new_n456_));
  XOR2_X1   g255(.A(G29gat), .B(G36gat), .Z(new_n457_));
  XOR2_X1   g256(.A(G43gat), .B(G50gat), .Z(new_n458_));
  XNOR2_X1  g257(.A(new_n457_), .B(new_n458_), .ZN(new_n459_));
  XNOR2_X1  g258(.A(KEYINPUT76), .B(KEYINPUT15), .ZN(new_n460_));
  XNOR2_X1  g259(.A(new_n459_), .B(new_n460_), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  XNOR2_X1  g261(.A(G15gat), .B(G22gat), .ZN(new_n463_));
  INV_X1    g262(.A(G1gat), .ZN(new_n464_));
  INV_X1    g263(.A(G8gat), .ZN(new_n465_));
  OAI21_X1  g264(.A(KEYINPUT14), .B1(new_n464_), .B2(new_n465_), .ZN(new_n466_));
  NAND2_X1  g265(.A1(new_n463_), .A2(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G1gat), .B(G8gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n467_), .B(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n462_), .A2(new_n469_), .ZN(new_n470_));
  XOR2_X1   g269(.A(new_n459_), .B(KEYINPUT80), .Z(new_n471_));
  OAI21_X1  g270(.A(new_n470_), .B1(new_n469_), .B2(new_n471_), .ZN(new_n472_));
  NAND2_X1  g271(.A1(G229gat), .A2(G233gat), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  NOR2_X1   g273(.A1(new_n472_), .A2(new_n474_), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n471_), .B(new_n469_), .ZN(new_n476_));
  AOI21_X1  g275(.A(new_n475_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n477_));
  XOR2_X1   g276(.A(G113gat), .B(G141gat), .Z(new_n478_));
  XNOR2_X1  g277(.A(G169gat), .B(G197gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(new_n478_), .B(new_n479_), .ZN(new_n480_));
  OR2_X1    g279(.A1(new_n477_), .A2(new_n480_), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n477_), .A2(new_n480_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n481_), .A2(new_n482_), .ZN(new_n483_));
  INV_X1    g282(.A(new_n483_), .ZN(new_n484_));
  NOR2_X1   g283(.A1(new_n456_), .A2(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(new_n485_), .B(KEYINPUT103), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT37), .ZN(new_n487_));
  XOR2_X1   g286(.A(G85gat), .B(G92gat), .Z(new_n488_));
  INV_X1    g287(.A(KEYINPUT7), .ZN(new_n489_));
  NAND2_X1  g288(.A1(new_n489_), .A2(KEYINPUT66), .ZN(new_n490_));
  NOR2_X1   g289(.A1(G99gat), .A2(G106gat), .ZN(new_n491_));
  XNOR2_X1  g290(.A(new_n490_), .B(new_n491_), .ZN(new_n492_));
  NAND2_X1  g291(.A1(G99gat), .A2(G106gat), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n493_), .A2(KEYINPUT6), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n495_));
  NAND3_X1  g294(.A1(new_n495_), .A2(G99gat), .A3(G106gat), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n494_), .A2(new_n496_), .ZN(new_n497_));
  OAI21_X1  g296(.A(new_n492_), .B1(KEYINPUT70), .B2(new_n497_), .ZN(new_n498_));
  AND2_X1   g297(.A1(new_n497_), .A2(KEYINPUT70), .ZN(new_n499_));
  OAI21_X1  g298(.A(new_n488_), .B1(new_n498_), .B2(new_n499_), .ZN(new_n500_));
  NAND2_X1  g299(.A1(new_n500_), .A2(KEYINPUT8), .ZN(new_n501_));
  INV_X1    g300(.A(KEYINPUT69), .ZN(new_n502_));
  AOI21_X1  g301(.A(KEYINPUT65), .B1(new_n494_), .B2(new_n496_), .ZN(new_n503_));
  INV_X1    g302(.A(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n494_), .A2(new_n496_), .A3(KEYINPUT65), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(new_n492_), .A3(new_n505_), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT67), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n506_), .A2(new_n507_), .ZN(new_n508_));
  INV_X1    g307(.A(new_n505_), .ZN(new_n509_));
  NOR2_X1   g308(.A1(new_n509_), .A2(new_n503_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n510_), .A2(KEYINPUT67), .A3(new_n492_), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n508_), .A2(new_n511_), .ZN(new_n512_));
  INV_X1    g311(.A(KEYINPUT8), .ZN(new_n513_));
  AND2_X1   g312(.A1(new_n513_), .A2(KEYINPUT68), .ZN(new_n514_));
  NOR2_X1   g313(.A1(new_n513_), .A2(KEYINPUT68), .ZN(new_n515_));
  OR2_X1    g314(.A1(new_n514_), .A2(new_n515_), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n516_), .A2(new_n488_), .ZN(new_n517_));
  INV_X1    g316(.A(new_n517_), .ZN(new_n518_));
  AOI21_X1  g317(.A(new_n502_), .B1(new_n512_), .B2(new_n518_), .ZN(new_n519_));
  AOI211_X1 g318(.A(KEYINPUT69), .B(new_n517_), .C1(new_n508_), .C2(new_n511_), .ZN(new_n520_));
  OAI21_X1  g319(.A(new_n501_), .B1(new_n519_), .B2(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n488_), .A2(KEYINPUT9), .ZN(new_n522_));
  NAND2_X1  g321(.A1(G85gat), .A2(G92gat), .ZN(new_n523_));
  XOR2_X1   g322(.A(KEYINPUT10), .B(G99gat), .Z(new_n524_));
  INV_X1    g323(.A(new_n524_), .ZN(new_n525_));
  OAI221_X1 g324(.A(new_n522_), .B1(KEYINPUT9), .B2(new_n523_), .C1(new_n525_), .C2(G106gat), .ZN(new_n526_));
  INV_X1    g325(.A(new_n510_), .ZN(new_n527_));
  NOR2_X1   g326(.A1(new_n526_), .A2(new_n527_), .ZN(new_n528_));
  INV_X1    g327(.A(new_n528_), .ZN(new_n529_));
  AND3_X1   g328(.A1(new_n521_), .A2(new_n459_), .A3(new_n529_), .ZN(new_n530_));
  INV_X1    g329(.A(new_n530_), .ZN(new_n531_));
  XNOR2_X1  g330(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n532_));
  NAND2_X1  g331(.A1(G232gat), .A2(G233gat), .ZN(new_n533_));
  XNOR2_X1  g332(.A(new_n532_), .B(new_n533_), .ZN(new_n534_));
  NAND2_X1  g333(.A1(new_n534_), .A2(KEYINPUT35), .ZN(new_n535_));
  XNOR2_X1  g334(.A(new_n528_), .B(KEYINPUT72), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n461_), .B1(new_n521_), .B2(new_n536_), .ZN(new_n537_));
  INV_X1    g336(.A(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n534_), .A2(KEYINPUT35), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n531_), .A2(new_n535_), .A3(new_n538_), .A4(new_n539_), .ZN(new_n540_));
  OAI211_X1 g339(.A(KEYINPUT35), .B(new_n534_), .C1(new_n530_), .C2(new_n537_), .ZN(new_n541_));
  NAND2_X1  g340(.A1(new_n540_), .A2(new_n541_), .ZN(new_n542_));
  XNOR2_X1  g341(.A(G190gat), .B(G218gat), .ZN(new_n543_));
  XNOR2_X1  g342(.A(G134gat), .B(G162gat), .ZN(new_n544_));
  XNOR2_X1  g343(.A(new_n543_), .B(new_n544_), .ZN(new_n545_));
  XOR2_X1   g344(.A(new_n545_), .B(KEYINPUT36), .Z(new_n546_));
  NAND2_X1  g345(.A1(new_n542_), .A2(new_n546_), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n487_), .B1(new_n547_), .B2(KEYINPUT77), .ZN(new_n548_));
  OR2_X1    g347(.A1(new_n545_), .A2(KEYINPUT36), .ZN(new_n549_));
  OAI21_X1  g348(.A(new_n547_), .B1(new_n549_), .B2(new_n542_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n548_), .A2(new_n550_), .ZN(new_n551_));
  OAI221_X1 g350(.A(new_n547_), .B1(KEYINPUT77), .B2(new_n487_), .C1(new_n549_), .C2(new_n542_), .ZN(new_n552_));
  NAND2_X1  g351(.A1(new_n551_), .A2(new_n552_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(KEYINPUT67), .B1(new_n510_), .B2(new_n492_), .ZN(new_n555_));
  AND4_X1   g354(.A1(KEYINPUT67), .A2(new_n504_), .A3(new_n492_), .A4(new_n505_), .ZN(new_n556_));
  OAI21_X1  g355(.A(new_n518_), .B1(new_n555_), .B2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT69), .ZN(new_n558_));
  NAND3_X1  g357(.A1(new_n512_), .A2(new_n502_), .A3(new_n518_), .ZN(new_n559_));
  AOI22_X1  g358(.A1(new_n558_), .A2(new_n559_), .B1(KEYINPUT8), .B2(new_n500_), .ZN(new_n560_));
  NOR2_X1   g359(.A1(new_n560_), .A2(new_n528_), .ZN(new_n561_));
  XNOR2_X1  g360(.A(G57gat), .B(G64gat), .ZN(new_n562_));
  NAND2_X1  g361(.A1(new_n562_), .A2(KEYINPUT11), .ZN(new_n563_));
  XOR2_X1   g362(.A(G71gat), .B(G78gat), .Z(new_n564_));
  OR2_X1    g363(.A1(new_n563_), .A2(new_n564_), .ZN(new_n565_));
  NOR2_X1   g364(.A1(new_n562_), .A2(KEYINPUT11), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n564_), .ZN(new_n567_));
  OAI21_X1  g366(.A(new_n565_), .B1(new_n566_), .B2(new_n567_), .ZN(new_n568_));
  XOR2_X1   g367(.A(new_n568_), .B(KEYINPUT71), .Z(new_n569_));
  NAND2_X1  g368(.A1(new_n521_), .A2(new_n536_), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT12), .ZN(new_n571_));
  OR2_X1    g370(.A1(new_n568_), .A2(new_n571_), .ZN(new_n572_));
  INV_X1    g371(.A(new_n572_), .ZN(new_n573_));
  AOI22_X1  g372(.A1(new_n561_), .A2(new_n569_), .B1(new_n570_), .B2(new_n573_), .ZN(new_n574_));
  OAI21_X1  g373(.A(new_n571_), .B1(new_n561_), .B2(new_n569_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(G230gat), .A2(G233gat), .ZN(new_n576_));
  XNOR2_X1  g375(.A(new_n576_), .B(KEYINPUT64), .ZN(new_n577_));
  NAND3_X1  g376(.A1(new_n574_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n578_));
  INV_X1    g377(.A(new_n577_), .ZN(new_n579_));
  NAND3_X1  g378(.A1(new_n521_), .A2(new_n569_), .A3(new_n529_), .ZN(new_n580_));
  INV_X1    g379(.A(new_n580_), .ZN(new_n581_));
  AOI21_X1  g380(.A(new_n569_), .B1(new_n521_), .B2(new_n529_), .ZN(new_n582_));
  OAI21_X1  g381(.A(new_n579_), .B1(new_n581_), .B2(new_n582_), .ZN(new_n583_));
  NAND2_X1  g382(.A1(new_n578_), .A2(new_n583_), .ZN(new_n584_));
  XOR2_X1   g383(.A(G120gat), .B(G148gat), .Z(new_n585_));
  XNOR2_X1  g384(.A(G176gat), .B(G204gat), .ZN(new_n586_));
  XNOR2_X1  g385(.A(new_n585_), .B(new_n586_), .ZN(new_n587_));
  XNOR2_X1  g386(.A(KEYINPUT73), .B(KEYINPUT5), .ZN(new_n588_));
  XNOR2_X1  g387(.A(new_n587_), .B(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(new_n589_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n584_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n578_), .A2(new_n583_), .A3(new_n589_), .ZN(new_n592_));
  NAND2_X1  g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  XOR2_X1   g392(.A(KEYINPUT74), .B(KEYINPUT13), .Z(new_n594_));
  NAND2_X1  g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(KEYINPUT13), .ZN(new_n596_));
  OAI211_X1 g395(.A(new_n591_), .B(new_n592_), .C1(KEYINPUT74), .C2(new_n596_), .ZN(new_n597_));
  NAND2_X1  g396(.A1(new_n595_), .A2(new_n597_), .ZN(new_n598_));
  INV_X1    g397(.A(new_n598_), .ZN(new_n599_));
  XOR2_X1   g398(.A(G127gat), .B(G155gat), .Z(new_n600_));
  XNOR2_X1  g399(.A(G183gat), .B(G211gat), .ZN(new_n601_));
  XNOR2_X1  g400(.A(new_n600_), .B(new_n601_), .ZN(new_n602_));
  XNOR2_X1  g401(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n603_));
  XNOR2_X1  g402(.A(new_n602_), .B(new_n603_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT17), .ZN(new_n605_));
  OR2_X1    g404(.A1(new_n604_), .A2(new_n605_), .ZN(new_n606_));
  XNOR2_X1  g405(.A(new_n606_), .B(KEYINPUT79), .ZN(new_n607_));
  NAND2_X1  g406(.A1(G231gat), .A2(G233gat), .ZN(new_n608_));
  XOR2_X1   g407(.A(new_n469_), .B(new_n608_), .Z(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(new_n568_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n607_), .A2(new_n610_), .ZN(new_n611_));
  OR2_X1    g410(.A1(new_n569_), .A2(new_n609_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n569_), .A2(new_n609_), .ZN(new_n613_));
  NAND2_X1  g412(.A1(new_n604_), .A2(new_n605_), .ZN(new_n614_));
  NAND4_X1  g413(.A1(new_n612_), .A2(new_n613_), .A3(new_n606_), .A4(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n611_), .A2(new_n615_), .ZN(new_n616_));
  NOR3_X1   g415(.A1(new_n554_), .A2(new_n599_), .A3(new_n616_), .ZN(new_n617_));
  AND2_X1   g416(.A1(new_n486_), .A2(new_n617_), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n618_), .A2(new_n464_), .A3(new_n365_), .ZN(new_n619_));
  INV_X1    g418(.A(KEYINPUT38), .ZN(new_n620_));
  OR2_X1    g419(.A1(new_n619_), .A2(new_n620_), .ZN(new_n621_));
  INV_X1    g420(.A(new_n550_), .ZN(new_n622_));
  NOR2_X1   g421(.A1(new_n456_), .A2(new_n622_), .ZN(new_n623_));
  NAND2_X1  g422(.A1(new_n598_), .A2(new_n483_), .ZN(new_n624_));
  NOR2_X1   g423(.A1(new_n624_), .A2(new_n616_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  OAI21_X1  g425(.A(G1gat), .B1(new_n626_), .B2(new_n429_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n619_), .A2(new_n620_), .ZN(new_n628_));
  NAND3_X1  g427(.A1(new_n621_), .A2(new_n627_), .A3(new_n628_), .ZN(G1324gat));
  NAND3_X1  g428(.A1(new_n618_), .A2(new_n465_), .A3(new_n450_), .ZN(new_n630_));
  OAI21_X1  g429(.A(G8gat), .B1(new_n626_), .B2(new_n451_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT39), .ZN(new_n632_));
  NAND2_X1  g431(.A1(new_n630_), .A2(new_n632_), .ZN(new_n633_));
  INV_X1    g432(.A(KEYINPUT40), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n633_), .B(new_n634_), .ZN(G1325gat));
  OAI21_X1  g434(.A(G15gat), .B1(new_n626_), .B2(new_n448_), .ZN(new_n636_));
  XOR2_X1   g435(.A(new_n636_), .B(KEYINPUT41), .Z(new_n637_));
  INV_X1    g436(.A(G15gat), .ZN(new_n638_));
  NAND3_X1  g437(.A1(new_n618_), .A2(new_n638_), .A3(new_n447_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n637_), .A2(new_n639_), .ZN(new_n640_));
  INV_X1    g439(.A(KEYINPUT104), .ZN(new_n641_));
  XNOR2_X1  g440(.A(new_n640_), .B(new_n641_), .ZN(G1326gat));
  INV_X1    g441(.A(G22gat), .ZN(new_n643_));
  NAND3_X1  g442(.A1(new_n618_), .A2(new_n643_), .A3(new_n417_), .ZN(new_n644_));
  OAI21_X1  g443(.A(G22gat), .B1(new_n626_), .B2(new_n421_), .ZN(new_n645_));
  XNOR2_X1  g444(.A(new_n645_), .B(KEYINPUT42), .ZN(new_n646_));
  NAND2_X1  g445(.A1(new_n644_), .A2(new_n646_), .ZN(new_n647_));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n648_));
  XNOR2_X1  g447(.A(new_n647_), .B(new_n648_), .ZN(G1327gat));
  INV_X1    g448(.A(new_n616_), .ZN(new_n650_));
  NOR2_X1   g449(.A1(new_n550_), .A2(new_n650_), .ZN(new_n651_));
  INV_X1    g450(.A(new_n651_), .ZN(new_n652_));
  NOR2_X1   g451(.A1(new_n599_), .A2(new_n652_), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n486_), .A2(new_n653_), .ZN(new_n654_));
  OR2_X1    g453(.A1(new_n429_), .A2(G29gat), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n654_), .A2(new_n655_), .ZN(new_n656_));
  NOR2_X1   g455(.A1(new_n624_), .A2(new_n650_), .ZN(new_n657_));
  INV_X1    g456(.A(KEYINPUT43), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n658_), .B(new_n554_), .C1(new_n454_), .C2(new_n455_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n659_), .ZN(new_n660_));
  NAND2_X1  g459(.A1(new_n435_), .A2(new_n448_), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n661_), .A2(KEYINPUT102), .ZN(new_n662_));
  NAND3_X1  g461(.A1(new_n662_), .A2(new_n453_), .A3(new_n449_), .ZN(new_n663_));
  AOI21_X1  g462(.A(new_n658_), .B1(new_n663_), .B2(new_n554_), .ZN(new_n664_));
  OAI21_X1  g463(.A(new_n657_), .B1(new_n660_), .B2(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n665_), .A2(KEYINPUT106), .ZN(new_n666_));
  INV_X1    g465(.A(KEYINPUT44), .ZN(new_n667_));
  INV_X1    g466(.A(new_n657_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n554_), .B1(new_n454_), .B2(new_n455_), .ZN(new_n669_));
  NAND2_X1  g468(.A1(new_n669_), .A2(KEYINPUT43), .ZN(new_n670_));
  AOI21_X1  g469(.A(new_n668_), .B1(new_n670_), .B2(new_n659_), .ZN(new_n671_));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n672_));
  NAND2_X1  g471(.A1(new_n671_), .A2(new_n672_), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n666_), .A2(new_n667_), .A3(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n671_), .A2(KEYINPUT44), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n674_), .A2(new_n365_), .A3(new_n675_), .ZN(new_n676_));
  AOI21_X1  g475(.A(new_n656_), .B1(new_n676_), .B2(G29gat), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n678_));
  NOR2_X1   g477(.A1(new_n677_), .A2(new_n678_), .ZN(new_n679_));
  AOI211_X1 g478(.A(KEYINPUT107), .B(new_n656_), .C1(new_n676_), .C2(G29gat), .ZN(new_n680_));
  NOR2_X1   g479(.A1(new_n679_), .A2(new_n680_), .ZN(G1328gat));
  NOR2_X1   g480(.A1(new_n451_), .A2(G36gat), .ZN(new_n682_));
  NAND3_X1  g481(.A1(new_n486_), .A2(new_n653_), .A3(new_n682_), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n683_), .A2(KEYINPUT45), .ZN(new_n684_));
  INV_X1    g483(.A(KEYINPUT45), .ZN(new_n685_));
  NAND4_X1  g484(.A1(new_n486_), .A2(new_n685_), .A3(new_n653_), .A4(new_n682_), .ZN(new_n686_));
  NAND2_X1  g485(.A1(new_n684_), .A2(new_n686_), .ZN(new_n687_));
  AOI21_X1  g486(.A(new_n451_), .B1(new_n671_), .B2(KEYINPUT44), .ZN(new_n688_));
  OAI21_X1  g487(.A(new_n667_), .B1(new_n671_), .B2(new_n672_), .ZN(new_n689_));
  AOI211_X1 g488(.A(KEYINPUT106), .B(new_n668_), .C1(new_n670_), .C2(new_n659_), .ZN(new_n690_));
  OAI211_X1 g489(.A(KEYINPUT108), .B(new_n688_), .C1(new_n689_), .C2(new_n690_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n691_), .A2(G36gat), .ZN(new_n692_));
  AOI21_X1  g491(.A(KEYINPUT108), .B1(new_n674_), .B2(new_n688_), .ZN(new_n693_));
  OAI21_X1  g492(.A(new_n687_), .B1(new_n692_), .B2(new_n693_), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT46), .ZN(new_n695_));
  NAND2_X1  g494(.A1(new_n694_), .A2(new_n695_), .ZN(new_n696_));
  OAI211_X1 g495(.A(new_n687_), .B(KEYINPUT46), .C1(new_n692_), .C2(new_n693_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n696_), .A2(new_n697_), .ZN(G1329gat));
  NAND4_X1  g497(.A1(new_n674_), .A2(G43gat), .A3(new_n447_), .A4(new_n675_), .ZN(new_n699_));
  INV_X1    g498(.A(G43gat), .ZN(new_n700_));
  OAI21_X1  g499(.A(new_n700_), .B1(new_n654_), .B2(new_n448_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n699_), .A2(new_n701_), .ZN(new_n702_));
  XNOR2_X1  g501(.A(new_n702_), .B(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g502(.A1(new_n674_), .A2(new_n417_), .A3(new_n675_), .ZN(new_n704_));
  NAND2_X1  g503(.A1(new_n704_), .A2(G50gat), .ZN(new_n705_));
  NOR2_X1   g504(.A1(new_n421_), .A2(G50gat), .ZN(new_n706_));
  XNOR2_X1  g505(.A(new_n706_), .B(KEYINPUT109), .ZN(new_n707_));
  OAI21_X1  g506(.A(new_n705_), .B1(new_n654_), .B2(new_n707_), .ZN(G1331gat));
  NOR2_X1   g507(.A1(new_n456_), .A2(new_n483_), .ZN(new_n709_));
  NAND4_X1  g508(.A1(new_n709_), .A2(new_n599_), .A3(new_n650_), .A4(new_n553_), .ZN(new_n710_));
  XNOR2_X1  g509(.A(new_n710_), .B(KEYINPUT110), .ZN(new_n711_));
  INV_X1    g510(.A(G57gat), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n711_), .A2(new_n712_), .A3(new_n365_), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n483_), .A2(new_n616_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n623_), .A2(new_n599_), .A3(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(G57gat), .B1(new_n715_), .B2(new_n429_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n713_), .A2(new_n716_), .ZN(G1332gat));
  OAI21_X1  g516(.A(G64gat), .B1(new_n715_), .B2(new_n451_), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n718_), .B(KEYINPUT48), .ZN(new_n719_));
  INV_X1    g518(.A(G64gat), .ZN(new_n720_));
  NAND3_X1  g519(.A1(new_n711_), .A2(new_n720_), .A3(new_n450_), .ZN(new_n721_));
  NAND2_X1  g520(.A1(new_n719_), .A2(new_n721_), .ZN(G1333gat));
  OAI21_X1  g521(.A(G71gat), .B1(new_n715_), .B2(new_n448_), .ZN(new_n723_));
  XNOR2_X1  g522(.A(new_n723_), .B(KEYINPUT49), .ZN(new_n724_));
  INV_X1    g523(.A(G71gat), .ZN(new_n725_));
  NAND3_X1  g524(.A1(new_n711_), .A2(new_n725_), .A3(new_n447_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1334gat));
  OAI21_X1  g526(.A(G78gat), .B1(new_n715_), .B2(new_n421_), .ZN(new_n728_));
  XNOR2_X1  g527(.A(new_n728_), .B(KEYINPUT50), .ZN(new_n729_));
  INV_X1    g528(.A(G78gat), .ZN(new_n730_));
  NAND3_X1  g529(.A1(new_n711_), .A2(new_n730_), .A3(new_n417_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n729_), .A2(new_n731_), .ZN(G1335gat));
  NOR2_X1   g531(.A1(new_n652_), .A2(new_n598_), .ZN(new_n733_));
  NAND2_X1  g532(.A1(new_n709_), .A2(new_n733_), .ZN(new_n734_));
  NOR3_X1   g533(.A1(new_n734_), .A2(G85gat), .A3(new_n429_), .ZN(new_n735_));
  NAND3_X1  g534(.A1(new_n599_), .A2(new_n484_), .A3(new_n616_), .ZN(new_n736_));
  NOR2_X1   g535(.A1(new_n660_), .A2(new_n664_), .ZN(new_n737_));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n738_));
  NAND2_X1  g537(.A1(new_n737_), .A2(new_n738_), .ZN(new_n739_));
  OAI21_X1  g538(.A(KEYINPUT111), .B1(new_n660_), .B2(new_n664_), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n736_), .B1(new_n739_), .B2(new_n740_), .ZN(new_n741_));
  NAND2_X1  g540(.A1(new_n741_), .A2(new_n365_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n735_), .B1(new_n742_), .B2(G85gat), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n744_));
  XNOR2_X1  g543(.A(new_n743_), .B(new_n744_), .ZN(G1336gat));
  NAND3_X1  g544(.A1(new_n741_), .A2(G92gat), .A3(new_n450_), .ZN(new_n746_));
  INV_X1    g545(.A(G92gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n747_), .B1(new_n734_), .B2(new_n451_), .ZN(new_n748_));
  XNOR2_X1  g547(.A(new_n748_), .B(KEYINPUT113), .ZN(new_n749_));
  AND2_X1   g548(.A1(new_n746_), .A2(new_n749_), .ZN(G1337gat));
  INV_X1    g549(.A(G99gat), .ZN(new_n751_));
  AOI21_X1  g550(.A(new_n751_), .B1(new_n741_), .B2(new_n447_), .ZN(new_n752_));
  INV_X1    g551(.A(new_n752_), .ZN(new_n753_));
  INV_X1    g552(.A(KEYINPUT114), .ZN(new_n754_));
  NOR3_X1   g553(.A1(new_n734_), .A2(new_n448_), .A3(new_n525_), .ZN(new_n755_));
  INV_X1    g554(.A(new_n755_), .ZN(new_n756_));
  NAND4_X1  g555(.A1(new_n753_), .A2(new_n754_), .A3(KEYINPUT51), .A4(new_n756_), .ZN(new_n757_));
  OR2_X1    g556(.A1(new_n754_), .A2(KEYINPUT51), .ZN(new_n758_));
  NAND2_X1  g557(.A1(new_n754_), .A2(KEYINPUT51), .ZN(new_n759_));
  OAI211_X1 g558(.A(new_n758_), .B(new_n759_), .C1(new_n752_), .C2(new_n755_), .ZN(new_n760_));
  AND2_X1   g559(.A1(new_n757_), .A2(new_n760_), .ZN(G1338gat));
  NOR2_X1   g560(.A1(new_n736_), .A2(new_n421_), .ZN(new_n762_));
  INV_X1    g561(.A(new_n762_), .ZN(new_n763_));
  OAI21_X1  g562(.A(G106gat), .B1(new_n737_), .B2(new_n763_), .ZN(new_n764_));
  XNOR2_X1  g563(.A(new_n764_), .B(KEYINPUT52), .ZN(new_n765_));
  OR3_X1    g564(.A1(new_n734_), .A2(G106gat), .A3(new_n421_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n765_), .A2(new_n766_), .ZN(new_n767_));
  XNOR2_X1  g566(.A(new_n767_), .B(KEYINPUT53), .ZN(G1339gat));
  NAND3_X1  g567(.A1(new_n598_), .A2(KEYINPUT115), .A3(new_n714_), .ZN(new_n769_));
  NAND2_X1  g568(.A1(new_n769_), .A2(new_n553_), .ZN(new_n770_));
  AOI21_X1  g569(.A(KEYINPUT115), .B1(new_n598_), .B2(new_n714_), .ZN(new_n771_));
  OAI21_X1  g570(.A(KEYINPUT54), .B1(new_n770_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n771_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT54), .ZN(new_n774_));
  NAND4_X1  g573(.A1(new_n773_), .A2(new_n774_), .A3(new_n553_), .A4(new_n769_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n772_), .A2(new_n775_), .ZN(new_n776_));
  NAND2_X1  g575(.A1(new_n483_), .A2(new_n592_), .ZN(new_n777_));
  INV_X1    g576(.A(KEYINPUT55), .ZN(new_n778_));
  INV_X1    g577(.A(new_n536_), .ZN(new_n779_));
  OAI21_X1  g578(.A(new_n573_), .B1(new_n779_), .B2(new_n560_), .ZN(new_n780_));
  OAI211_X1 g579(.A(new_n780_), .B(new_n580_), .C1(new_n582_), .C2(KEYINPUT12), .ZN(new_n781_));
  OAI21_X1  g580(.A(new_n778_), .B1(new_n781_), .B2(new_n579_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n579_), .ZN(new_n783_));
  NAND4_X1  g582(.A1(new_n574_), .A2(new_n575_), .A3(KEYINPUT55), .A4(new_n577_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n782_), .A2(new_n783_), .A3(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n785_), .A2(new_n590_), .ZN(new_n786_));
  INV_X1    g585(.A(KEYINPUT56), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  NAND3_X1  g587(.A1(new_n785_), .A2(KEYINPUT56), .A3(new_n590_), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n777_), .B1(new_n788_), .B2(new_n789_), .ZN(new_n790_));
  AOI21_X1  g589(.A(new_n473_), .B1(new_n472_), .B2(KEYINPUT116), .ZN(new_n791_));
  OAI21_X1  g590(.A(new_n791_), .B1(KEYINPUT116), .B2(new_n472_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n480_), .B1(new_n476_), .B2(new_n473_), .ZN(new_n793_));
  AOI22_X1  g592(.A1(new_n792_), .A2(new_n793_), .B1(new_n477_), .B2(new_n480_), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n593_), .A2(new_n794_), .ZN(new_n795_));
  INV_X1    g594(.A(new_n795_), .ZN(new_n796_));
  OAI21_X1  g595(.A(new_n550_), .B1(new_n790_), .B2(new_n796_), .ZN(new_n797_));
  NAND2_X1  g596(.A1(new_n797_), .A2(KEYINPUT57), .ZN(new_n798_));
  INV_X1    g597(.A(KEYINPUT57), .ZN(new_n799_));
  OAI211_X1 g598(.A(new_n799_), .B(new_n550_), .C1(new_n790_), .C2(new_n796_), .ZN(new_n800_));
  AND2_X1   g599(.A1(new_n794_), .A2(new_n592_), .ZN(new_n801_));
  INV_X1    g600(.A(new_n789_), .ZN(new_n802_));
  AOI21_X1  g601(.A(KEYINPUT56), .B1(new_n785_), .B2(new_n590_), .ZN(new_n803_));
  OAI21_X1  g602(.A(new_n801_), .B1(new_n802_), .B2(new_n803_), .ZN(new_n804_));
  INV_X1    g603(.A(KEYINPUT58), .ZN(new_n805_));
  OR2_X1    g604(.A1(new_n804_), .A2(new_n805_), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n553_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n807_));
  AOI22_X1  g606(.A1(new_n798_), .A2(new_n800_), .B1(new_n806_), .B2(new_n807_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n616_), .B1(new_n808_), .B2(KEYINPUT117), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n806_), .A2(new_n807_), .ZN(new_n810_));
  OAI211_X1 g609(.A(new_n483_), .B(new_n592_), .C1(new_n802_), .C2(new_n803_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n811_), .A2(new_n795_), .ZN(new_n812_));
  AOI21_X1  g611(.A(new_n799_), .B1(new_n812_), .B2(new_n550_), .ZN(new_n813_));
  INV_X1    g612(.A(new_n800_), .ZN(new_n814_));
  OAI211_X1 g613(.A(KEYINPUT117), .B(new_n810_), .C1(new_n813_), .C2(new_n814_), .ZN(new_n815_));
  INV_X1    g614(.A(new_n815_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n776_), .B1(new_n809_), .B2(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  OAI211_X1 g618(.A(KEYINPUT118), .B(new_n776_), .C1(new_n809_), .C2(new_n816_), .ZN(new_n820_));
  NOR4_X1   g619(.A1(new_n450_), .A2(new_n417_), .A3(new_n448_), .A4(new_n429_), .ZN(new_n821_));
  NAND3_X1  g620(.A1(new_n819_), .A2(new_n820_), .A3(new_n821_), .ZN(new_n822_));
  INV_X1    g621(.A(new_n822_), .ZN(new_n823_));
  INV_X1    g622(.A(G113gat), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n483_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n776_), .B1(new_n808_), .B2(new_n650_), .ZN(new_n826_));
  INV_X1    g625(.A(KEYINPUT59), .ZN(new_n827_));
  NAND2_X1  g626(.A1(new_n821_), .A2(new_n827_), .ZN(new_n828_));
  INV_X1    g627(.A(new_n828_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n826_), .A2(KEYINPUT119), .A3(new_n829_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT119), .B1(new_n826_), .B2(new_n829_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n832_), .B1(new_n822_), .B2(KEYINPUT59), .ZN(new_n833_));
  AND2_X1   g632(.A1(new_n833_), .A2(new_n483_), .ZN(new_n834_));
  OAI21_X1  g633(.A(new_n825_), .B1(new_n834_), .B2(new_n824_), .ZN(G1340gat));
  INV_X1    g634(.A(G120gat), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n836_), .B1(new_n833_), .B2(new_n599_), .ZN(new_n837_));
  OAI21_X1  g636(.A(new_n836_), .B1(new_n598_), .B2(KEYINPUT60), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n838_), .B1(KEYINPUT60), .B2(new_n836_), .ZN(new_n839_));
  NOR2_X1   g638(.A1(new_n822_), .A2(new_n839_), .ZN(new_n840_));
  OAI21_X1  g639(.A(KEYINPUT120), .B1(new_n837_), .B2(new_n840_), .ZN(new_n841_));
  INV_X1    g640(.A(KEYINPUT120), .ZN(new_n842_));
  INV_X1    g641(.A(new_n840_), .ZN(new_n843_));
  AOI211_X1 g642(.A(new_n598_), .B(new_n832_), .C1(new_n822_), .C2(KEYINPUT59), .ZN(new_n844_));
  OAI211_X1 g643(.A(new_n842_), .B(new_n843_), .C1(new_n844_), .C2(new_n836_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n841_), .A2(new_n845_), .ZN(G1341gat));
  INV_X1    g645(.A(G127gat), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n823_), .A2(new_n847_), .A3(new_n650_), .ZN(new_n848_));
  AND2_X1   g647(.A1(new_n833_), .A2(new_n650_), .ZN(new_n849_));
  OAI21_X1  g648(.A(new_n848_), .B1(new_n849_), .B2(new_n847_), .ZN(G1342gat));
  INV_X1    g649(.A(G134gat), .ZN(new_n851_));
  NAND3_X1  g650(.A1(new_n823_), .A2(new_n851_), .A3(new_n622_), .ZN(new_n852_));
  AND2_X1   g651(.A1(new_n833_), .A2(new_n554_), .ZN(new_n853_));
  OAI21_X1  g652(.A(new_n852_), .B1(new_n853_), .B2(new_n851_), .ZN(G1343gat));
  AND2_X1   g653(.A1(new_n819_), .A2(new_n820_), .ZN(new_n855_));
  NAND2_X1  g654(.A1(new_n417_), .A2(new_n448_), .ZN(new_n856_));
  NOR3_X1   g655(.A1(new_n856_), .A2(new_n429_), .A3(new_n450_), .ZN(new_n857_));
  AND2_X1   g656(.A1(new_n855_), .A2(new_n857_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n858_), .A2(new_n483_), .ZN(new_n859_));
  XOR2_X1   g658(.A(KEYINPUT121), .B(G141gat), .Z(new_n860_));
  XNOR2_X1  g659(.A(new_n859_), .B(new_n860_), .ZN(G1344gat));
  NAND2_X1  g660(.A1(new_n858_), .A2(new_n599_), .ZN(new_n862_));
  XNOR2_X1  g661(.A(new_n862_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g662(.A1(new_n858_), .A2(new_n650_), .ZN(new_n864_));
  XNOR2_X1  g663(.A(KEYINPUT61), .B(G155gat), .ZN(new_n865_));
  XNOR2_X1  g664(.A(new_n864_), .B(new_n865_), .ZN(G1346gat));
  INV_X1    g665(.A(G162gat), .ZN(new_n867_));
  NAND3_X1  g666(.A1(new_n858_), .A2(new_n867_), .A3(new_n622_), .ZN(new_n868_));
  AND2_X1   g667(.A1(new_n858_), .A2(new_n554_), .ZN(new_n869_));
  OAI21_X1  g668(.A(new_n868_), .B1(new_n869_), .B2(new_n867_), .ZN(G1347gat));
  NAND2_X1  g669(.A1(new_n452_), .A2(new_n450_), .ZN(new_n871_));
  NOR2_X1   g670(.A1(new_n871_), .A2(new_n417_), .ZN(new_n872_));
  NAND2_X1  g671(.A1(new_n826_), .A2(new_n872_), .ZN(new_n873_));
  OAI21_X1  g672(.A(G169gat), .B1(new_n873_), .B2(new_n484_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(KEYINPUT122), .B(KEYINPUT62), .ZN(new_n875_));
  NOR2_X1   g674(.A1(new_n873_), .A2(new_n484_), .ZN(new_n876_));
  AOI22_X1  g675(.A1(new_n874_), .A2(new_n875_), .B1(new_n876_), .B2(new_n240_), .ZN(new_n877_));
  OAI21_X1  g676(.A(new_n877_), .B1(new_n874_), .B2(new_n875_), .ZN(G1348gat));
  INV_X1    g677(.A(new_n873_), .ZN(new_n879_));
  AOI21_X1  g678(.A(G176gat), .B1(new_n879_), .B2(new_n599_), .ZN(new_n880_));
  AND2_X1   g679(.A1(new_n855_), .A2(new_n421_), .ZN(new_n881_));
  NOR3_X1   g680(.A1(new_n598_), .A2(new_n871_), .A3(new_n280_), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n880_), .B1(new_n881_), .B2(new_n882_), .ZN(G1349gat));
  NOR3_X1   g682(.A1(new_n873_), .A2(new_n266_), .A3(new_n616_), .ZN(new_n884_));
  NAND4_X1  g683(.A1(new_n881_), .A2(new_n450_), .A3(new_n452_), .A4(new_n650_), .ZN(new_n885_));
  AOI21_X1  g684(.A(new_n884_), .B1(new_n885_), .B2(new_n259_), .ZN(G1350gat));
  OAI21_X1  g685(.A(G190gat), .B1(new_n873_), .B2(new_n553_), .ZN(new_n887_));
  XOR2_X1   g686(.A(new_n887_), .B(KEYINPUT123), .Z(new_n888_));
  NAND3_X1  g687(.A1(new_n879_), .A2(new_n267_), .A3(new_n622_), .ZN(new_n889_));
  NAND2_X1  g688(.A1(new_n888_), .A2(new_n889_), .ZN(G1351gat));
  NOR3_X1   g689(.A1(new_n856_), .A2(new_n451_), .A3(new_n365_), .ZN(new_n891_));
  AND2_X1   g690(.A1(new_n855_), .A2(new_n891_), .ZN(new_n892_));
  NAND4_X1  g691(.A1(new_n892_), .A2(KEYINPUT124), .A3(G197gat), .A4(new_n483_), .ZN(new_n893_));
  INV_X1    g692(.A(KEYINPUT124), .ZN(new_n894_));
  NAND3_X1  g693(.A1(new_n855_), .A2(new_n483_), .A3(new_n891_), .ZN(new_n895_));
  OAI21_X1  g694(.A(new_n894_), .B1(new_n895_), .B2(new_n221_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n895_), .A2(new_n221_), .ZN(new_n897_));
  AND3_X1   g696(.A1(new_n893_), .A2(new_n896_), .A3(new_n897_), .ZN(G1352gat));
  NAND2_X1  g697(.A1(new_n855_), .A2(new_n891_), .ZN(new_n899_));
  NOR4_X1   g698(.A1(new_n899_), .A2(KEYINPUT125), .A3(new_n289_), .A4(new_n598_), .ZN(new_n900_));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n901_));
  NOR2_X1   g700(.A1(new_n899_), .A2(new_n598_), .ZN(new_n902_));
  INV_X1    g701(.A(new_n289_), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n901_), .B1(new_n902_), .B2(new_n903_), .ZN(new_n904_));
  OAI21_X1  g703(.A(G204gat), .B1(new_n899_), .B2(new_n598_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n900_), .B1(new_n904_), .B2(new_n905_), .ZN(G1353gat));
  AOI211_X1 g705(.A(KEYINPUT63), .B(G211gat), .C1(new_n892_), .C2(new_n650_), .ZN(new_n907_));
  XNOR2_X1  g706(.A(KEYINPUT63), .B(G211gat), .ZN(new_n908_));
  NOR3_X1   g707(.A1(new_n899_), .A2(new_n616_), .A3(new_n908_), .ZN(new_n909_));
  NOR2_X1   g708(.A1(new_n907_), .A2(new_n909_), .ZN(G1354gat));
  XOR2_X1   g709(.A(KEYINPUT126), .B(G218gat), .Z(new_n911_));
  NOR3_X1   g710(.A1(new_n899_), .A2(new_n553_), .A3(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n892_), .A2(new_n622_), .ZN(new_n913_));
  AOI21_X1  g712(.A(new_n912_), .B1(new_n913_), .B2(new_n911_), .ZN(G1355gat));
endmodule


