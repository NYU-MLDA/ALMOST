//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n665_, new_n666_,
    new_n667_, new_n668_, new_n669_, new_n670_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n733_, new_n734_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n775_, new_n776_, new_n777_, new_n779_,
    new_n780_, new_n781_, new_n782_, new_n783_, new_n784_, new_n785_,
    new_n786_, new_n788_, new_n789_, new_n790_, new_n791_, new_n792_,
    new_n793_, new_n794_, new_n795_, new_n796_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n866_, new_n867_, new_n868_,
    new_n870_, new_n871_, new_n872_, new_n874_, new_n876_, new_n877_,
    new_n878_, new_n880_, new_n881_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n894_, new_n895_, new_n897_, new_n898_, new_n900_,
    new_n901_, new_n902_, new_n904_, new_n905_, new_n906_, new_n907_,
    new_n909_, new_n910_, new_n911_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n918_, new_n919_;
  INV_X1    g000(.A(KEYINPUT102), .ZN(new_n202_));
  XNOR2_X1  g001(.A(KEYINPUT95), .B(G106gat), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  XOR2_X1   g003(.A(KEYINPUT93), .B(KEYINPUT28), .Z(new_n205_));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206_));
  NOR2_X1   g005(.A1(new_n206_), .A2(KEYINPUT1), .ZN(new_n207_));
  NOR2_X1   g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208_));
  OAI21_X1  g007(.A(new_n206_), .B1(new_n208_), .B2(KEYINPUT1), .ZN(new_n209_));
  AOI21_X1  g008(.A(new_n207_), .B1(new_n209_), .B2(KEYINPUT91), .ZN(new_n210_));
  INV_X1    g009(.A(KEYINPUT91), .ZN(new_n211_));
  OAI211_X1 g010(.A(new_n211_), .B(new_n206_), .C1(new_n208_), .C2(KEYINPUT1), .ZN(new_n212_));
  NAND2_X1  g011(.A1(new_n210_), .A2(new_n212_), .ZN(new_n213_));
  NAND2_X1  g012(.A1(G141gat), .A2(G148gat), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216_));
  NOR2_X1   g015(.A1(new_n215_), .A2(new_n216_), .ZN(new_n217_));
  NAND2_X1  g016(.A1(new_n213_), .A2(new_n217_), .ZN(new_n218_));
  INV_X1    g017(.A(KEYINPUT3), .ZN(new_n219_));
  NAND2_X1  g018(.A1(new_n216_), .A2(new_n219_), .ZN(new_n220_));
  INV_X1    g019(.A(KEYINPUT2), .ZN(new_n221_));
  NAND2_X1  g020(.A1(new_n214_), .A2(new_n221_), .ZN(new_n222_));
  NAND3_X1  g021(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n223_));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n224_));
  NAND4_X1  g023(.A1(new_n220_), .A2(new_n222_), .A3(new_n223_), .A4(new_n224_), .ZN(new_n225_));
  INV_X1    g024(.A(new_n206_), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n226_), .A2(new_n208_), .ZN(new_n227_));
  AOI21_X1  g026(.A(KEYINPUT92), .B1(new_n225_), .B2(new_n227_), .ZN(new_n228_));
  AND3_X1   g027(.A1(new_n225_), .A2(KEYINPUT92), .A3(new_n227_), .ZN(new_n229_));
  OAI21_X1  g028(.A(new_n218_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n205_), .B1(new_n230_), .B2(KEYINPUT29), .ZN(new_n231_));
  OR2_X1    g030(.A1(new_n229_), .A2(new_n228_), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT29), .ZN(new_n233_));
  INV_X1    g032(.A(new_n205_), .ZN(new_n234_));
  NAND4_X1  g033(.A1(new_n232_), .A2(new_n233_), .A3(new_n218_), .A4(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n231_), .A2(new_n235_), .ZN(new_n236_));
  XOR2_X1   g035(.A(G22gat), .B(G50gat), .Z(new_n237_));
  INV_X1    g036(.A(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n230_), .A2(KEYINPUT29), .ZN(new_n239_));
  INV_X1    g038(.A(KEYINPUT21), .ZN(new_n240_));
  XNOR2_X1  g039(.A(KEYINPUT94), .B(G204gat), .ZN(new_n241_));
  INV_X1    g040(.A(G197gat), .ZN(new_n242_));
  NOR2_X1   g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  NOR2_X1   g042(.A1(G197gat), .A2(G204gat), .ZN(new_n244_));
  OAI21_X1  g043(.A(new_n240_), .B1(new_n243_), .B2(new_n244_), .ZN(new_n245_));
  XNOR2_X1  g044(.A(G211gat), .B(G218gat), .ZN(new_n246_));
  INV_X1    g045(.A(new_n246_), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n241_), .A2(new_n242_), .ZN(new_n248_));
  AOI21_X1  g047(.A(new_n240_), .B1(G197gat), .B2(G204gat), .ZN(new_n249_));
  AOI21_X1  g048(.A(new_n247_), .B1(new_n248_), .B2(new_n249_), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n243_), .A2(new_n244_), .ZN(new_n251_));
  NOR2_X1   g050(.A1(new_n246_), .A2(new_n240_), .ZN(new_n252_));
  AOI22_X1  g051(.A1(new_n245_), .A2(new_n250_), .B1(new_n251_), .B2(new_n252_), .ZN(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  AOI21_X1  g053(.A(new_n238_), .B1(new_n239_), .B2(new_n254_), .ZN(new_n255_));
  AOI211_X1 g054(.A(new_n237_), .B(new_n253_), .C1(new_n230_), .C2(KEYINPUT29), .ZN(new_n256_));
  OAI21_X1  g055(.A(new_n236_), .B1(new_n255_), .B2(new_n256_), .ZN(new_n257_));
  AOI21_X1  g056(.A(new_n233_), .B1(new_n232_), .B2(new_n218_), .ZN(new_n258_));
  OAI21_X1  g057(.A(new_n237_), .B1(new_n258_), .B2(new_n253_), .ZN(new_n259_));
  NAND3_X1  g058(.A1(new_n239_), .A2(new_n254_), .A3(new_n238_), .ZN(new_n260_));
  NAND4_X1  g059(.A1(new_n259_), .A2(new_n235_), .A3(new_n231_), .A4(new_n260_), .ZN(new_n261_));
  NAND2_X1  g060(.A1(G228gat), .A2(G233gat), .ZN(new_n262_));
  INV_X1    g061(.A(G78gat), .ZN(new_n263_));
  XNOR2_X1  g062(.A(new_n262_), .B(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  AND3_X1   g064(.A1(new_n257_), .A2(new_n261_), .A3(new_n265_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n265_), .B1(new_n257_), .B2(new_n261_), .ZN(new_n267_));
  OAI21_X1  g066(.A(new_n204_), .B1(new_n266_), .B2(new_n267_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n257_), .A2(new_n261_), .ZN(new_n269_));
  NAND2_X1  g068(.A1(new_n269_), .A2(new_n264_), .ZN(new_n270_));
  NAND3_X1  g069(.A1(new_n257_), .A2(new_n261_), .A3(new_n265_), .ZN(new_n271_));
  NAND3_X1  g070(.A1(new_n270_), .A2(new_n203_), .A3(new_n271_), .ZN(new_n272_));
  NAND2_X1  g071(.A1(new_n268_), .A2(new_n272_), .ZN(new_n273_));
  NAND2_X1  g072(.A1(G226gat), .A2(G233gat), .ZN(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT19), .ZN(new_n275_));
  INV_X1    g074(.A(new_n275_), .ZN(new_n276_));
  INV_X1    g075(.A(KEYINPUT20), .ZN(new_n277_));
  XNOR2_X1  g076(.A(KEYINPUT25), .B(G183gat), .ZN(new_n278_));
  XNOR2_X1  g077(.A(KEYINPUT26), .B(G190gat), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n278_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT24), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(G169gat), .B2(G176gat), .ZN(new_n282_));
  INV_X1    g081(.A(G169gat), .ZN(new_n283_));
  INV_X1    g082(.A(G176gat), .ZN(new_n284_));
  NAND3_X1  g083(.A1(new_n283_), .A2(new_n284_), .A3(KEYINPUT84), .ZN(new_n285_));
  INV_X1    g084(.A(KEYINPUT84), .ZN(new_n286_));
  OAI21_X1  g085(.A(new_n286_), .B1(G169gat), .B2(G176gat), .ZN(new_n287_));
  NAND3_X1  g086(.A1(new_n282_), .A2(new_n285_), .A3(new_n287_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n280_), .A2(new_n288_), .ZN(new_n289_));
  OR2_X1    g088(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n290_));
  AND2_X1   g089(.A1(G183gat), .A2(G190gat), .ZN(new_n291_));
  NAND2_X1  g090(.A1(KEYINPUT85), .A2(KEYINPUT23), .ZN(new_n292_));
  NAND3_X1  g091(.A1(new_n290_), .A2(new_n291_), .A3(new_n292_), .ZN(new_n293_));
  NAND2_X1  g092(.A1(new_n293_), .A2(KEYINPUT89), .ZN(new_n294_));
  INV_X1    g093(.A(KEYINPUT89), .ZN(new_n295_));
  NAND4_X1  g094(.A1(new_n290_), .A2(new_n291_), .A3(new_n295_), .A4(new_n292_), .ZN(new_n296_));
  INV_X1    g095(.A(new_n291_), .ZN(new_n297_));
  NAND2_X1  g096(.A1(new_n297_), .A2(KEYINPUT23), .ZN(new_n298_));
  NAND3_X1  g097(.A1(new_n294_), .A2(new_n296_), .A3(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(new_n285_), .A2(new_n287_), .ZN(new_n300_));
  NAND2_X1  g099(.A1(new_n300_), .A2(new_n281_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  AOI21_X1  g101(.A(new_n289_), .B1(new_n302_), .B2(KEYINPUT96), .ZN(new_n303_));
  AOI22_X1  g102(.A1(new_n293_), .A2(KEYINPUT89), .B1(KEYINPUT23), .B2(new_n297_), .ZN(new_n304_));
  AOI22_X1  g103(.A1(new_n304_), .A2(new_n296_), .B1(new_n281_), .B2(new_n300_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT96), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n305_), .A2(new_n306_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n291_), .B1(new_n290_), .B2(new_n292_), .ZN(new_n308_));
  INV_X1    g107(.A(KEYINPUT86), .ZN(new_n309_));
  NAND2_X1  g108(.A1(new_n308_), .A2(new_n309_), .ZN(new_n310_));
  OAI21_X1  g109(.A(KEYINPUT86), .B1(new_n297_), .B2(KEYINPUT23), .ZN(new_n311_));
  OAI21_X1  g110(.A(new_n310_), .B1(new_n308_), .B2(new_n311_), .ZN(new_n312_));
  NOR2_X1   g111(.A1(G183gat), .A2(G190gat), .ZN(new_n313_));
  OR2_X1    g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(KEYINPUT87), .B(G176gat), .ZN(new_n315_));
  XNOR2_X1  g114(.A(KEYINPUT22), .B(G169gat), .ZN(new_n316_));
  AOI22_X1  g115(.A1(new_n315_), .A2(new_n316_), .B1(G169gat), .B2(G176gat), .ZN(new_n317_));
  AOI22_X1  g116(.A1(new_n303_), .A2(new_n307_), .B1(new_n314_), .B2(new_n317_), .ZN(new_n318_));
  AOI21_X1  g117(.A(new_n277_), .B1(new_n318_), .B2(new_n253_), .ZN(new_n319_));
  INV_X1    g118(.A(KEYINPUT97), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n315_), .A2(new_n316_), .ZN(new_n321_));
  OR2_X1    g120(.A1(new_n321_), .A2(KEYINPUT88), .ZN(new_n322_));
  NAND2_X1  g121(.A1(new_n321_), .A2(KEYINPUT88), .ZN(new_n323_));
  AOI22_X1  g122(.A1(new_n322_), .A2(new_n323_), .B1(G169gat), .B2(G176gat), .ZN(new_n324_));
  INV_X1    g123(.A(KEYINPUT90), .ZN(new_n325_));
  AOI211_X1 g124(.A(new_n325_), .B(new_n313_), .C1(new_n304_), .C2(new_n296_), .ZN(new_n326_));
  INV_X1    g125(.A(new_n313_), .ZN(new_n327_));
  AOI21_X1  g126(.A(KEYINPUT90), .B1(new_n299_), .B2(new_n327_), .ZN(new_n328_));
  OAI21_X1  g127(.A(new_n324_), .B1(new_n326_), .B2(new_n328_), .ZN(new_n329_));
  NOR2_X1   g128(.A1(new_n278_), .A2(KEYINPUT83), .ZN(new_n330_));
  INV_X1    g129(.A(G183gat), .ZN(new_n331_));
  OAI21_X1  g130(.A(KEYINPUT83), .B1(new_n331_), .B2(KEYINPUT25), .ZN(new_n332_));
  NAND2_X1  g131(.A1(new_n279_), .A2(new_n332_), .ZN(new_n333_));
  NOR2_X1   g132(.A1(new_n330_), .A2(new_n333_), .ZN(new_n334_));
  NAND2_X1  g133(.A1(new_n301_), .A2(new_n288_), .ZN(new_n335_));
  NOR3_X1   g134(.A1(new_n312_), .A2(new_n334_), .A3(new_n335_), .ZN(new_n336_));
  INV_X1    g135(.A(new_n336_), .ZN(new_n337_));
  NAND2_X1  g136(.A1(new_n329_), .A2(new_n337_), .ZN(new_n338_));
  AOI21_X1  g137(.A(new_n320_), .B1(new_n338_), .B2(new_n254_), .ZN(new_n339_));
  AOI211_X1 g138(.A(KEYINPUT97), .B(new_n253_), .C1(new_n329_), .C2(new_n337_), .ZN(new_n340_));
  OAI211_X1 g139(.A(new_n276_), .B(new_n319_), .C1(new_n339_), .C2(new_n340_), .ZN(new_n341_));
  NAND3_X1  g140(.A1(new_n329_), .A2(new_n253_), .A3(new_n337_), .ZN(new_n342_));
  OAI211_X1 g141(.A(new_n342_), .B(KEYINPUT20), .C1(new_n253_), .C2(new_n318_), .ZN(new_n343_));
  NAND2_X1  g142(.A1(new_n343_), .A2(new_n275_), .ZN(new_n344_));
  XNOR2_X1  g143(.A(G8gat), .B(G36gat), .ZN(new_n345_));
  XNOR2_X1  g144(.A(new_n345_), .B(KEYINPUT18), .ZN(new_n346_));
  XNOR2_X1  g145(.A(G64gat), .B(G92gat), .ZN(new_n347_));
  XOR2_X1   g146(.A(new_n346_), .B(new_n347_), .Z(new_n348_));
  NAND3_X1  g147(.A1(new_n341_), .A2(new_n344_), .A3(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n349_), .A2(KEYINPUT27), .ZN(new_n350_));
  OAI21_X1  g149(.A(new_n317_), .B1(new_n312_), .B2(new_n313_), .ZN(new_n351_));
  OAI211_X1 g150(.A(new_n288_), .B(new_n280_), .C1(new_n305_), .C2(new_n306_), .ZN(new_n352_));
  NOR2_X1   g151(.A1(new_n302_), .A2(KEYINPUT96), .ZN(new_n353_));
  OAI21_X1  g152(.A(new_n351_), .B1(new_n352_), .B2(new_n353_), .ZN(new_n354_));
  OAI21_X1  g153(.A(KEYINPUT20), .B1(new_n354_), .B2(new_n254_), .ZN(new_n355_));
  NAND2_X1  g154(.A1(new_n299_), .A2(new_n327_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n356_), .A2(new_n325_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(new_n299_), .A2(KEYINPUT90), .A3(new_n327_), .ZN(new_n358_));
  NAND2_X1  g157(.A1(new_n357_), .A2(new_n358_), .ZN(new_n359_));
  AOI21_X1  g158(.A(new_n336_), .B1(new_n359_), .B2(new_n324_), .ZN(new_n360_));
  OAI21_X1  g159(.A(KEYINPUT97), .B1(new_n360_), .B2(new_n253_), .ZN(new_n361_));
  NAND3_X1  g160(.A1(new_n338_), .A2(new_n320_), .A3(new_n254_), .ZN(new_n362_));
  AOI21_X1  g161(.A(new_n355_), .B1(new_n361_), .B2(new_n362_), .ZN(new_n363_));
  OAI21_X1  g162(.A(KEYINPUT100), .B1(new_n363_), .B2(new_n276_), .ZN(new_n364_));
  OAI21_X1  g163(.A(new_n319_), .B1(new_n339_), .B2(new_n340_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT100), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n365_), .A2(new_n366_), .A3(new_n275_), .ZN(new_n367_));
  NOR2_X1   g166(.A1(new_n343_), .A2(new_n275_), .ZN(new_n368_));
  INV_X1    g167(.A(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n364_), .A2(new_n367_), .A3(new_n369_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n348_), .ZN(new_n371_));
  AOI21_X1  g170(.A(new_n350_), .B1(new_n370_), .B2(new_n371_), .ZN(new_n372_));
  AOI21_X1  g171(.A(new_n348_), .B1(new_n341_), .B2(new_n344_), .ZN(new_n373_));
  INV_X1    g172(.A(new_n373_), .ZN(new_n374_));
  AOI21_X1  g173(.A(KEYINPUT27), .B1(new_n374_), .B2(new_n349_), .ZN(new_n375_));
  OAI21_X1  g174(.A(KEYINPUT101), .B1(new_n372_), .B2(new_n375_), .ZN(new_n376_));
  INV_X1    g175(.A(KEYINPUT101), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT27), .ZN(new_n378_));
  INV_X1    g177(.A(new_n349_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n378_), .B1(new_n379_), .B2(new_n373_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n365_), .A2(new_n275_), .ZN(new_n381_));
  AOI21_X1  g180(.A(new_n368_), .B1(new_n381_), .B2(KEYINPUT100), .ZN(new_n382_));
  AOI21_X1  g181(.A(new_n348_), .B1(new_n382_), .B2(new_n367_), .ZN(new_n383_));
  OAI211_X1 g182(.A(new_n377_), .B(new_n380_), .C1(new_n383_), .C2(new_n350_), .ZN(new_n384_));
  AOI21_X1  g183(.A(new_n273_), .B1(new_n376_), .B2(new_n384_), .ZN(new_n385_));
  XNOR2_X1  g184(.A(G71gat), .B(G99gat), .ZN(new_n386_));
  XNOR2_X1  g185(.A(new_n386_), .B(G43gat), .ZN(new_n387_));
  XNOR2_X1  g186(.A(new_n338_), .B(new_n387_), .ZN(new_n388_));
  XOR2_X1   g187(.A(G127gat), .B(G134gat), .Z(new_n389_));
  XOR2_X1   g188(.A(G113gat), .B(G120gat), .Z(new_n390_));
  XNOR2_X1  g189(.A(new_n389_), .B(new_n390_), .ZN(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  XNOR2_X1  g191(.A(new_n388_), .B(new_n392_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(G227gat), .A2(G233gat), .ZN(new_n394_));
  INV_X1    g193(.A(G15gat), .ZN(new_n395_));
  XNOR2_X1  g194(.A(new_n394_), .B(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(new_n396_), .B(KEYINPUT30), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(KEYINPUT31), .ZN(new_n398_));
  OR2_X1    g197(.A1(new_n393_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G1gat), .B(G29gat), .ZN(new_n400_));
  XNOR2_X1  g199(.A(new_n400_), .B(G85gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT0), .B(G57gat), .ZN(new_n402_));
  XOR2_X1   g201(.A(new_n401_), .B(new_n402_), .Z(new_n403_));
  INV_X1    g202(.A(new_n403_), .ZN(new_n404_));
  NAND2_X1  g203(.A1(G225gat), .A2(G233gat), .ZN(new_n405_));
  INV_X1    g204(.A(new_n405_), .ZN(new_n406_));
  NOR2_X1   g205(.A1(new_n229_), .A2(new_n228_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n217_), .ZN(new_n408_));
  AOI21_X1  g207(.A(new_n408_), .B1(new_n210_), .B2(new_n212_), .ZN(new_n409_));
  OAI21_X1  g208(.A(new_n392_), .B1(new_n407_), .B2(new_n409_), .ZN(new_n410_));
  OAI211_X1 g209(.A(new_n218_), .B(new_n391_), .C1(new_n228_), .C2(new_n229_), .ZN(new_n411_));
  NAND3_X1  g210(.A1(new_n410_), .A2(new_n411_), .A3(KEYINPUT4), .ZN(new_n412_));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n413_));
  OAI211_X1 g212(.A(new_n413_), .B(new_n392_), .C1(new_n407_), .C2(new_n409_), .ZN(new_n414_));
  INV_X1    g213(.A(KEYINPUT98), .ZN(new_n415_));
  NAND2_X1  g214(.A1(new_n414_), .A2(new_n415_), .ZN(new_n416_));
  NAND4_X1  g215(.A1(new_n230_), .A2(KEYINPUT98), .A3(new_n413_), .A4(new_n392_), .ZN(new_n417_));
  AND4_X1   g216(.A1(new_n406_), .A2(new_n412_), .A3(new_n416_), .A4(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n410_), .A2(new_n411_), .A3(new_n405_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT99), .ZN(new_n420_));
  INV_X1    g219(.A(KEYINPUT99), .ZN(new_n421_));
  NAND4_X1  g220(.A1(new_n410_), .A2(new_n411_), .A3(new_n421_), .A4(new_n405_), .ZN(new_n422_));
  NAND2_X1  g221(.A1(new_n420_), .A2(new_n422_), .ZN(new_n423_));
  OAI21_X1  g222(.A(new_n404_), .B1(new_n418_), .B2(new_n423_), .ZN(new_n424_));
  NAND4_X1  g223(.A1(new_n412_), .A2(new_n416_), .A3(new_n417_), .A4(new_n406_), .ZN(new_n425_));
  NAND4_X1  g224(.A1(new_n425_), .A2(new_n403_), .A3(new_n420_), .A4(new_n422_), .ZN(new_n426_));
  NAND2_X1  g225(.A1(new_n424_), .A2(new_n426_), .ZN(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n393_), .A2(new_n398_), .ZN(new_n429_));
  NAND3_X1  g228(.A1(new_n399_), .A2(new_n428_), .A3(new_n429_), .ZN(new_n430_));
  INV_X1    g229(.A(new_n430_), .ZN(new_n431_));
  INV_X1    g230(.A(new_n273_), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n348_), .A2(KEYINPUT32), .ZN(new_n433_));
  NAND3_X1  g232(.A1(new_n341_), .A2(new_n344_), .A3(new_n433_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n427_), .A2(new_n434_), .ZN(new_n435_));
  INV_X1    g234(.A(new_n433_), .ZN(new_n436_));
  AOI21_X1  g235(.A(new_n435_), .B1(new_n370_), .B2(new_n436_), .ZN(new_n437_));
  INV_X1    g236(.A(new_n423_), .ZN(new_n438_));
  NAND4_X1  g237(.A1(new_n438_), .A2(KEYINPUT33), .A3(new_n403_), .A4(new_n425_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT33), .ZN(new_n440_));
  NAND2_X1  g239(.A1(new_n426_), .A2(new_n440_), .ZN(new_n441_));
  NAND4_X1  g240(.A1(new_n412_), .A2(new_n416_), .A3(new_n417_), .A4(new_n405_), .ZN(new_n442_));
  NAND2_X1  g241(.A1(new_n410_), .A2(new_n411_), .ZN(new_n443_));
  OAI211_X1 g242(.A(new_n442_), .B(new_n404_), .C1(new_n405_), .C2(new_n443_), .ZN(new_n444_));
  NAND3_X1  g243(.A1(new_n439_), .A2(new_n441_), .A3(new_n444_), .ZN(new_n445_));
  NOR3_X1   g244(.A1(new_n445_), .A2(new_n379_), .A3(new_n373_), .ZN(new_n446_));
  OAI21_X1  g245(.A(new_n432_), .B1(new_n437_), .B2(new_n446_), .ZN(new_n447_));
  AOI21_X1  g246(.A(new_n427_), .B1(new_n268_), .B2(new_n272_), .ZN(new_n448_));
  OAI211_X1 g247(.A(new_n448_), .B(new_n380_), .C1(new_n383_), .C2(new_n350_), .ZN(new_n449_));
  NAND2_X1  g248(.A1(new_n447_), .A2(new_n449_), .ZN(new_n450_));
  NAND2_X1  g249(.A1(new_n399_), .A2(new_n429_), .ZN(new_n451_));
  AOI22_X1  g250(.A1(new_n385_), .A2(new_n431_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  INV_X1    g251(.A(new_n452_), .ZN(new_n453_));
  XNOR2_X1  g252(.A(G15gat), .B(G22gat), .ZN(new_n454_));
  INV_X1    g253(.A(G1gat), .ZN(new_n455_));
  INV_X1    g254(.A(G8gat), .ZN(new_n456_));
  OAI21_X1  g255(.A(KEYINPUT14), .B1(new_n455_), .B2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n454_), .A2(new_n457_), .ZN(new_n458_));
  XOR2_X1   g257(.A(G1gat), .B(G8gat), .Z(new_n459_));
  XNOR2_X1  g258(.A(new_n458_), .B(new_n459_), .ZN(new_n460_));
  XNOR2_X1  g259(.A(KEYINPUT79), .B(KEYINPUT80), .ZN(new_n461_));
  INV_X1    g260(.A(new_n461_), .ZN(new_n462_));
  OR2_X1    g261(.A1(new_n460_), .A2(new_n462_), .ZN(new_n463_));
  NAND2_X1  g262(.A1(new_n460_), .A2(new_n462_), .ZN(new_n464_));
  NAND2_X1  g263(.A1(new_n463_), .A2(new_n464_), .ZN(new_n465_));
  XNOR2_X1  g264(.A(G29gat), .B(G36gat), .ZN(new_n466_));
  XNOR2_X1  g265(.A(G43gat), .B(G50gat), .ZN(new_n467_));
  XNOR2_X1  g266(.A(new_n466_), .B(new_n467_), .ZN(new_n468_));
  INV_X1    g267(.A(new_n468_), .ZN(new_n469_));
  NOR2_X1   g268(.A1(new_n465_), .A2(new_n469_), .ZN(new_n470_));
  XNOR2_X1  g269(.A(new_n470_), .B(KEYINPUT82), .ZN(new_n471_));
  NAND2_X1  g270(.A1(G229gat), .A2(G233gat), .ZN(new_n472_));
  XNOR2_X1  g271(.A(new_n468_), .B(KEYINPUT15), .ZN(new_n473_));
  NAND2_X1  g272(.A1(new_n465_), .A2(new_n473_), .ZN(new_n474_));
  NAND3_X1  g273(.A1(new_n471_), .A2(new_n472_), .A3(new_n474_), .ZN(new_n475_));
  NAND2_X1  g274(.A1(new_n465_), .A2(new_n469_), .ZN(new_n476_));
  AND2_X1   g275(.A1(new_n471_), .A2(new_n476_), .ZN(new_n477_));
  OAI21_X1  g276(.A(new_n475_), .B1(new_n477_), .B2(new_n472_), .ZN(new_n478_));
  XNOR2_X1  g277(.A(G113gat), .B(G141gat), .ZN(new_n479_));
  XNOR2_X1  g278(.A(G169gat), .B(G197gat), .ZN(new_n480_));
  XOR2_X1   g279(.A(new_n479_), .B(new_n480_), .Z(new_n481_));
  INV_X1    g280(.A(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(new_n478_), .A2(new_n482_), .ZN(new_n483_));
  OAI211_X1 g282(.A(new_n475_), .B(new_n481_), .C1(new_n477_), .C2(new_n472_), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  AOI21_X1  g284(.A(new_n202_), .B1(new_n453_), .B2(new_n485_), .ZN(new_n486_));
  INV_X1    g285(.A(new_n485_), .ZN(new_n487_));
  NOR3_X1   g286(.A1(new_n452_), .A2(KEYINPUT102), .A3(new_n487_), .ZN(new_n488_));
  NOR2_X1   g287(.A1(new_n486_), .A2(new_n488_), .ZN(new_n489_));
  XNOR2_X1  g288(.A(KEYINPUT75), .B(KEYINPUT13), .ZN(new_n490_));
  XOR2_X1   g289(.A(G120gat), .B(G148gat), .Z(new_n491_));
  XNOR2_X1  g290(.A(new_n491_), .B(KEYINPUT72), .ZN(new_n492_));
  XOR2_X1   g291(.A(G176gat), .B(G204gat), .Z(new_n493_));
  XNOR2_X1  g292(.A(new_n492_), .B(new_n493_), .ZN(new_n494_));
  XOR2_X1   g293(.A(KEYINPUT71), .B(KEYINPUT5), .Z(new_n495_));
  XNOR2_X1  g294(.A(new_n494_), .B(new_n495_), .ZN(new_n496_));
  XNOR2_X1  g295(.A(new_n496_), .B(KEYINPUT73), .ZN(new_n497_));
  NAND2_X1  g296(.A1(G99gat), .A2(G106gat), .ZN(new_n498_));
  INV_X1    g297(.A(KEYINPUT6), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n498_), .A2(new_n499_), .ZN(new_n500_));
  NAND3_X1  g299(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n501_));
  OAI21_X1  g300(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n502_));
  NAND3_X1  g301(.A1(new_n500_), .A2(new_n501_), .A3(new_n502_), .ZN(new_n503_));
  NOR4_X1   g302(.A1(KEYINPUT65), .A2(KEYINPUT7), .A3(G99gat), .A4(G106gat), .ZN(new_n504_));
  INV_X1    g303(.A(KEYINPUT65), .ZN(new_n505_));
  NOR2_X1   g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506_));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n507_));
  AOI21_X1  g306(.A(new_n505_), .B1(new_n506_), .B2(new_n507_), .ZN(new_n508_));
  NOR3_X1   g307(.A1(new_n503_), .A2(new_n504_), .A3(new_n508_), .ZN(new_n509_));
  INV_X1    g308(.A(G85gat), .ZN(new_n510_));
  INV_X1    g309(.A(G92gat), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n510_), .A2(new_n511_), .ZN(new_n512_));
  NAND2_X1  g311(.A1(G85gat), .A2(G92gat), .ZN(new_n513_));
  NAND2_X1  g312(.A1(new_n512_), .A2(new_n513_), .ZN(new_n514_));
  OAI21_X1  g313(.A(KEYINPUT8), .B1(new_n509_), .B2(new_n514_), .ZN(new_n515_));
  INV_X1    g314(.A(new_n508_), .ZN(new_n516_));
  INV_X1    g315(.A(new_n501_), .ZN(new_n517_));
  AOI21_X1  g316(.A(KEYINPUT6), .B1(G99gat), .B2(G106gat), .ZN(new_n518_));
  NOR2_X1   g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  NAND3_X1  g318(.A1(new_n506_), .A2(new_n505_), .A3(new_n507_), .ZN(new_n520_));
  NAND4_X1  g319(.A1(new_n516_), .A2(new_n519_), .A3(new_n502_), .A4(new_n520_), .ZN(new_n521_));
  INV_X1    g320(.A(KEYINPUT8), .ZN(new_n522_));
  INV_X1    g321(.A(new_n514_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n522_), .A3(new_n523_), .ZN(new_n524_));
  NAND2_X1  g323(.A1(new_n515_), .A2(new_n524_), .ZN(new_n525_));
  OR2_X1    g324(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n526_));
  INV_X1    g325(.A(G106gat), .ZN(new_n527_));
  NAND2_X1  g326(.A1(KEYINPUT10), .A2(G99gat), .ZN(new_n528_));
  NAND3_X1  g327(.A1(new_n526_), .A2(new_n527_), .A3(new_n528_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n512_), .A2(KEYINPUT9), .A3(new_n513_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n529_), .A2(new_n530_), .ZN(new_n531_));
  INV_X1    g330(.A(KEYINPUT9), .ZN(new_n532_));
  NAND3_X1  g331(.A1(new_n532_), .A2(G85gat), .A3(G92gat), .ZN(new_n533_));
  NAND3_X1  g332(.A1(new_n500_), .A2(new_n533_), .A3(new_n501_), .ZN(new_n534_));
  OAI21_X1  g333(.A(KEYINPUT64), .B1(new_n531_), .B2(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n534_), .ZN(new_n536_));
  INV_X1    g335(.A(KEYINPUT64), .ZN(new_n537_));
  NAND4_X1  g336(.A1(new_n536_), .A2(new_n537_), .A3(new_n529_), .A4(new_n530_), .ZN(new_n538_));
  AND2_X1   g337(.A1(new_n535_), .A2(new_n538_), .ZN(new_n539_));
  XNOR2_X1  g338(.A(G57gat), .B(G64gat), .ZN(new_n540_));
  NAND2_X1  g339(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n541_));
  XOR2_X1   g340(.A(G71gat), .B(G78gat), .Z(new_n542_));
  AND2_X1   g341(.A1(new_n541_), .A2(new_n542_), .ZN(new_n543_));
  OR2_X1    g342(.A1(new_n540_), .A2(KEYINPUT11), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n543_), .A2(new_n544_), .ZN(new_n545_));
  NOR2_X1   g344(.A1(new_n541_), .A2(new_n542_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n546_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n545_), .A2(new_n547_), .ZN(new_n548_));
  NAND3_X1  g347(.A1(new_n525_), .A2(new_n539_), .A3(new_n548_), .ZN(new_n549_));
  AOI21_X1  g348(.A(new_n548_), .B1(new_n525_), .B2(new_n539_), .ZN(new_n550_));
  INV_X1    g349(.A(KEYINPUT66), .ZN(new_n551_));
  OAI21_X1  g350(.A(new_n549_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND4_X1  g351(.A1(new_n525_), .A2(new_n548_), .A3(new_n539_), .A4(KEYINPUT66), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n552_), .A2(new_n553_), .ZN(new_n554_));
  NAND2_X1  g353(.A1(G230gat), .A2(G233gat), .ZN(new_n555_));
  INV_X1    g354(.A(new_n555_), .ZN(new_n556_));
  NAND2_X1  g355(.A1(new_n554_), .A2(new_n556_), .ZN(new_n557_));
  NAND2_X1  g356(.A1(new_n557_), .A2(KEYINPUT67), .ZN(new_n558_));
  INV_X1    g357(.A(KEYINPUT67), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n554_), .A2(new_n559_), .A3(new_n556_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n546_), .B1(new_n543_), .B2(new_n544_), .ZN(new_n561_));
  NAND2_X1  g360(.A1(new_n561_), .A2(KEYINPUT12), .ZN(new_n562_));
  INV_X1    g361(.A(new_n562_), .ZN(new_n563_));
  NAND3_X1  g362(.A1(new_n535_), .A2(new_n538_), .A3(KEYINPUT68), .ZN(new_n564_));
  NOR3_X1   g363(.A1(new_n509_), .A2(KEYINPUT8), .A3(new_n514_), .ZN(new_n565_));
  AOI21_X1  g364(.A(new_n522_), .B1(new_n521_), .B2(new_n523_), .ZN(new_n566_));
  OAI21_X1  g365(.A(new_n564_), .B1(new_n565_), .B2(new_n566_), .ZN(new_n567_));
  AOI21_X1  g366(.A(KEYINPUT68), .B1(new_n535_), .B2(new_n538_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n563_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT69), .ZN(new_n570_));
  XNOR2_X1  g369(.A(KEYINPUT70), .B(KEYINPUT12), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n549_), .A2(new_n571_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n525_), .A2(new_n539_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n573_), .A2(new_n561_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n572_), .A2(new_n574_), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT69), .ZN(new_n576_));
  OAI211_X1 g375(.A(new_n563_), .B(new_n576_), .C1(new_n567_), .C2(new_n568_), .ZN(new_n577_));
  NAND4_X1  g376(.A1(new_n570_), .A2(new_n575_), .A3(new_n555_), .A4(new_n577_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n558_), .A2(new_n560_), .A3(new_n578_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n558_), .A2(new_n496_), .A3(new_n560_), .A4(new_n578_), .ZN(new_n580_));
  NAND2_X1  g379(.A1(new_n580_), .A2(KEYINPUT74), .ZN(new_n581_));
  AND4_X1   g380(.A1(new_n555_), .A2(new_n570_), .A3(new_n575_), .A4(new_n577_), .ZN(new_n582_));
  AOI21_X1  g381(.A(new_n559_), .B1(new_n554_), .B2(new_n556_), .ZN(new_n583_));
  NOR2_X1   g382(.A1(new_n582_), .A2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(KEYINPUT74), .ZN(new_n585_));
  NAND4_X1  g384(.A1(new_n584_), .A2(new_n585_), .A3(new_n496_), .A4(new_n560_), .ZN(new_n586_));
  AOI221_X4 g385(.A(new_n490_), .B1(new_n497_), .B2(new_n579_), .C1(new_n581_), .C2(new_n586_), .ZN(new_n587_));
  INV_X1    g386(.A(KEYINPUT75), .ZN(new_n588_));
  NOR2_X1   g387(.A1(new_n588_), .A2(KEYINPUT13), .ZN(new_n589_));
  NAND2_X1  g388(.A1(new_n581_), .A2(new_n586_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n579_), .A2(new_n497_), .ZN(new_n591_));
  AOI21_X1  g390(.A(new_n589_), .B1(new_n590_), .B2(new_n591_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n587_), .A2(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(new_n593_), .ZN(new_n594_));
  OAI21_X1  g393(.A(new_n473_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n595_));
  NAND2_X1  g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596_));
  XNOR2_X1  g395(.A(new_n596_), .B(KEYINPUT34), .ZN(new_n597_));
  OAI221_X1 g396(.A(new_n595_), .B1(KEYINPUT35), .B2(new_n597_), .C1(new_n469_), .C2(new_n573_), .ZN(new_n598_));
  NAND2_X1  g397(.A1(new_n597_), .A2(KEYINPUT35), .ZN(new_n599_));
  XNOR2_X1  g398(.A(new_n599_), .B(KEYINPUT76), .ZN(new_n600_));
  XNOR2_X1  g399(.A(new_n598_), .B(new_n600_), .ZN(new_n601_));
  XOR2_X1   g400(.A(G190gat), .B(G218gat), .Z(new_n602_));
  XNOR2_X1  g401(.A(new_n602_), .B(KEYINPUT77), .ZN(new_n603_));
  XOR2_X1   g402(.A(G134gat), .B(G162gat), .Z(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  INV_X1    g404(.A(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(new_n606_), .A2(KEYINPUT36), .ZN(new_n607_));
  AND2_X1   g406(.A1(new_n601_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(new_n605_), .B(KEYINPUT36), .ZN(new_n609_));
  INV_X1    g408(.A(new_n609_), .ZN(new_n610_));
  NOR2_X1   g409(.A1(new_n601_), .A2(new_n610_), .ZN(new_n611_));
  NOR2_X1   g410(.A1(new_n608_), .A2(new_n611_), .ZN(new_n612_));
  XNOR2_X1  g411(.A(KEYINPUT78), .B(KEYINPUT37), .ZN(new_n613_));
  XNOR2_X1  g412(.A(new_n612_), .B(new_n613_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(G231gat), .A2(G233gat), .ZN(new_n615_));
  XNOR2_X1  g414(.A(new_n465_), .B(new_n615_), .ZN(new_n616_));
  XNOR2_X1  g415(.A(new_n616_), .B(new_n561_), .ZN(new_n617_));
  XOR2_X1   g416(.A(G127gat), .B(G155gat), .Z(new_n618_));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619_));
  XNOR2_X1  g418(.A(new_n618_), .B(new_n619_), .ZN(new_n620_));
  XOR2_X1   g419(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n621_));
  XNOR2_X1  g420(.A(new_n620_), .B(new_n621_), .ZN(new_n622_));
  XNOR2_X1  g421(.A(new_n622_), .B(KEYINPUT17), .ZN(new_n623_));
  OR2_X1    g422(.A1(new_n617_), .A2(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n617_), .A2(KEYINPUT17), .A3(new_n622_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n624_), .A2(new_n625_), .ZN(new_n626_));
  INV_X1    g425(.A(new_n626_), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n614_), .A2(new_n627_), .ZN(new_n628_));
  NOR3_X1   g427(.A1(new_n489_), .A2(new_n594_), .A3(new_n628_), .ZN(new_n629_));
  XOR2_X1   g428(.A(new_n427_), .B(KEYINPUT103), .Z(new_n630_));
  NAND3_X1  g429(.A1(new_n629_), .A2(new_n455_), .A3(new_n630_), .ZN(new_n631_));
  XNOR2_X1  g430(.A(new_n631_), .B(KEYINPUT38), .ZN(new_n632_));
  INV_X1    g431(.A(new_n612_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n453_), .A2(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(new_n634_), .B(KEYINPUT105), .ZN(new_n635_));
  OAI21_X1  g434(.A(new_n485_), .B1(new_n587_), .B2(new_n592_), .ZN(new_n636_));
  INV_X1    g435(.A(KEYINPUT104), .ZN(new_n637_));
  NAND2_X1  g436(.A1(new_n636_), .A2(new_n637_), .ZN(new_n638_));
  OAI211_X1 g437(.A(KEYINPUT104), .B(new_n485_), .C1(new_n587_), .C2(new_n592_), .ZN(new_n639_));
  AND3_X1   g438(.A1(new_n638_), .A2(new_n627_), .A3(new_n639_), .ZN(new_n640_));
  AOI21_X1  g439(.A(KEYINPUT106), .B1(new_n635_), .B2(new_n640_), .ZN(new_n641_));
  INV_X1    g440(.A(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n635_), .A2(KEYINPUT106), .A3(new_n640_), .ZN(new_n643_));
  AOI21_X1  g442(.A(new_n428_), .B1(new_n642_), .B2(new_n643_), .ZN(new_n644_));
  OAI21_X1  g443(.A(new_n632_), .B1(new_n455_), .B2(new_n644_), .ZN(G1324gat));
  NAND2_X1  g444(.A1(new_n376_), .A2(new_n384_), .ZN(new_n646_));
  INV_X1    g445(.A(new_n646_), .ZN(new_n647_));
  NAND3_X1  g446(.A1(new_n629_), .A2(new_n456_), .A3(new_n647_), .ZN(new_n648_));
  NAND3_X1  g447(.A1(new_n635_), .A2(new_n647_), .A3(new_n640_), .ZN(new_n649_));
  INV_X1    g448(.A(KEYINPUT39), .ZN(new_n650_));
  AND3_X1   g449(.A1(new_n649_), .A2(new_n650_), .A3(G8gat), .ZN(new_n651_));
  AOI21_X1  g450(.A(new_n650_), .B1(new_n649_), .B2(G8gat), .ZN(new_n652_));
  OAI21_X1  g451(.A(new_n648_), .B1(new_n651_), .B2(new_n652_), .ZN(new_n653_));
  INV_X1    g452(.A(KEYINPUT40), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n653_), .A2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(KEYINPUT40), .B(new_n648_), .C1(new_n651_), .C2(new_n652_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n655_), .A2(new_n656_), .ZN(G1325gat));
  INV_X1    g456(.A(new_n451_), .ZN(new_n658_));
  NAND3_X1  g457(.A1(new_n629_), .A2(new_n395_), .A3(new_n658_), .ZN(new_n659_));
  INV_X1    g458(.A(new_n643_), .ZN(new_n660_));
  OAI21_X1  g459(.A(new_n658_), .B1(new_n660_), .B2(new_n641_), .ZN(new_n661_));
  AND3_X1   g460(.A1(new_n661_), .A2(KEYINPUT41), .A3(G15gat), .ZN(new_n662_));
  AOI21_X1  g461(.A(KEYINPUT41), .B1(new_n661_), .B2(G15gat), .ZN(new_n663_));
  OAI21_X1  g462(.A(new_n659_), .B1(new_n662_), .B2(new_n663_), .ZN(G1326gat));
  INV_X1    g463(.A(G22gat), .ZN(new_n665_));
  NAND3_X1  g464(.A1(new_n629_), .A2(new_n665_), .A3(new_n273_), .ZN(new_n666_));
  OAI21_X1  g465(.A(new_n273_), .B1(new_n660_), .B2(new_n641_), .ZN(new_n667_));
  INV_X1    g466(.A(KEYINPUT42), .ZN(new_n668_));
  AND3_X1   g467(.A1(new_n667_), .A2(new_n668_), .A3(G22gat), .ZN(new_n669_));
  AOI21_X1  g468(.A(new_n668_), .B1(new_n667_), .B2(G22gat), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(G1327gat));
  NOR2_X1   g470(.A1(new_n633_), .A2(new_n627_), .ZN(new_n672_));
  OAI211_X1 g471(.A(new_n593_), .B(new_n672_), .C1(new_n486_), .C2(new_n488_), .ZN(new_n673_));
  INV_X1    g472(.A(new_n673_), .ZN(new_n674_));
  AOI21_X1  g473(.A(G29gat), .B1(new_n674_), .B2(new_n427_), .ZN(new_n675_));
  NAND3_X1  g474(.A1(new_n638_), .A2(new_n626_), .A3(new_n639_), .ZN(new_n676_));
  NAND2_X1  g475(.A1(new_n676_), .A2(KEYINPUT107), .ZN(new_n677_));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n638_), .A2(new_n678_), .A3(new_n626_), .A4(new_n639_), .ZN(new_n679_));
  OAI21_X1  g478(.A(KEYINPUT43), .B1(new_n452_), .B2(new_n614_), .ZN(new_n680_));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n681_));
  XOR2_X1   g480(.A(new_n612_), .B(new_n613_), .Z(new_n682_));
  AOI211_X1 g481(.A(new_n273_), .B(new_n430_), .C1(new_n376_), .C2(new_n384_), .ZN(new_n683_));
  AOI21_X1  g482(.A(new_n658_), .B1(new_n447_), .B2(new_n449_), .ZN(new_n684_));
  OAI211_X1 g483(.A(new_n681_), .B(new_n682_), .C1(new_n683_), .C2(new_n684_), .ZN(new_n685_));
  AOI22_X1  g484(.A1(new_n677_), .A2(new_n679_), .B1(new_n680_), .B2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n686_), .A2(KEYINPUT44), .ZN(new_n687_));
  INV_X1    g486(.A(G29gat), .ZN(new_n688_));
  INV_X1    g487(.A(new_n630_), .ZN(new_n689_));
  NOR3_X1   g488(.A1(new_n687_), .A2(new_n688_), .A3(new_n689_), .ZN(new_n690_));
  NAND2_X1  g489(.A1(new_n677_), .A2(new_n679_), .ZN(new_n691_));
  NAND2_X1  g490(.A1(new_n680_), .A2(new_n685_), .ZN(new_n692_));
  NAND3_X1  g491(.A1(new_n691_), .A2(KEYINPUT44), .A3(new_n692_), .ZN(new_n693_));
  NAND2_X1  g492(.A1(new_n693_), .A2(KEYINPUT108), .ZN(new_n694_));
  INV_X1    g493(.A(KEYINPUT108), .ZN(new_n695_));
  NAND3_X1  g494(.A1(new_n686_), .A2(new_n695_), .A3(KEYINPUT44), .ZN(new_n696_));
  NAND2_X1  g495(.A1(new_n694_), .A2(new_n696_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n675_), .B1(new_n690_), .B2(new_n697_), .ZN(G1328gat));
  NOR3_X1   g497(.A1(new_n673_), .A2(G36gat), .A3(new_n646_), .ZN(new_n699_));
  XNOR2_X1  g498(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n700_));
  INV_X1    g499(.A(new_n700_), .ZN(new_n701_));
  XNOR2_X1  g500(.A(new_n699_), .B(new_n701_), .ZN(new_n702_));
  AOI21_X1  g501(.A(new_n687_), .B1(new_n694_), .B2(new_n696_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(new_n647_), .ZN(new_n704_));
  INV_X1    g503(.A(G36gat), .ZN(new_n705_));
  OAI211_X1 g504(.A(new_n702_), .B(KEYINPUT46), .C1(new_n704_), .C2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT46), .ZN(new_n707_));
  XNOR2_X1  g506(.A(new_n699_), .B(new_n700_), .ZN(new_n708_));
  AOI21_X1  g507(.A(new_n705_), .B1(new_n703_), .B2(new_n647_), .ZN(new_n709_));
  OAI21_X1  g508(.A(new_n707_), .B1(new_n708_), .B2(new_n709_), .ZN(new_n710_));
  NAND2_X1  g509(.A1(new_n706_), .A2(new_n710_), .ZN(G1329gat));
  INV_X1    g510(.A(G43gat), .ZN(new_n712_));
  OAI21_X1  g511(.A(new_n712_), .B1(new_n673_), .B2(new_n451_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n658_), .A2(G43gat), .ZN(new_n714_));
  NAND2_X1  g513(.A1(new_n691_), .A2(new_n692_), .ZN(new_n715_));
  INV_X1    g514(.A(KEYINPUT44), .ZN(new_n716_));
  AOI21_X1  g515(.A(new_n714_), .B1(new_n715_), .B2(new_n716_), .ZN(new_n717_));
  AND4_X1   g516(.A1(new_n695_), .A2(new_n691_), .A3(KEYINPUT44), .A4(new_n692_), .ZN(new_n718_));
  AOI21_X1  g517(.A(new_n695_), .B1(new_n686_), .B2(KEYINPUT44), .ZN(new_n719_));
  OAI211_X1 g518(.A(KEYINPUT110), .B(new_n717_), .C1(new_n718_), .C2(new_n719_), .ZN(new_n720_));
  INV_X1    g519(.A(new_n720_), .ZN(new_n721_));
  AOI21_X1  g520(.A(KEYINPUT110), .B1(new_n697_), .B2(new_n717_), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n713_), .B1(new_n721_), .B2(new_n722_), .ZN(new_n723_));
  NAND2_X1  g522(.A1(new_n723_), .A2(KEYINPUT47), .ZN(new_n724_));
  INV_X1    g523(.A(KEYINPUT47), .ZN(new_n725_));
  OAI211_X1 g524(.A(new_n725_), .B(new_n713_), .C1(new_n721_), .C2(new_n722_), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n724_), .A2(new_n726_), .ZN(G1330gat));
  AND2_X1   g526(.A1(new_n703_), .A2(new_n273_), .ZN(new_n728_));
  INV_X1    g527(.A(G50gat), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n273_), .A2(new_n729_), .ZN(new_n730_));
  XNOR2_X1  g529(.A(new_n730_), .B(KEYINPUT111), .ZN(new_n731_));
  OAI22_X1  g530(.A1(new_n728_), .A2(new_n729_), .B1(new_n673_), .B2(new_n731_), .ZN(G1331gat));
  NOR4_X1   g531(.A1(new_n452_), .A2(new_n628_), .A3(new_n485_), .A4(new_n593_), .ZN(new_n733_));
  INV_X1    g532(.A(G57gat), .ZN(new_n734_));
  NAND3_X1  g533(.A1(new_n733_), .A2(new_n734_), .A3(new_n630_), .ZN(new_n735_));
  INV_X1    g534(.A(new_n635_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n594_), .A2(new_n487_), .ZN(new_n737_));
  NOR2_X1   g536(.A1(new_n737_), .A2(new_n626_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  NOR3_X1   g538(.A1(new_n736_), .A2(new_n428_), .A3(new_n739_), .ZN(new_n740_));
  OAI21_X1  g539(.A(new_n735_), .B1(new_n740_), .B2(new_n734_), .ZN(G1332gat));
  INV_X1    g540(.A(G64gat), .ZN(new_n742_));
  NAND3_X1  g541(.A1(new_n733_), .A2(new_n742_), .A3(new_n647_), .ZN(new_n743_));
  NOR2_X1   g542(.A1(new_n736_), .A2(new_n739_), .ZN(new_n744_));
  NAND2_X1  g543(.A1(new_n744_), .A2(new_n647_), .ZN(new_n745_));
  XNOR2_X1  g544(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n746_));
  AND3_X1   g545(.A1(new_n745_), .A2(G64gat), .A3(new_n746_), .ZN(new_n747_));
  AOI21_X1  g546(.A(new_n746_), .B1(new_n745_), .B2(G64gat), .ZN(new_n748_));
  OAI21_X1  g547(.A(new_n743_), .B1(new_n747_), .B2(new_n748_), .ZN(G1333gat));
  INV_X1    g548(.A(G71gat), .ZN(new_n750_));
  NAND3_X1  g549(.A1(new_n733_), .A2(new_n750_), .A3(new_n658_), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT49), .ZN(new_n752_));
  NAND2_X1  g551(.A1(new_n744_), .A2(new_n658_), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n752_), .B1(new_n753_), .B2(G71gat), .ZN(new_n754_));
  AOI211_X1 g553(.A(KEYINPUT49), .B(new_n750_), .C1(new_n744_), .C2(new_n658_), .ZN(new_n755_));
  OAI21_X1  g554(.A(new_n751_), .B1(new_n754_), .B2(new_n755_), .ZN(G1334gat));
  NAND3_X1  g555(.A1(new_n733_), .A2(new_n263_), .A3(new_n273_), .ZN(new_n757_));
  NAND3_X1  g556(.A1(new_n635_), .A2(new_n273_), .A3(new_n738_), .ZN(new_n758_));
  INV_X1    g557(.A(KEYINPUT50), .ZN(new_n759_));
  AND3_X1   g558(.A1(new_n758_), .A2(new_n759_), .A3(G78gat), .ZN(new_n760_));
  AOI21_X1  g559(.A(new_n759_), .B1(new_n758_), .B2(G78gat), .ZN(new_n761_));
  OAI21_X1  g560(.A(new_n757_), .B1(new_n760_), .B2(new_n761_), .ZN(new_n762_));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n762_), .A2(new_n763_), .ZN(new_n764_));
  OAI211_X1 g563(.A(KEYINPUT113), .B(new_n757_), .C1(new_n760_), .C2(new_n761_), .ZN(new_n765_));
  NAND2_X1  g564(.A1(new_n764_), .A2(new_n765_), .ZN(G1335gat));
  NOR2_X1   g565(.A1(new_n452_), .A2(new_n485_), .ZN(new_n767_));
  NOR3_X1   g566(.A1(new_n593_), .A2(new_n633_), .A3(new_n627_), .ZN(new_n768_));
  NAND2_X1  g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(new_n769_), .ZN(new_n770_));
  NAND3_X1  g569(.A1(new_n770_), .A2(new_n510_), .A3(new_n630_), .ZN(new_n771_));
  AOI211_X1 g570(.A(new_n627_), .B(new_n737_), .C1(new_n680_), .C2(new_n685_), .ZN(new_n772_));
  AND2_X1   g571(.A1(new_n772_), .A2(new_n427_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n771_), .B1(new_n773_), .B2(new_n510_), .ZN(G1336gat));
  NOR3_X1   g573(.A1(new_n769_), .A2(G92gat), .A3(new_n646_), .ZN(new_n775_));
  NAND2_X1  g574(.A1(new_n772_), .A2(new_n647_), .ZN(new_n776_));
  AOI21_X1  g575(.A(new_n775_), .B1(new_n776_), .B2(G92gat), .ZN(new_n777_));
  XNOR2_X1  g576(.A(new_n777_), .B(KEYINPUT114), .ZN(G1337gat));
  NAND3_X1  g577(.A1(new_n658_), .A2(new_n526_), .A3(new_n528_), .ZN(new_n779_));
  NOR2_X1   g578(.A1(new_n769_), .A2(new_n779_), .ZN(new_n780_));
  XNOR2_X1  g579(.A(new_n780_), .B(KEYINPUT116), .ZN(new_n781_));
  NAND2_X1  g580(.A1(new_n772_), .A2(new_n658_), .ZN(new_n782_));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783_));
  AND3_X1   g582(.A1(new_n782_), .A2(new_n783_), .A3(G99gat), .ZN(new_n784_));
  AOI21_X1  g583(.A(new_n783_), .B1(new_n782_), .B2(G99gat), .ZN(new_n785_));
  OAI21_X1  g584(.A(new_n781_), .B1(new_n784_), .B2(new_n785_), .ZN(new_n786_));
  XNOR2_X1  g585(.A(new_n786_), .B(KEYINPUT51), .ZN(G1338gat));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n788_));
  OAI21_X1  g587(.A(G106gat), .B1(new_n788_), .B2(KEYINPUT118), .ZN(new_n789_));
  AOI21_X1  g588(.A(new_n789_), .B1(new_n772_), .B2(new_n273_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n788_), .A2(KEYINPUT118), .ZN(new_n791_));
  OR2_X1    g590(.A1(new_n790_), .A2(new_n791_), .ZN(new_n792_));
  NOR3_X1   g591(.A1(new_n769_), .A2(G106gat), .A3(new_n432_), .ZN(new_n793_));
  XNOR2_X1  g592(.A(new_n793_), .B(KEYINPUT117), .ZN(new_n794_));
  NAND2_X1  g593(.A1(new_n790_), .A2(new_n791_), .ZN(new_n795_));
  NAND3_X1  g594(.A1(new_n792_), .A2(new_n794_), .A3(new_n795_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g596(.A(KEYINPUT120), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n798_), .A2(KEYINPUT55), .ZN(new_n799_));
  OR2_X1    g598(.A1(new_n578_), .A2(new_n799_), .ZN(new_n800_));
  NAND3_X1  g599(.A1(new_n570_), .A2(new_n575_), .A3(new_n577_), .ZN(new_n801_));
  NAND2_X1  g600(.A1(new_n801_), .A2(new_n556_), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n802_), .A2(KEYINPUT119), .ZN(new_n803_));
  NOR2_X1   g602(.A1(new_n798_), .A2(KEYINPUT55), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n799_), .B1(new_n578_), .B2(new_n804_), .ZN(new_n805_));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n801_), .A2(new_n806_), .A3(new_n556_), .ZN(new_n807_));
  NAND4_X1  g606(.A1(new_n800_), .A2(new_n803_), .A3(new_n805_), .A4(new_n807_), .ZN(new_n808_));
  NAND2_X1  g607(.A1(new_n808_), .A2(new_n497_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n809_), .A2(KEYINPUT56), .ZN(new_n810_));
  INV_X1    g609(.A(new_n472_), .ZN(new_n811_));
  NAND3_X1  g610(.A1(new_n471_), .A2(new_n811_), .A3(new_n474_), .ZN(new_n812_));
  OAI211_X1 g611(.A(new_n482_), .B(new_n812_), .C1(new_n477_), .C2(new_n811_), .ZN(new_n813_));
  AND2_X1   g612(.A1(new_n484_), .A2(new_n813_), .ZN(new_n814_));
  INV_X1    g613(.A(KEYINPUT56), .ZN(new_n815_));
  NAND3_X1  g614(.A1(new_n808_), .A2(new_n815_), .A3(new_n497_), .ZN(new_n816_));
  NAND4_X1  g615(.A1(new_n810_), .A2(new_n814_), .A3(new_n590_), .A4(new_n816_), .ZN(new_n817_));
  INV_X1    g616(.A(KEYINPUT58), .ZN(new_n818_));
  NAND2_X1  g617(.A1(new_n817_), .A2(new_n818_), .ZN(new_n819_));
  NAND2_X1  g618(.A1(new_n682_), .A2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821_));
  NAND2_X1  g620(.A1(new_n820_), .A2(new_n821_), .ZN(new_n822_));
  NAND3_X1  g621(.A1(new_n682_), .A2(new_n819_), .A3(KEYINPUT121), .ZN(new_n823_));
  OR2_X1    g622(.A1(new_n817_), .A2(new_n818_), .ZN(new_n824_));
  NAND3_X1  g623(.A1(new_n822_), .A2(new_n823_), .A3(new_n824_), .ZN(new_n825_));
  NAND2_X1  g624(.A1(new_n590_), .A2(new_n591_), .ZN(new_n826_));
  NAND2_X1  g625(.A1(new_n826_), .A2(new_n814_), .ZN(new_n827_));
  NAND3_X1  g626(.A1(new_n810_), .A2(new_n590_), .A3(new_n816_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n827_), .B1(new_n828_), .B2(new_n487_), .ZN(new_n829_));
  AND3_X1   g628(.A1(new_n829_), .A2(KEYINPUT57), .A3(new_n633_), .ZN(new_n830_));
  AOI21_X1  g629(.A(KEYINPUT57), .B1(new_n829_), .B2(new_n633_), .ZN(new_n831_));
  NOR2_X1   g630(.A1(new_n830_), .A2(new_n831_), .ZN(new_n832_));
  AOI21_X1  g631(.A(new_n627_), .B1(new_n825_), .B2(new_n832_), .ZN(new_n833_));
  NAND4_X1  g632(.A1(new_n593_), .A2(new_n627_), .A3(new_n487_), .A4(new_n614_), .ZN(new_n834_));
  XOR2_X1   g633(.A(new_n834_), .B(KEYINPUT54), .Z(new_n835_));
  NOR2_X1   g634(.A1(new_n833_), .A2(new_n835_), .ZN(new_n836_));
  NAND3_X1  g635(.A1(new_n385_), .A2(new_n658_), .A3(new_n630_), .ZN(new_n837_));
  NOR2_X1   g636(.A1(new_n836_), .A2(new_n837_), .ZN(new_n838_));
  AOI21_X1  g637(.A(G113gat), .B1(new_n838_), .B2(new_n485_), .ZN(new_n839_));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n840_));
  OAI21_X1  g639(.A(new_n840_), .B1(new_n836_), .B2(new_n837_), .ZN(new_n841_));
  INV_X1    g640(.A(new_n837_), .ZN(new_n842_));
  OAI211_X1 g641(.A(KEYINPUT59), .B(new_n842_), .C1(new_n833_), .C2(new_n835_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n841_), .A2(new_n843_), .ZN(new_n844_));
  NOR2_X1   g643(.A1(new_n487_), .A2(KEYINPUT122), .ZN(new_n845_));
  MUX2_X1   g644(.A(KEYINPUT122), .B(new_n845_), .S(G113gat), .Z(new_n846_));
  AOI21_X1  g645(.A(new_n839_), .B1(new_n844_), .B2(new_n846_), .ZN(G1340gat));
  INV_X1    g646(.A(G120gat), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n593_), .B2(KEYINPUT60), .ZN(new_n849_));
  OAI211_X1 g648(.A(new_n838_), .B(new_n849_), .C1(KEYINPUT60), .C2(new_n848_), .ZN(new_n850_));
  AOI21_X1  g649(.A(new_n593_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n851_));
  OAI21_X1  g650(.A(new_n850_), .B1(new_n851_), .B2(new_n848_), .ZN(G1341gat));
  XNOR2_X1  g651(.A(KEYINPUT124), .B(G127gat), .ZN(new_n853_));
  NAND2_X1  g652(.A1(new_n627_), .A2(new_n853_), .ZN(new_n854_));
  AOI21_X1  g653(.A(new_n854_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n855_));
  INV_X1    g654(.A(new_n855_), .ZN(new_n856_));
  INV_X1    g655(.A(KEYINPUT125), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n627_), .B(new_n842_), .C1(new_n833_), .C2(new_n835_), .ZN(new_n858_));
  INV_X1    g657(.A(G127gat), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT123), .B1(new_n858_), .B2(new_n859_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n858_), .A2(KEYINPUT123), .A3(new_n859_), .ZN(new_n861_));
  OAI211_X1 g660(.A(new_n856_), .B(new_n857_), .C1(new_n860_), .C2(new_n861_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n861_), .A2(new_n860_), .ZN(new_n863_));
  OAI21_X1  g662(.A(KEYINPUT125), .B1(new_n863_), .B2(new_n855_), .ZN(new_n864_));
  NAND2_X1  g663(.A1(new_n862_), .A2(new_n864_), .ZN(G1342gat));
  INV_X1    g664(.A(G134gat), .ZN(new_n866_));
  NAND3_X1  g665(.A1(new_n838_), .A2(new_n866_), .A3(new_n612_), .ZN(new_n867_));
  AOI21_X1  g666(.A(new_n614_), .B1(new_n841_), .B2(new_n843_), .ZN(new_n868_));
  OAI21_X1  g667(.A(new_n867_), .B1(new_n868_), .B2(new_n866_), .ZN(G1343gat));
  NOR2_X1   g668(.A1(new_n836_), .A2(new_n658_), .ZN(new_n870_));
  NOR3_X1   g669(.A1(new_n647_), .A2(new_n432_), .A3(new_n689_), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n870_), .A2(new_n485_), .A3(new_n871_), .ZN(new_n872_));
  XNOR2_X1  g671(.A(new_n872_), .B(G141gat), .ZN(G1344gat));
  NAND3_X1  g672(.A1(new_n870_), .A2(new_n594_), .A3(new_n871_), .ZN(new_n874_));
  XNOR2_X1  g673(.A(new_n874_), .B(G148gat), .ZN(G1345gat));
  NAND2_X1  g674(.A1(new_n870_), .A2(new_n871_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n876_), .A2(new_n626_), .ZN(new_n877_));
  XOR2_X1   g676(.A(KEYINPUT61), .B(G155gat), .Z(new_n878_));
  XNOR2_X1  g677(.A(new_n877_), .B(new_n878_), .ZN(G1346gat));
  OAI21_X1  g678(.A(G162gat), .B1(new_n876_), .B2(new_n614_), .ZN(new_n880_));
  OR2_X1    g679(.A1(new_n633_), .A2(G162gat), .ZN(new_n881_));
  OAI21_X1  g680(.A(new_n880_), .B1(new_n876_), .B2(new_n881_), .ZN(G1347gat));
  NAND4_X1  g681(.A1(new_n647_), .A2(new_n432_), .A3(new_n658_), .A4(new_n689_), .ZN(new_n883_));
  NOR2_X1   g682(.A1(new_n836_), .A2(new_n883_), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n884_), .A2(new_n485_), .ZN(new_n885_));
  INV_X1    g684(.A(KEYINPUT126), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n283_), .B1(new_n886_), .B2(KEYINPUT62), .ZN(new_n887_));
  NAND2_X1  g686(.A1(new_n885_), .A2(new_n887_), .ZN(new_n888_));
  INV_X1    g687(.A(KEYINPUT62), .ZN(new_n889_));
  NAND3_X1  g688(.A1(new_n888_), .A2(KEYINPUT126), .A3(new_n889_), .ZN(new_n890_));
  OAI211_X1 g689(.A(new_n885_), .B(new_n887_), .C1(new_n886_), .C2(KEYINPUT62), .ZN(new_n891_));
  NAND3_X1  g690(.A1(new_n884_), .A2(new_n316_), .A3(new_n485_), .ZN(new_n892_));
  NAND3_X1  g691(.A1(new_n890_), .A2(new_n891_), .A3(new_n892_), .ZN(G1348gat));
  NAND2_X1  g692(.A1(new_n884_), .A2(new_n594_), .ZN(new_n894_));
  NOR2_X1   g693(.A1(new_n894_), .A2(new_n284_), .ZN(new_n895_));
  AOI21_X1  g694(.A(new_n895_), .B1(new_n315_), .B2(new_n894_), .ZN(G1349gat));
  NAND2_X1  g695(.A1(new_n884_), .A2(new_n627_), .ZN(new_n897_));
  NOR2_X1   g696(.A1(new_n897_), .A2(new_n278_), .ZN(new_n898_));
  AOI21_X1  g697(.A(new_n898_), .B1(new_n331_), .B2(new_n897_), .ZN(G1350gat));
  NAND3_X1  g698(.A1(new_n884_), .A2(new_n279_), .A3(new_n612_), .ZN(new_n900_));
  NOR3_X1   g699(.A1(new_n836_), .A2(new_n614_), .A3(new_n883_), .ZN(new_n901_));
  INV_X1    g700(.A(G190gat), .ZN(new_n902_));
  OAI21_X1  g701(.A(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(G1351gat));
  NOR3_X1   g702(.A1(new_n646_), .A2(new_n427_), .A3(new_n432_), .ZN(new_n904_));
  NAND2_X1  g703(.A1(new_n870_), .A2(new_n904_), .ZN(new_n905_));
  NOR2_X1   g704(.A1(new_n905_), .A2(new_n487_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(KEYINPUT127), .B(G197gat), .ZN(new_n907_));
  XNOR2_X1  g706(.A(new_n906_), .B(new_n907_), .ZN(G1352gat));
  INV_X1    g707(.A(new_n905_), .ZN(new_n909_));
  AOI21_X1  g708(.A(G204gat), .B1(new_n909_), .B2(new_n594_), .ZN(new_n910_));
  NOR3_X1   g709(.A1(new_n905_), .A2(new_n241_), .A3(new_n593_), .ZN(new_n911_));
  NOR2_X1   g710(.A1(new_n910_), .A2(new_n911_), .ZN(G1353gat));
  XOR2_X1   g711(.A(KEYINPUT63), .B(G211gat), .Z(new_n913_));
  NAND3_X1  g712(.A1(new_n909_), .A2(new_n627_), .A3(new_n913_), .ZN(new_n914_));
  NOR2_X1   g713(.A1(KEYINPUT63), .A2(G211gat), .ZN(new_n915_));
  OAI21_X1  g714(.A(new_n915_), .B1(new_n905_), .B2(new_n626_), .ZN(new_n916_));
  AND2_X1   g715(.A1(new_n914_), .A2(new_n916_), .ZN(G1354gat));
  OR3_X1    g716(.A1(new_n905_), .A2(G218gat), .A3(new_n633_), .ZN(new_n918_));
  OAI21_X1  g717(.A(G218gat), .B1(new_n905_), .B2(new_n614_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n918_), .A2(new_n919_), .ZN(G1355gat));
endmodule


