//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n628_, new_n629_,
    new_n630_, new_n632_, new_n633_, new_n634_, new_n635_, new_n636_,
    new_n637_, new_n638_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n695_, new_n696_, new_n697_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n708_,
    new_n709_, new_n710_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n720_, new_n721_, new_n722_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n736_, new_n737_,
    new_n738_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n834_, new_n835_, new_n836_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n854_, new_n855_, new_n856_, new_n857_,
    new_n859_, new_n861_, new_n862_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n892_,
    new_n893_, new_n895_, new_n896_, new_n897_, new_n899_, new_n900_,
    new_n902_, new_n903_, new_n904_, new_n906_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n915_, new_n916_;
  NAND2_X1  g000(.A1(G183gat), .A2(G190gat), .ZN(new_n202_));
  INV_X1    g001(.A(KEYINPUT82), .ZN(new_n203_));
  XNOR2_X1  g002(.A(new_n202_), .B(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT23), .ZN(new_n205_));
  OAI211_X1 g004(.A(new_n205_), .B(KEYINPUT84), .C1(KEYINPUT23), .C2(new_n202_), .ZN(new_n206_));
  XOR2_X1   g005(.A(KEYINPUT79), .B(G183gat), .Z(new_n207_));
  INV_X1    g006(.A(G190gat), .ZN(new_n208_));
  NAND2_X1  g007(.A1(new_n207_), .A2(new_n208_), .ZN(new_n209_));
  INV_X1    g008(.A(KEYINPUT84), .ZN(new_n210_));
  NAND3_X1  g009(.A1(new_n204_), .A2(new_n210_), .A3(KEYINPUT23), .ZN(new_n211_));
  NAND3_X1  g010(.A1(new_n206_), .A2(new_n209_), .A3(new_n211_), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT85), .ZN(new_n213_));
  NAND2_X1  g012(.A1(new_n212_), .A2(new_n213_), .ZN(new_n214_));
  NAND4_X1  g013(.A1(new_n206_), .A2(KEYINPUT85), .A3(new_n209_), .A4(new_n211_), .ZN(new_n215_));
  NOR2_X1   g014(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n216_));
  XNOR2_X1  g015(.A(new_n216_), .B(G169gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n214_), .A2(new_n215_), .A3(new_n217_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n207_), .A2(KEYINPUT25), .ZN(new_n219_));
  XNOR2_X1  g018(.A(new_n219_), .B(KEYINPUT80), .ZN(new_n220_));
  XOR2_X1   g019(.A(KEYINPUT26), .B(G190gat), .Z(new_n221_));
  INV_X1    g020(.A(KEYINPUT25), .ZN(new_n222_));
  AOI21_X1  g021(.A(new_n221_), .B1(new_n222_), .B2(G183gat), .ZN(new_n223_));
  XOR2_X1   g022(.A(G169gat), .B(G176gat), .Z(new_n224_));
  AOI22_X1  g023(.A1(new_n220_), .A2(new_n223_), .B1(KEYINPUT24), .B2(new_n224_), .ZN(new_n225_));
  NAND2_X1  g024(.A1(new_n202_), .A2(KEYINPUT23), .ZN(new_n226_));
  XNOR2_X1  g025(.A(new_n226_), .B(KEYINPUT81), .ZN(new_n227_));
  OAI21_X1  g026(.A(new_n227_), .B1(KEYINPUT23), .B2(new_n204_), .ZN(new_n228_));
  NOR2_X1   g027(.A1(G169gat), .A2(G176gat), .ZN(new_n229_));
  INV_X1    g028(.A(new_n229_), .ZN(new_n230_));
  OAI21_X1  g029(.A(new_n228_), .B1(KEYINPUT24), .B2(new_n230_), .ZN(new_n231_));
  INV_X1    g030(.A(KEYINPUT83), .ZN(new_n232_));
  NAND2_X1  g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  OAI211_X1 g032(.A(new_n228_), .B(KEYINPUT83), .C1(KEYINPUT24), .C2(new_n230_), .ZN(new_n234_));
  NAND3_X1  g033(.A1(new_n225_), .A2(new_n233_), .A3(new_n234_), .ZN(new_n235_));
  NAND2_X1  g034(.A1(new_n218_), .A2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(KEYINPUT30), .ZN(new_n237_));
  XNOR2_X1  g036(.A(new_n236_), .B(new_n237_), .ZN(new_n238_));
  NAND2_X1  g037(.A1(new_n238_), .A2(KEYINPUT86), .ZN(new_n239_));
  XNOR2_X1  g038(.A(G71gat), .B(G99gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G43gat), .ZN(new_n241_));
  NAND2_X1  g040(.A1(G227gat), .A2(G233gat), .ZN(new_n242_));
  INV_X1    g041(.A(G15gat), .ZN(new_n243_));
  XNOR2_X1  g042(.A(new_n242_), .B(new_n243_), .ZN(new_n244_));
  XNOR2_X1  g043(.A(new_n241_), .B(new_n244_), .ZN(new_n245_));
  NAND2_X1  g044(.A1(new_n239_), .A2(new_n245_), .ZN(new_n246_));
  XNOR2_X1  g045(.A(G127gat), .B(G134gat), .ZN(new_n247_));
  XNOR2_X1  g046(.A(G113gat), .B(G120gat), .ZN(new_n248_));
  XNOR2_X1  g047(.A(new_n247_), .B(new_n248_), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n249_), .A2(KEYINPUT87), .ZN(new_n250_));
  NOR2_X1   g049(.A1(new_n247_), .A2(new_n248_), .ZN(new_n251_));
  OAI21_X1  g050(.A(new_n250_), .B1(KEYINPUT87), .B2(new_n251_), .ZN(new_n252_));
  XOR2_X1   g051(.A(new_n252_), .B(KEYINPUT31), .Z(new_n253_));
  INV_X1    g052(.A(new_n253_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(KEYINPUT88), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n246_), .A2(new_n255_), .ZN(new_n256_));
  XNOR2_X1  g055(.A(new_n236_), .B(KEYINPUT30), .ZN(new_n257_));
  INV_X1    g056(.A(KEYINPUT86), .ZN(new_n258_));
  NAND2_X1  g057(.A1(new_n257_), .A2(new_n258_), .ZN(new_n259_));
  AOI21_X1  g058(.A(new_n245_), .B1(new_n259_), .B2(new_n239_), .ZN(new_n260_));
  NOR2_X1   g059(.A1(new_n254_), .A2(KEYINPUT88), .ZN(new_n261_));
  OR3_X1    g060(.A1(new_n256_), .A2(new_n260_), .A3(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n261_), .B1(new_n256_), .B2(new_n260_), .ZN(new_n263_));
  NAND2_X1  g062(.A1(new_n262_), .A2(new_n263_), .ZN(new_n264_));
  INV_X1    g063(.A(new_n264_), .ZN(new_n265_));
  XNOR2_X1  g064(.A(G8gat), .B(G36gat), .ZN(new_n266_));
  XNOR2_X1  g065(.A(new_n266_), .B(KEYINPUT18), .ZN(new_n267_));
  XNOR2_X1  g066(.A(G64gat), .B(G92gat), .ZN(new_n268_));
  XOR2_X1   g067(.A(new_n267_), .B(new_n268_), .Z(new_n269_));
  NAND2_X1  g068(.A1(G226gat), .A2(G233gat), .ZN(new_n270_));
  XNOR2_X1  g069(.A(new_n270_), .B(KEYINPUT19), .ZN(new_n271_));
  INV_X1    g070(.A(KEYINPUT20), .ZN(new_n272_));
  NOR2_X1   g071(.A1(G197gat), .A2(G204gat), .ZN(new_n273_));
  XNOR2_X1  g072(.A(KEYINPUT91), .B(G197gat), .ZN(new_n274_));
  AOI21_X1  g073(.A(new_n273_), .B1(new_n274_), .B2(G204gat), .ZN(new_n275_));
  XOR2_X1   g074(.A(G211gat), .B(G218gat), .Z(new_n276_));
  NAND3_X1  g075(.A1(new_n275_), .A2(KEYINPUT21), .A3(new_n276_), .ZN(new_n277_));
  INV_X1    g076(.A(KEYINPUT92), .ZN(new_n278_));
  XNOR2_X1  g077(.A(new_n277_), .B(new_n278_), .ZN(new_n279_));
  OR2_X1    g078(.A1(new_n274_), .A2(G204gat), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT21), .ZN(new_n281_));
  AOI21_X1  g080(.A(new_n281_), .B1(G197gat), .B2(G204gat), .ZN(new_n282_));
  AOI21_X1  g081(.A(new_n276_), .B1(new_n280_), .B2(new_n282_), .ZN(new_n283_));
  OAI21_X1  g082(.A(new_n283_), .B1(KEYINPUT21), .B2(new_n275_), .ZN(new_n284_));
  NAND2_X1  g083(.A1(new_n279_), .A2(new_n284_), .ZN(new_n285_));
  AOI21_X1  g084(.A(new_n272_), .B1(new_n236_), .B2(new_n285_), .ZN(new_n286_));
  XNOR2_X1  g085(.A(KEYINPUT25), .B(G183gat), .ZN(new_n287_));
  XNOR2_X1  g086(.A(new_n287_), .B(KEYINPUT96), .ZN(new_n288_));
  OR2_X1    g087(.A1(new_n288_), .A2(new_n221_), .ZN(new_n289_));
  XNOR2_X1  g088(.A(KEYINPUT97), .B(KEYINPUT24), .ZN(new_n290_));
  NOR2_X1   g089(.A1(new_n290_), .A2(new_n230_), .ZN(new_n291_));
  AOI21_X1  g090(.A(new_n291_), .B1(new_n224_), .B2(new_n290_), .ZN(new_n292_));
  NAND4_X1  g091(.A1(new_n289_), .A2(new_n206_), .A3(new_n211_), .A4(new_n292_), .ZN(new_n293_));
  OAI21_X1  g092(.A(new_n228_), .B1(G183gat), .B2(G190gat), .ZN(new_n294_));
  NAND2_X1  g093(.A1(new_n294_), .A2(new_n217_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n293_), .A2(new_n295_), .ZN(new_n296_));
  NOR2_X1   g095(.A1(new_n296_), .A2(new_n285_), .ZN(new_n297_));
  INV_X1    g096(.A(new_n297_), .ZN(new_n298_));
  AOI21_X1  g097(.A(new_n271_), .B1(new_n286_), .B2(new_n298_), .ZN(new_n299_));
  INV_X1    g098(.A(new_n285_), .ZN(new_n300_));
  NAND3_X1  g099(.A1(new_n218_), .A2(new_n300_), .A3(new_n235_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n272_), .B1(new_n296_), .B2(new_n285_), .ZN(new_n302_));
  NAND3_X1  g101(.A1(new_n301_), .A2(new_n302_), .A3(new_n271_), .ZN(new_n303_));
  INV_X1    g102(.A(new_n303_), .ZN(new_n304_));
  OAI21_X1  g103(.A(new_n269_), .B1(new_n299_), .B2(new_n304_), .ZN(new_n305_));
  INV_X1    g104(.A(KEYINPUT98), .ZN(new_n306_));
  INV_X1    g105(.A(new_n269_), .ZN(new_n307_));
  AOI21_X1  g106(.A(new_n300_), .B1(new_n218_), .B2(new_n235_), .ZN(new_n308_));
  NOR3_X1   g107(.A1(new_n308_), .A2(new_n297_), .A3(new_n272_), .ZN(new_n309_));
  OAI211_X1 g108(.A(new_n307_), .B(new_n303_), .C1(new_n309_), .C2(new_n271_), .ZN(new_n310_));
  NAND3_X1  g109(.A1(new_n305_), .A2(new_n306_), .A3(new_n310_), .ZN(new_n311_));
  INV_X1    g110(.A(KEYINPUT27), .ZN(new_n312_));
  NOR2_X1   g111(.A1(new_n299_), .A2(new_n304_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n313_), .A2(KEYINPUT98), .A3(new_n307_), .ZN(new_n314_));
  NAND3_X1  g113(.A1(new_n311_), .A2(new_n312_), .A3(new_n314_), .ZN(new_n315_));
  INV_X1    g114(.A(new_n315_), .ZN(new_n316_));
  XOR2_X1   g115(.A(new_n269_), .B(KEYINPUT103), .Z(new_n317_));
  INV_X1    g116(.A(new_n317_), .ZN(new_n318_));
  NAND2_X1  g117(.A1(new_n301_), .A2(new_n302_), .ZN(new_n319_));
  NOR2_X1   g118(.A1(new_n319_), .A2(new_n271_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(new_n296_), .A2(KEYINPUT100), .ZN(new_n321_));
  INV_X1    g120(.A(KEYINPUT100), .ZN(new_n322_));
  NAND3_X1  g121(.A1(new_n293_), .A2(new_n295_), .A3(new_n322_), .ZN(new_n323_));
  NAND3_X1  g122(.A1(new_n321_), .A2(new_n323_), .A3(new_n300_), .ZN(new_n324_));
  NAND2_X1  g123(.A1(new_n286_), .A2(new_n324_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n325_), .A2(new_n271_), .ZN(new_n326_));
  AOI21_X1  g125(.A(new_n320_), .B1(new_n326_), .B2(KEYINPUT101), .ZN(new_n327_));
  INV_X1    g126(.A(new_n271_), .ZN(new_n328_));
  AOI211_X1 g127(.A(KEYINPUT101), .B(new_n328_), .C1(new_n286_), .C2(new_n324_), .ZN(new_n329_));
  INV_X1    g128(.A(new_n329_), .ZN(new_n330_));
  AOI21_X1  g129(.A(new_n318_), .B1(new_n327_), .B2(new_n330_), .ZN(new_n331_));
  OAI21_X1  g130(.A(new_n303_), .B1(new_n309_), .B2(new_n271_), .ZN(new_n332_));
  AOI21_X1  g131(.A(new_n312_), .B1(new_n332_), .B2(new_n269_), .ZN(new_n333_));
  INV_X1    g132(.A(new_n333_), .ZN(new_n334_));
  OAI21_X1  g133(.A(KEYINPUT104), .B1(new_n331_), .B2(new_n334_), .ZN(new_n335_));
  AOI21_X1  g134(.A(new_n328_), .B1(new_n286_), .B2(new_n324_), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT101), .ZN(new_n337_));
  OAI22_X1  g136(.A1(new_n336_), .A2(new_n337_), .B1(new_n271_), .B2(new_n319_), .ZN(new_n338_));
  OAI21_X1  g137(.A(new_n317_), .B1(new_n338_), .B2(new_n329_), .ZN(new_n339_));
  INV_X1    g138(.A(KEYINPUT104), .ZN(new_n340_));
  NAND3_X1  g139(.A1(new_n339_), .A2(new_n333_), .A3(new_n340_), .ZN(new_n341_));
  AOI21_X1  g140(.A(new_n316_), .B1(new_n335_), .B2(new_n341_), .ZN(new_n342_));
  NAND3_X1  g141(.A1(KEYINPUT93), .A2(G228gat), .A3(G233gat), .ZN(new_n343_));
  XOR2_X1   g142(.A(G155gat), .B(G162gat), .Z(new_n344_));
  OR3_X1    g143(.A1(KEYINPUT3), .A2(G141gat), .A3(G148gat), .ZN(new_n345_));
  OAI21_X1  g144(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n346_));
  NAND2_X1  g145(.A1(G141gat), .A2(G148gat), .ZN(new_n347_));
  INV_X1    g146(.A(KEYINPUT89), .ZN(new_n348_));
  NAND2_X1  g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  OAI211_X1 g148(.A(new_n345_), .B(new_n346_), .C1(new_n349_), .C2(KEYINPUT2), .ZN(new_n350_));
  AND2_X1   g149(.A1(new_n349_), .A2(KEYINPUT2), .ZN(new_n351_));
  OAI21_X1  g150(.A(new_n344_), .B1(new_n350_), .B2(new_n351_), .ZN(new_n352_));
  INV_X1    g151(.A(KEYINPUT1), .ZN(new_n353_));
  NAND2_X1  g152(.A1(new_n344_), .A2(new_n353_), .ZN(new_n354_));
  INV_X1    g153(.A(G141gat), .ZN(new_n355_));
  INV_X1    g154(.A(G148gat), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n355_), .A2(new_n356_), .ZN(new_n357_));
  NAND3_X1  g156(.A1(KEYINPUT1), .A2(G155gat), .A3(G162gat), .ZN(new_n358_));
  NAND4_X1  g157(.A1(new_n354_), .A2(new_n347_), .A3(new_n357_), .A4(new_n358_), .ZN(new_n359_));
  AND2_X1   g158(.A1(new_n352_), .A2(new_n359_), .ZN(new_n360_));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361_));
  OAI21_X1  g160(.A(new_n343_), .B1(new_n360_), .B2(new_n361_), .ZN(new_n362_));
  NOR2_X1   g161(.A1(new_n300_), .A2(new_n362_), .ZN(new_n363_));
  XNOR2_X1  g162(.A(new_n363_), .B(KEYINPUT95), .ZN(new_n364_));
  INV_X1    g163(.A(new_n364_), .ZN(new_n365_));
  NAND2_X1  g164(.A1(new_n360_), .A2(new_n361_), .ZN(new_n366_));
  XNOR2_X1  g165(.A(KEYINPUT90), .B(KEYINPUT28), .ZN(new_n367_));
  XNOR2_X1  g166(.A(new_n366_), .B(new_n367_), .ZN(new_n368_));
  XOR2_X1   g167(.A(G22gat), .B(G50gat), .Z(new_n369_));
  AOI21_X1  g168(.A(KEYINPUT93), .B1(G228gat), .B2(G233gat), .ZN(new_n370_));
  XNOR2_X1  g169(.A(new_n369_), .B(new_n370_), .ZN(new_n371_));
  OR2_X1    g170(.A1(new_n368_), .A2(new_n371_), .ZN(new_n372_));
  NAND2_X1  g171(.A1(new_n368_), .A2(new_n371_), .ZN(new_n373_));
  XNOR2_X1  g172(.A(G78gat), .B(G106gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(new_n374_), .B(KEYINPUT94), .ZN(new_n375_));
  INV_X1    g174(.A(new_n375_), .ZN(new_n376_));
  NAND3_X1  g175(.A1(new_n372_), .A2(new_n373_), .A3(new_n376_), .ZN(new_n377_));
  INV_X1    g176(.A(new_n377_), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n376_), .B1(new_n372_), .B2(new_n373_), .ZN(new_n379_));
  OAI21_X1  g178(.A(new_n365_), .B1(new_n378_), .B2(new_n379_), .ZN(new_n380_));
  NAND2_X1  g179(.A1(new_n372_), .A2(new_n373_), .ZN(new_n381_));
  NAND2_X1  g180(.A1(new_n381_), .A2(new_n375_), .ZN(new_n382_));
  NAND3_X1  g181(.A1(new_n382_), .A2(new_n364_), .A3(new_n377_), .ZN(new_n383_));
  AND2_X1   g182(.A1(new_n380_), .A2(new_n383_), .ZN(new_n384_));
  OR2_X1    g183(.A1(new_n252_), .A2(new_n360_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n360_), .A2(new_n249_), .ZN(new_n386_));
  NAND3_X1  g185(.A1(new_n385_), .A2(KEYINPUT4), .A3(new_n386_), .ZN(new_n387_));
  NAND2_X1  g186(.A1(G225gat), .A2(G233gat), .ZN(new_n388_));
  NOR2_X1   g187(.A1(new_n252_), .A2(new_n360_), .ZN(new_n389_));
  INV_X1    g188(.A(KEYINPUT4), .ZN(new_n390_));
  AOI21_X1  g189(.A(new_n388_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n391_));
  NAND3_X1  g190(.A1(new_n387_), .A2(KEYINPUT99), .A3(new_n391_), .ZN(new_n392_));
  NAND3_X1  g191(.A1(new_n385_), .A2(new_n386_), .A3(new_n388_), .ZN(new_n393_));
  NAND2_X1  g192(.A1(new_n392_), .A2(new_n393_), .ZN(new_n394_));
  AOI21_X1  g193(.A(KEYINPUT99), .B1(new_n387_), .B2(new_n391_), .ZN(new_n395_));
  NOR2_X1   g194(.A1(new_n394_), .A2(new_n395_), .ZN(new_n396_));
  XNOR2_X1  g195(.A(G1gat), .B(G29gat), .ZN(new_n397_));
  XNOR2_X1  g196(.A(new_n397_), .B(G85gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(KEYINPUT0), .B(G57gat), .ZN(new_n399_));
  XOR2_X1   g198(.A(new_n398_), .B(new_n399_), .Z(new_n400_));
  NAND3_X1  g199(.A1(new_n396_), .A2(KEYINPUT102), .A3(new_n400_), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n387_), .A2(new_n391_), .ZN(new_n402_));
  INV_X1    g201(.A(KEYINPUT99), .ZN(new_n403_));
  NAND2_X1  g202(.A1(new_n402_), .A2(new_n403_), .ZN(new_n404_));
  NAND4_X1  g203(.A1(new_n404_), .A2(new_n400_), .A3(new_n393_), .A4(new_n392_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT102), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  INV_X1    g206(.A(new_n400_), .ZN(new_n408_));
  OAI21_X1  g207(.A(new_n408_), .B1(new_n394_), .B2(new_n395_), .ZN(new_n409_));
  NAND3_X1  g208(.A1(new_n401_), .A2(new_n407_), .A3(new_n409_), .ZN(new_n410_));
  INV_X1    g209(.A(new_n410_), .ZN(new_n411_));
  NAND4_X1  g210(.A1(new_n265_), .A2(new_n342_), .A3(new_n384_), .A4(new_n411_), .ZN(new_n412_));
  NOR2_X1   g211(.A1(new_n384_), .A2(new_n410_), .ZN(new_n413_));
  NAND2_X1  g212(.A1(new_n269_), .A2(KEYINPUT32), .ZN(new_n414_));
  INV_X1    g213(.A(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n415_), .B1(new_n338_), .B2(new_n329_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n332_), .A2(new_n414_), .ZN(new_n417_));
  NAND3_X1  g216(.A1(new_n416_), .A2(new_n410_), .A3(new_n417_), .ZN(new_n418_));
  AND2_X1   g217(.A1(new_n311_), .A2(new_n314_), .ZN(new_n419_));
  NAND3_X1  g218(.A1(new_n396_), .A2(KEYINPUT33), .A3(new_n400_), .ZN(new_n420_));
  NAND2_X1  g219(.A1(new_n385_), .A2(new_n386_), .ZN(new_n421_));
  INV_X1    g220(.A(new_n387_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n388_), .B1(new_n385_), .B2(KEYINPUT4), .ZN(new_n423_));
  OAI221_X1 g222(.A(new_n408_), .B1(new_n421_), .B2(new_n388_), .C1(new_n422_), .C2(new_n423_), .ZN(new_n424_));
  INV_X1    g223(.A(KEYINPUT33), .ZN(new_n425_));
  NAND2_X1  g224(.A1(new_n405_), .A2(new_n425_), .ZN(new_n426_));
  NAND3_X1  g225(.A1(new_n420_), .A2(new_n424_), .A3(new_n426_), .ZN(new_n427_));
  OAI21_X1  g226(.A(new_n418_), .B1(new_n419_), .B2(new_n427_), .ZN(new_n428_));
  AOI22_X1  g227(.A1(new_n342_), .A2(new_n413_), .B1(new_n428_), .B2(new_n384_), .ZN(new_n429_));
  OAI21_X1  g228(.A(new_n412_), .B1(new_n429_), .B2(new_n265_), .ZN(new_n430_));
  XOR2_X1   g229(.A(G29gat), .B(G36gat), .Z(new_n431_));
  XOR2_X1   g230(.A(G43gat), .B(G50gat), .Z(new_n432_));
  XOR2_X1   g231(.A(new_n431_), .B(new_n432_), .Z(new_n433_));
  XOR2_X1   g232(.A(new_n433_), .B(KEYINPUT15), .Z(new_n434_));
  INV_X1    g233(.A(KEYINPUT14), .ZN(new_n435_));
  XOR2_X1   g234(.A(KEYINPUT76), .B(G8gat), .Z(new_n436_));
  XNOR2_X1  g235(.A(KEYINPUT75), .B(G1gat), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n435_), .B1(new_n436_), .B2(new_n437_), .ZN(new_n438_));
  XOR2_X1   g237(.A(G15gat), .B(G22gat), .Z(new_n439_));
  XNOR2_X1  g238(.A(G1gat), .B(G8gat), .ZN(new_n440_));
  INV_X1    g239(.A(new_n440_), .ZN(new_n441_));
  OR3_X1    g240(.A1(new_n438_), .A2(new_n439_), .A3(new_n441_), .ZN(new_n442_));
  OAI21_X1  g241(.A(new_n441_), .B1(new_n438_), .B2(new_n439_), .ZN(new_n443_));
  NAND2_X1  g242(.A1(new_n442_), .A2(new_n443_), .ZN(new_n444_));
  INV_X1    g243(.A(new_n444_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n434_), .A2(new_n445_), .ZN(new_n446_));
  NAND2_X1  g245(.A1(G229gat), .A2(G233gat), .ZN(new_n447_));
  INV_X1    g246(.A(new_n433_), .ZN(new_n448_));
  NAND2_X1  g247(.A1(new_n444_), .A2(new_n448_), .ZN(new_n449_));
  NAND3_X1  g248(.A1(new_n446_), .A2(new_n447_), .A3(new_n449_), .ZN(new_n450_));
  XNOR2_X1  g249(.A(new_n444_), .B(new_n448_), .ZN(new_n451_));
  NAND3_X1  g250(.A1(new_n451_), .A2(G229gat), .A3(G233gat), .ZN(new_n452_));
  AND2_X1   g251(.A1(new_n450_), .A2(new_n452_), .ZN(new_n453_));
  XOR2_X1   g252(.A(G113gat), .B(G141gat), .Z(new_n454_));
  XNOR2_X1  g253(.A(G169gat), .B(G197gat), .ZN(new_n455_));
  XNOR2_X1  g254(.A(new_n454_), .B(new_n455_), .ZN(new_n456_));
  NAND2_X1  g255(.A1(new_n453_), .A2(new_n456_), .ZN(new_n457_));
  NAND2_X1  g256(.A1(new_n457_), .A2(KEYINPUT78), .ZN(new_n458_));
  INV_X1    g257(.A(KEYINPUT78), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n453_), .A2(new_n459_), .A3(new_n456_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n458_), .A2(new_n460_), .ZN(new_n461_));
  OR2_X1    g260(.A1(new_n453_), .A2(new_n456_), .ZN(new_n462_));
  NAND2_X1  g261(.A1(new_n461_), .A2(new_n462_), .ZN(new_n463_));
  AND2_X1   g262(.A1(new_n430_), .A2(new_n463_), .ZN(new_n464_));
  XNOR2_X1  g263(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n465_));
  INV_X1    g264(.A(new_n465_), .ZN(new_n466_));
  XOR2_X1   g265(.A(KEYINPUT71), .B(KEYINPUT12), .Z(new_n467_));
  XNOR2_X1  g266(.A(KEYINPUT10), .B(G99gat), .ZN(new_n468_));
  XNOR2_X1  g267(.A(new_n468_), .B(KEYINPUT64), .ZN(new_n469_));
  INV_X1    g268(.A(G106gat), .ZN(new_n470_));
  AND2_X1   g269(.A1(new_n469_), .A2(new_n470_), .ZN(new_n471_));
  XNOR2_X1  g270(.A(KEYINPUT65), .B(G85gat), .ZN(new_n472_));
  INV_X1    g271(.A(KEYINPUT9), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(new_n473_), .A3(G92gat), .ZN(new_n474_));
  NAND2_X1  g273(.A1(G99gat), .A2(G106gat), .ZN(new_n475_));
  XNOR2_X1  g274(.A(new_n475_), .B(KEYINPUT6), .ZN(new_n476_));
  XOR2_X1   g275(.A(G85gat), .B(G92gat), .Z(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  OAI211_X1 g277(.A(new_n474_), .B(new_n476_), .C1(new_n473_), .C2(new_n478_), .ZN(new_n479_));
  NOR2_X1   g278(.A1(new_n471_), .A2(new_n479_), .ZN(new_n480_));
  INV_X1    g279(.A(KEYINPUT7), .ZN(new_n481_));
  INV_X1    g280(.A(G99gat), .ZN(new_n482_));
  NAND3_X1  g281(.A1(new_n481_), .A2(new_n482_), .A3(new_n470_), .ZN(new_n483_));
  OAI21_X1  g282(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n484_));
  NAND2_X1  g283(.A1(new_n483_), .A2(new_n484_), .ZN(new_n485_));
  INV_X1    g284(.A(new_n485_), .ZN(new_n486_));
  NAND2_X1  g285(.A1(new_n486_), .A2(new_n476_), .ZN(new_n487_));
  INV_X1    g286(.A(KEYINPUT8), .ZN(new_n488_));
  AND3_X1   g287(.A1(new_n487_), .A2(new_n488_), .A3(new_n477_), .ZN(new_n489_));
  INV_X1    g288(.A(KEYINPUT6), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(KEYINPUT66), .ZN(new_n491_));
  INV_X1    g290(.A(KEYINPUT66), .ZN(new_n492_));
  NAND2_X1  g291(.A1(new_n492_), .A2(KEYINPUT6), .ZN(new_n493_));
  AND3_X1   g292(.A1(new_n491_), .A2(new_n493_), .A3(new_n475_), .ZN(new_n494_));
  AOI21_X1  g293(.A(new_n475_), .B1(new_n491_), .B2(new_n493_), .ZN(new_n495_));
  NOR3_X1   g294(.A1(new_n494_), .A2(new_n495_), .A3(new_n485_), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT67), .B1(new_n496_), .B2(new_n478_), .ZN(new_n497_));
  INV_X1    g296(.A(KEYINPUT67), .ZN(new_n498_));
  XNOR2_X1  g297(.A(KEYINPUT66), .B(KEYINPUT6), .ZN(new_n499_));
  OAI211_X1 g298(.A(new_n483_), .B(new_n484_), .C1(new_n499_), .C2(new_n475_), .ZN(new_n500_));
  OAI211_X1 g299(.A(new_n498_), .B(new_n477_), .C1(new_n500_), .C2(new_n494_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n497_), .A2(KEYINPUT8), .A3(new_n501_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n489_), .B1(new_n502_), .B2(KEYINPUT68), .ZN(new_n503_));
  INV_X1    g302(.A(KEYINPUT68), .ZN(new_n504_));
  NAND4_X1  g303(.A1(new_n497_), .A2(new_n504_), .A3(KEYINPUT8), .A4(new_n501_), .ZN(new_n505_));
  AOI21_X1  g304(.A(new_n480_), .B1(new_n503_), .B2(new_n505_), .ZN(new_n506_));
  XNOR2_X1  g305(.A(G57gat), .B(G64gat), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n507_), .A2(KEYINPUT11), .ZN(new_n508_));
  XOR2_X1   g307(.A(G71gat), .B(G78gat), .Z(new_n509_));
  OR2_X1    g308(.A1(new_n508_), .A2(new_n509_), .ZN(new_n510_));
  NOR2_X1   g309(.A1(new_n507_), .A2(KEYINPUT11), .ZN(new_n511_));
  NAND2_X1  g310(.A1(new_n508_), .A2(new_n509_), .ZN(new_n512_));
  OAI21_X1  g311(.A(new_n510_), .B1(new_n511_), .B2(new_n512_), .ZN(new_n513_));
  XOR2_X1   g312(.A(new_n513_), .B(KEYINPUT69), .Z(new_n514_));
  OAI21_X1  g313(.A(new_n467_), .B1(new_n506_), .B2(new_n514_), .ZN(new_n515_));
  NAND2_X1  g314(.A1(G230gat), .A2(G233gat), .ZN(new_n516_));
  NAND2_X1  g315(.A1(new_n501_), .A2(KEYINPUT8), .ZN(new_n517_));
  NOR2_X1   g316(.A1(new_n495_), .A2(new_n485_), .ZN(new_n518_));
  INV_X1    g317(.A(new_n494_), .ZN(new_n519_));
  NAND2_X1  g318(.A1(new_n518_), .A2(new_n519_), .ZN(new_n520_));
  AOI21_X1  g319(.A(new_n498_), .B1(new_n520_), .B2(new_n477_), .ZN(new_n521_));
  OAI21_X1  g320(.A(KEYINPUT68), .B1(new_n517_), .B2(new_n521_), .ZN(new_n522_));
  INV_X1    g321(.A(new_n489_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n522_), .A2(new_n505_), .A3(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(new_n480_), .ZN(new_n525_));
  NAND3_X1  g324(.A1(new_n524_), .A2(new_n514_), .A3(new_n525_), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n524_), .A2(new_n525_), .ZN(new_n527_));
  INV_X1    g326(.A(KEYINPUT12), .ZN(new_n528_));
  OR2_X1    g327(.A1(new_n513_), .A2(new_n528_), .ZN(new_n529_));
  INV_X1    g328(.A(new_n529_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n527_), .A2(new_n530_), .ZN(new_n531_));
  NAND4_X1  g330(.A1(new_n515_), .A2(new_n516_), .A3(new_n526_), .A4(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(new_n516_), .ZN(new_n533_));
  AND3_X1   g332(.A1(new_n524_), .A2(new_n514_), .A3(new_n525_), .ZN(new_n534_));
  AOI21_X1  g333(.A(new_n514_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n535_));
  OAI21_X1  g334(.A(new_n533_), .B1(new_n534_), .B2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(new_n532_), .A2(KEYINPUT70), .A3(new_n536_), .ZN(new_n537_));
  OR2_X1    g336(.A1(new_n536_), .A2(KEYINPUT70), .ZN(new_n538_));
  XNOR2_X1  g337(.A(G120gat), .B(G148gat), .ZN(new_n539_));
  XNOR2_X1  g338(.A(new_n539_), .B(KEYINPUT5), .ZN(new_n540_));
  XNOR2_X1  g339(.A(G176gat), .B(G204gat), .ZN(new_n541_));
  XOR2_X1   g340(.A(new_n540_), .B(new_n541_), .Z(new_n542_));
  NAND3_X1  g341(.A1(new_n537_), .A2(new_n538_), .A3(new_n542_), .ZN(new_n543_));
  INV_X1    g342(.A(new_n543_), .ZN(new_n544_));
  AOI21_X1  g343(.A(new_n542_), .B1(new_n537_), .B2(new_n538_), .ZN(new_n545_));
  OAI21_X1  g344(.A(new_n466_), .B1(new_n544_), .B2(new_n545_), .ZN(new_n546_));
  INV_X1    g345(.A(new_n545_), .ZN(new_n547_));
  NAND2_X1  g346(.A1(new_n547_), .A2(new_n543_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT13), .ZN(new_n549_));
  NOR2_X1   g348(.A1(new_n549_), .A2(KEYINPUT72), .ZN(new_n550_));
  OAI21_X1  g349(.A(new_n546_), .B1(new_n548_), .B2(new_n550_), .ZN(new_n551_));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552_));
  XOR2_X1   g351(.A(new_n444_), .B(new_n552_), .Z(new_n553_));
  XNOR2_X1  g352(.A(new_n553_), .B(new_n514_), .ZN(new_n554_));
  XOR2_X1   g353(.A(G127gat), .B(G155gat), .Z(new_n555_));
  XNOR2_X1  g354(.A(new_n555_), .B(KEYINPUT16), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G183gat), .B(G211gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n556_), .B(new_n557_), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(KEYINPUT17), .ZN(new_n559_));
  NAND2_X1  g358(.A1(new_n554_), .A2(new_n559_), .ZN(new_n560_));
  XNOR2_X1  g359(.A(new_n560_), .B(KEYINPUT77), .ZN(new_n561_));
  AND2_X1   g360(.A1(new_n553_), .A2(new_n513_), .ZN(new_n562_));
  INV_X1    g361(.A(KEYINPUT17), .ZN(new_n563_));
  NOR3_X1   g362(.A1(new_n562_), .A2(new_n563_), .A3(new_n558_), .ZN(new_n564_));
  OAI21_X1  g363(.A(new_n564_), .B1(new_n513_), .B2(new_n553_), .ZN(new_n565_));
  NAND2_X1  g364(.A1(new_n561_), .A2(new_n565_), .ZN(new_n566_));
  INV_X1    g365(.A(new_n566_), .ZN(new_n567_));
  XOR2_X1   g366(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n568_));
  NAND2_X1  g367(.A1(G232gat), .A2(G233gat), .ZN(new_n569_));
  XNOR2_X1  g368(.A(new_n568_), .B(new_n569_), .ZN(new_n570_));
  INV_X1    g369(.A(new_n434_), .ZN(new_n571_));
  NOR2_X1   g370(.A1(new_n506_), .A2(new_n571_), .ZN(new_n572_));
  NOR2_X1   g371(.A1(new_n527_), .A2(new_n433_), .ZN(new_n573_));
  OAI211_X1 g372(.A(KEYINPUT35), .B(new_n570_), .C1(new_n572_), .C2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n506_), .A2(new_n448_), .ZN(new_n575_));
  NAND2_X1  g374(.A1(new_n527_), .A2(new_n434_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n570_), .A2(KEYINPUT35), .ZN(new_n577_));
  OR2_X1    g376(.A1(new_n570_), .A2(KEYINPUT35), .ZN(new_n578_));
  NAND4_X1  g377(.A1(new_n575_), .A2(new_n576_), .A3(new_n577_), .A4(new_n578_), .ZN(new_n579_));
  NAND2_X1  g378(.A1(new_n574_), .A2(new_n579_), .ZN(new_n580_));
  XNOR2_X1  g379(.A(G190gat), .B(G218gat), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G134gat), .B(G162gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(new_n581_), .B(new_n582_), .ZN(new_n583_));
  XOR2_X1   g382(.A(new_n583_), .B(KEYINPUT36), .Z(new_n584_));
  NAND2_X1  g383(.A1(new_n580_), .A2(new_n584_), .ZN(new_n585_));
  NOR2_X1   g384(.A1(new_n583_), .A2(KEYINPUT36), .ZN(new_n586_));
  NAND3_X1  g385(.A1(new_n574_), .A2(new_n579_), .A3(new_n586_), .ZN(new_n587_));
  NAND3_X1  g386(.A1(new_n585_), .A2(KEYINPUT37), .A3(new_n587_), .ZN(new_n588_));
  INV_X1    g387(.A(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT74), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n585_), .A2(new_n590_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n580_), .A2(KEYINPUT74), .A3(new_n584_), .ZN(new_n592_));
  NAND3_X1  g391(.A1(new_n591_), .A2(new_n587_), .A3(new_n592_), .ZN(new_n593_));
  INV_X1    g392(.A(KEYINPUT37), .ZN(new_n594_));
  AOI21_X1  g393(.A(new_n589_), .B1(new_n593_), .B2(new_n594_), .ZN(new_n595_));
  NAND4_X1  g394(.A1(new_n464_), .A2(new_n551_), .A3(new_n567_), .A4(new_n595_), .ZN(new_n596_));
  OR3_X1    g395(.A1(new_n596_), .A2(new_n437_), .A3(new_n411_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT38), .ZN(new_n598_));
  OR2_X1    g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  AND2_X1   g398(.A1(new_n430_), .A2(new_n593_), .ZN(new_n600_));
  INV_X1    g399(.A(new_n551_), .ZN(new_n601_));
  INV_X1    g400(.A(new_n463_), .ZN(new_n602_));
  NOR2_X1   g401(.A1(new_n601_), .A2(new_n602_), .ZN(new_n603_));
  NAND3_X1  g402(.A1(new_n603_), .A2(KEYINPUT105), .A3(new_n567_), .ZN(new_n604_));
  INV_X1    g403(.A(KEYINPUT105), .ZN(new_n605_));
  INV_X1    g404(.A(new_n603_), .ZN(new_n606_));
  OAI21_X1  g405(.A(new_n605_), .B1(new_n606_), .B2(new_n566_), .ZN(new_n607_));
  AND3_X1   g406(.A1(new_n600_), .A2(new_n604_), .A3(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n608_), .ZN(new_n609_));
  OAI21_X1  g408(.A(G1gat), .B1(new_n609_), .B2(new_n411_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n597_), .A2(new_n598_), .ZN(new_n611_));
  NAND3_X1  g410(.A1(new_n599_), .A2(new_n610_), .A3(new_n611_), .ZN(G1324gat));
  XNOR2_X1  g411(.A(KEYINPUT106), .B(KEYINPUT40), .ZN(new_n613_));
  INV_X1    g412(.A(new_n342_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n608_), .A2(new_n614_), .ZN(new_n615_));
  NAND2_X1  g414(.A1(new_n615_), .A2(G8gat), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n616_), .A2(KEYINPUT39), .ZN(new_n617_));
  INV_X1    g416(.A(KEYINPUT39), .ZN(new_n618_));
  NAND3_X1  g417(.A1(new_n615_), .A2(new_n618_), .A3(G8gat), .ZN(new_n619_));
  NAND2_X1  g418(.A1(new_n617_), .A2(new_n619_), .ZN(new_n620_));
  OR3_X1    g419(.A1(new_n596_), .A2(new_n436_), .A3(new_n342_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n613_), .B1(new_n620_), .B2(new_n621_), .ZN(new_n622_));
  AND3_X1   g421(.A1(new_n615_), .A2(new_n618_), .A3(G8gat), .ZN(new_n623_));
  AOI21_X1  g422(.A(new_n618_), .B1(new_n615_), .B2(G8gat), .ZN(new_n624_));
  OAI211_X1 g423(.A(new_n621_), .B(new_n613_), .C1(new_n623_), .C2(new_n624_), .ZN(new_n625_));
  INV_X1    g424(.A(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n622_), .A2(new_n626_), .ZN(G1325gat));
  AOI21_X1  g426(.A(new_n243_), .B1(new_n608_), .B2(new_n265_), .ZN(new_n628_));
  XNOR2_X1  g427(.A(new_n628_), .B(KEYINPUT41), .ZN(new_n629_));
  NAND2_X1  g428(.A1(new_n265_), .A2(new_n243_), .ZN(new_n630_));
  OAI21_X1  g429(.A(new_n629_), .B1(new_n596_), .B2(new_n630_), .ZN(G1326gat));
  OR3_X1    g430(.A1(new_n596_), .A2(G22gat), .A3(new_n384_), .ZN(new_n632_));
  INV_X1    g431(.A(new_n384_), .ZN(new_n633_));
  NAND2_X1  g432(.A1(new_n608_), .A2(new_n633_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT42), .ZN(new_n635_));
  AND3_X1   g434(.A1(new_n634_), .A2(new_n635_), .A3(G22gat), .ZN(new_n636_));
  AOI21_X1  g435(.A(new_n635_), .B1(new_n634_), .B2(G22gat), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n632_), .B1(new_n636_), .B2(new_n637_), .ZN(new_n638_));
  XNOR2_X1  g437(.A(new_n638_), .B(KEYINPUT107), .ZN(G1327gat));
  INV_X1    g438(.A(new_n593_), .ZN(new_n640_));
  NAND2_X1  g439(.A1(new_n640_), .A2(new_n566_), .ZN(new_n641_));
  NOR2_X1   g440(.A1(new_n601_), .A2(new_n641_), .ZN(new_n642_));
  NAND3_X1  g441(.A1(new_n430_), .A2(new_n642_), .A3(new_n463_), .ZN(new_n643_));
  OR3_X1    g442(.A1(new_n643_), .A2(G29gat), .A3(new_n411_), .ZN(new_n644_));
  INV_X1    g443(.A(new_n595_), .ZN(new_n645_));
  NAND2_X1  g444(.A1(new_n645_), .A2(KEYINPUT108), .ZN(new_n646_));
  INV_X1    g445(.A(KEYINPUT108), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n595_), .A2(new_n647_), .ZN(new_n648_));
  AND3_X1   g447(.A1(new_n339_), .A2(new_n333_), .A3(new_n340_), .ZN(new_n649_));
  AOI21_X1  g448(.A(new_n340_), .B1(new_n339_), .B2(new_n333_), .ZN(new_n650_));
  OAI211_X1 g449(.A(new_n413_), .B(new_n315_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n651_));
  AND3_X1   g450(.A1(new_n416_), .A2(new_n410_), .A3(new_n417_), .ZN(new_n652_));
  AOI21_X1  g451(.A(new_n427_), .B1(new_n311_), .B2(new_n314_), .ZN(new_n653_));
  OAI21_X1  g452(.A(new_n384_), .B1(new_n652_), .B2(new_n653_), .ZN(new_n654_));
  AOI21_X1  g453(.A(new_n265_), .B1(new_n651_), .B2(new_n654_), .ZN(new_n655_));
  OAI211_X1 g454(.A(new_n384_), .B(new_n315_), .C1(new_n649_), .C2(new_n650_), .ZN(new_n656_));
  NAND3_X1  g455(.A1(new_n262_), .A2(new_n263_), .A3(new_n411_), .ZN(new_n657_));
  NOR2_X1   g456(.A1(new_n656_), .A2(new_n657_), .ZN(new_n658_));
  OAI211_X1 g457(.A(new_n646_), .B(new_n648_), .C1(new_n655_), .C2(new_n658_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n659_), .A2(KEYINPUT43), .ZN(new_n660_));
  NOR2_X1   g459(.A1(new_n595_), .A2(KEYINPUT43), .ZN(new_n661_));
  NAND2_X1  g460(.A1(new_n430_), .A2(new_n661_), .ZN(new_n662_));
  NAND2_X1  g461(.A1(new_n660_), .A2(new_n662_), .ZN(new_n663_));
  NOR2_X1   g462(.A1(new_n606_), .A2(new_n567_), .ZN(new_n664_));
  NAND3_X1  g463(.A1(new_n663_), .A2(KEYINPUT44), .A3(new_n664_), .ZN(new_n665_));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666_));
  AOI22_X1  g465(.A1(new_n659_), .A2(KEYINPUT43), .B1(new_n430_), .B2(new_n661_), .ZN(new_n667_));
  INV_X1    g466(.A(new_n664_), .ZN(new_n668_));
  OAI21_X1  g467(.A(new_n666_), .B1(new_n667_), .B2(new_n668_), .ZN(new_n669_));
  NAND3_X1  g468(.A1(new_n665_), .A2(new_n669_), .A3(new_n410_), .ZN(new_n670_));
  INV_X1    g469(.A(KEYINPUT109), .ZN(new_n671_));
  AND2_X1   g470(.A1(new_n670_), .A2(new_n671_), .ZN(new_n672_));
  OAI21_X1  g471(.A(G29gat), .B1(new_n670_), .B2(new_n671_), .ZN(new_n673_));
  OAI21_X1  g472(.A(new_n644_), .B1(new_n672_), .B2(new_n673_), .ZN(new_n674_));
  NAND2_X1  g473(.A1(new_n674_), .A2(KEYINPUT110), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT110), .ZN(new_n676_));
  OAI211_X1 g475(.A(new_n676_), .B(new_n644_), .C1(new_n672_), .C2(new_n673_), .ZN(new_n677_));
  NAND2_X1  g476(.A1(new_n675_), .A2(new_n677_), .ZN(G1328gat));
  OR2_X1    g477(.A1(new_n342_), .A2(G36gat), .ZN(new_n679_));
  OR3_X1    g478(.A1(new_n643_), .A2(KEYINPUT45), .A3(new_n679_), .ZN(new_n680_));
  OAI21_X1  g479(.A(KEYINPUT45), .B1(new_n643_), .B2(new_n679_), .ZN(new_n681_));
  INV_X1    g480(.A(KEYINPUT46), .ZN(new_n682_));
  AOI22_X1  g481(.A1(new_n680_), .A2(new_n681_), .B1(KEYINPUT111), .B2(new_n682_), .ZN(new_n683_));
  NAND3_X1  g482(.A1(new_n665_), .A2(new_n669_), .A3(new_n614_), .ZN(new_n684_));
  NAND2_X1  g483(.A1(new_n684_), .A2(G36gat), .ZN(new_n685_));
  AND2_X1   g484(.A1(new_n683_), .A2(new_n685_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n682_), .A2(KEYINPUT111), .ZN(new_n687_));
  XNOR2_X1  g486(.A(new_n686_), .B(new_n687_), .ZN(G1329gat));
  NAND2_X1  g487(.A1(new_n665_), .A2(new_n669_), .ZN(new_n689_));
  OAI21_X1  g488(.A(G43gat), .B1(new_n689_), .B2(new_n264_), .ZN(new_n690_));
  OR2_X1    g489(.A1(new_n264_), .A2(G43gat), .ZN(new_n691_));
  OAI21_X1  g490(.A(new_n690_), .B1(new_n643_), .B2(new_n691_), .ZN(new_n692_));
  INV_X1    g491(.A(KEYINPUT47), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n692_), .B(new_n693_), .ZN(G1330gat));
  INV_X1    g493(.A(G50gat), .ZN(new_n695_));
  NOR3_X1   g494(.A1(new_n689_), .A2(new_n695_), .A3(new_n384_), .ZN(new_n696_));
  NAND3_X1  g495(.A1(new_n464_), .A2(new_n633_), .A3(new_n642_), .ZN(new_n697_));
  AOI21_X1  g496(.A(new_n696_), .B1(new_n695_), .B2(new_n697_), .ZN(G1331gat));
  NOR3_X1   g497(.A1(new_n551_), .A2(new_n463_), .A3(new_n566_), .ZN(new_n699_));
  NAND2_X1  g498(.A1(new_n600_), .A2(new_n699_), .ZN(new_n700_));
  OAI21_X1  g499(.A(G57gat), .B1(new_n700_), .B2(new_n411_), .ZN(new_n701_));
  NAND2_X1  g500(.A1(new_n430_), .A2(new_n602_), .ZN(new_n702_));
  NAND2_X1  g501(.A1(new_n595_), .A2(new_n567_), .ZN(new_n703_));
  NOR3_X1   g502(.A1(new_n702_), .A2(new_n551_), .A3(new_n703_), .ZN(new_n704_));
  INV_X1    g503(.A(new_n704_), .ZN(new_n705_));
  OR2_X1    g504(.A1(new_n411_), .A2(G57gat), .ZN(new_n706_));
  OAI21_X1  g505(.A(new_n701_), .B1(new_n705_), .B2(new_n706_), .ZN(G1332gat));
  OAI21_X1  g506(.A(G64gat), .B1(new_n700_), .B2(new_n342_), .ZN(new_n708_));
  XNOR2_X1  g507(.A(new_n708_), .B(KEYINPUT48), .ZN(new_n709_));
  OR2_X1    g508(.A1(new_n342_), .A2(G64gat), .ZN(new_n710_));
  OAI21_X1  g509(.A(new_n709_), .B1(new_n705_), .B2(new_n710_), .ZN(G1333gat));
  OAI21_X1  g510(.A(G71gat), .B1(new_n700_), .B2(new_n264_), .ZN(new_n712_));
  XNOR2_X1  g511(.A(new_n712_), .B(KEYINPUT49), .ZN(new_n713_));
  NOR2_X1   g512(.A1(new_n264_), .A2(G71gat), .ZN(new_n714_));
  XNOR2_X1  g513(.A(new_n714_), .B(KEYINPUT112), .ZN(new_n715_));
  NAND2_X1  g514(.A1(new_n704_), .A2(new_n715_), .ZN(new_n716_));
  NAND2_X1  g515(.A1(new_n713_), .A2(new_n716_), .ZN(new_n717_));
  INV_X1    g516(.A(KEYINPUT113), .ZN(new_n718_));
  XNOR2_X1  g517(.A(new_n717_), .B(new_n718_), .ZN(G1334gat));
  OAI21_X1  g518(.A(G78gat), .B1(new_n700_), .B2(new_n384_), .ZN(new_n720_));
  XNOR2_X1  g519(.A(new_n720_), .B(KEYINPUT50), .ZN(new_n721_));
  OR2_X1    g520(.A1(new_n384_), .A2(G78gat), .ZN(new_n722_));
  OAI21_X1  g521(.A(new_n721_), .B1(new_n705_), .B2(new_n722_), .ZN(G1335gat));
  NOR3_X1   g522(.A1(new_n702_), .A2(new_n551_), .A3(new_n641_), .ZN(new_n724_));
  AOI21_X1  g523(.A(G85gat), .B1(new_n724_), .B2(new_n410_), .ZN(new_n725_));
  NOR3_X1   g524(.A1(new_n551_), .A2(new_n463_), .A3(new_n567_), .ZN(new_n726_));
  INV_X1    g525(.A(new_n726_), .ZN(new_n727_));
  AOI21_X1  g526(.A(new_n727_), .B1(new_n660_), .B2(new_n662_), .ZN(new_n728_));
  AND2_X1   g527(.A1(new_n410_), .A2(new_n472_), .ZN(new_n729_));
  AOI21_X1  g528(.A(new_n725_), .B1(new_n728_), .B2(new_n729_), .ZN(G1336gat));
  INV_X1    g529(.A(new_n728_), .ZN(new_n731_));
  OAI21_X1  g530(.A(G92gat), .B1(new_n731_), .B2(new_n342_), .ZN(new_n732_));
  INV_X1    g531(.A(G92gat), .ZN(new_n733_));
  NAND3_X1  g532(.A1(new_n724_), .A2(new_n733_), .A3(new_n614_), .ZN(new_n734_));
  NAND2_X1  g533(.A1(new_n732_), .A2(new_n734_), .ZN(G1337gat));
  OAI21_X1  g534(.A(G99gat), .B1(new_n731_), .B2(new_n264_), .ZN(new_n736_));
  NAND3_X1  g535(.A1(new_n724_), .A2(new_n265_), .A3(new_n469_), .ZN(new_n737_));
  NAND2_X1  g536(.A1(new_n736_), .A2(new_n737_), .ZN(new_n738_));
  XNOR2_X1  g537(.A(new_n738_), .B(KEYINPUT51), .ZN(G1338gat));
  NAND3_X1  g538(.A1(new_n724_), .A2(new_n470_), .A3(new_n633_), .ZN(new_n740_));
  INV_X1    g539(.A(KEYINPUT52), .ZN(new_n741_));
  NOR3_X1   g540(.A1(new_n667_), .A2(new_n384_), .A3(new_n727_), .ZN(new_n742_));
  AOI21_X1  g541(.A(new_n470_), .B1(new_n742_), .B2(KEYINPUT114), .ZN(new_n743_));
  AOI21_X1  g542(.A(KEYINPUT114), .B1(new_n728_), .B2(new_n633_), .ZN(new_n744_));
  INV_X1    g543(.A(new_n744_), .ZN(new_n745_));
  AOI21_X1  g544(.A(new_n741_), .B1(new_n743_), .B2(new_n745_), .ZN(new_n746_));
  NAND4_X1  g545(.A1(new_n663_), .A2(KEYINPUT114), .A3(new_n633_), .A4(new_n726_), .ZN(new_n747_));
  NAND2_X1  g546(.A1(new_n747_), .A2(G106gat), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n748_), .A2(KEYINPUT52), .A3(new_n744_), .ZN(new_n749_));
  OAI21_X1  g548(.A(new_n740_), .B1(new_n746_), .B2(new_n749_), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n750_), .A2(KEYINPUT53), .ZN(new_n751_));
  INV_X1    g550(.A(KEYINPUT53), .ZN(new_n752_));
  OAI211_X1 g551(.A(new_n752_), .B(new_n740_), .C1(new_n746_), .C2(new_n749_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n751_), .A2(new_n753_), .ZN(G1339gat));
  NAND4_X1  g553(.A1(new_n551_), .A2(new_n595_), .A3(new_n602_), .A4(new_n567_), .ZN(new_n755_));
  INV_X1    g554(.A(KEYINPUT54), .ZN(new_n756_));
  XNOR2_X1  g555(.A(new_n755_), .B(new_n756_), .ZN(new_n757_));
  INV_X1    g556(.A(KEYINPUT56), .ZN(new_n758_));
  OAI21_X1  g557(.A(new_n526_), .B1(new_n506_), .B2(new_n529_), .ZN(new_n759_));
  INV_X1    g558(.A(new_n467_), .ZN(new_n760_));
  INV_X1    g559(.A(new_n514_), .ZN(new_n761_));
  AOI21_X1  g560(.A(new_n760_), .B1(new_n527_), .B2(new_n761_), .ZN(new_n762_));
  OAI21_X1  g561(.A(new_n533_), .B1(new_n759_), .B2(new_n762_), .ZN(new_n763_));
  NAND2_X1  g562(.A1(new_n763_), .A2(KEYINPUT115), .ZN(new_n764_));
  INV_X1    g563(.A(KEYINPUT115), .ZN(new_n765_));
  OAI211_X1 g564(.A(new_n765_), .B(new_n533_), .C1(new_n759_), .C2(new_n762_), .ZN(new_n766_));
  NAND2_X1  g565(.A1(new_n532_), .A2(KEYINPUT55), .ZN(new_n767_));
  AOI21_X1  g566(.A(new_n529_), .B1(new_n524_), .B2(new_n525_), .ZN(new_n768_));
  NOR2_X1   g567(.A1(new_n534_), .A2(new_n768_), .ZN(new_n769_));
  INV_X1    g568(.A(KEYINPUT55), .ZN(new_n770_));
  NAND4_X1  g569(.A1(new_n769_), .A2(new_n770_), .A3(new_n516_), .A4(new_n515_), .ZN(new_n771_));
  AOI22_X1  g570(.A1(new_n764_), .A2(new_n766_), .B1(new_n767_), .B2(new_n771_), .ZN(new_n772_));
  INV_X1    g571(.A(new_n542_), .ZN(new_n773_));
  OAI21_X1  g572(.A(new_n758_), .B1(new_n772_), .B2(new_n773_), .ZN(new_n774_));
  NOR2_X1   g573(.A1(new_n773_), .A2(new_n758_), .ZN(new_n775_));
  INV_X1    g574(.A(new_n775_), .ZN(new_n776_));
  OAI21_X1  g575(.A(KEYINPUT116), .B1(new_n772_), .B2(new_n776_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n764_), .A2(new_n766_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n767_), .A2(new_n771_), .ZN(new_n779_));
  NAND2_X1  g578(.A1(new_n778_), .A2(new_n779_), .ZN(new_n780_));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n781_));
  NAND3_X1  g580(.A1(new_n780_), .A2(new_n781_), .A3(new_n775_), .ZN(new_n782_));
  NAND3_X1  g581(.A1(new_n774_), .A2(new_n777_), .A3(new_n782_), .ZN(new_n783_));
  NOR2_X1   g582(.A1(new_n602_), .A2(new_n545_), .ZN(new_n784_));
  NAND2_X1  g583(.A1(new_n783_), .A2(new_n784_), .ZN(new_n785_));
  NAND2_X1  g584(.A1(new_n446_), .A2(new_n449_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n447_), .B1(new_n786_), .B2(KEYINPUT117), .ZN(new_n787_));
  OAI21_X1  g586(.A(new_n787_), .B1(KEYINPUT117), .B2(new_n786_), .ZN(new_n788_));
  AOI21_X1  g587(.A(new_n456_), .B1(new_n451_), .B2(new_n447_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND2_X1  g589(.A1(new_n461_), .A2(new_n790_), .ZN(new_n791_));
  AOI21_X1  g590(.A(new_n791_), .B1(new_n547_), .B2(new_n543_), .ZN(new_n792_));
  INV_X1    g591(.A(new_n792_), .ZN(new_n793_));
  NAND2_X1  g592(.A1(new_n785_), .A2(new_n793_), .ZN(new_n794_));
  NAND3_X1  g593(.A1(new_n794_), .A2(KEYINPUT57), .A3(new_n593_), .ZN(new_n795_));
  NOR2_X1   g594(.A1(new_n791_), .A2(new_n545_), .ZN(new_n796_));
  AOI21_X1  g595(.A(KEYINPUT56), .B1(new_n780_), .B2(new_n542_), .ZN(new_n797_));
  NOR2_X1   g596(.A1(new_n772_), .A2(new_n776_), .ZN(new_n798_));
  OAI21_X1  g597(.A(new_n796_), .B1(new_n797_), .B2(new_n798_), .ZN(new_n799_));
  NOR2_X1   g598(.A1(KEYINPUT118), .A2(KEYINPUT58), .ZN(new_n800_));
  NAND2_X1  g599(.A1(new_n799_), .A2(new_n800_), .ZN(new_n801_));
  OAI221_X1 g600(.A(new_n796_), .B1(KEYINPUT118), .B2(KEYINPUT58), .C1(new_n797_), .C2(new_n798_), .ZN(new_n802_));
  NAND3_X1  g601(.A1(new_n801_), .A2(new_n802_), .A3(new_n645_), .ZN(new_n803_));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n804_));
  AOI21_X1  g603(.A(new_n792_), .B1(new_n783_), .B2(new_n784_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n804_), .B1(new_n805_), .B2(new_n640_), .ZN(new_n806_));
  NAND3_X1  g605(.A1(new_n795_), .A2(new_n803_), .A3(new_n806_), .ZN(new_n807_));
  AOI21_X1  g606(.A(new_n757_), .B1(new_n807_), .B2(new_n566_), .ZN(new_n808_));
  NOR3_X1   g607(.A1(new_n656_), .A2(new_n411_), .A3(new_n264_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n809_), .ZN(new_n810_));
  NOR2_X1   g609(.A1(new_n808_), .A2(new_n810_), .ZN(new_n811_));
  INV_X1    g610(.A(G113gat), .ZN(new_n812_));
  NAND3_X1  g611(.A1(new_n811_), .A2(new_n812_), .A3(new_n463_), .ZN(new_n813_));
  NAND2_X1  g612(.A1(new_n806_), .A2(new_n803_), .ZN(new_n814_));
  NOR3_X1   g613(.A1(new_n805_), .A2(new_n804_), .A3(new_n640_), .ZN(new_n815_));
  OAI21_X1  g614(.A(new_n566_), .B1(new_n814_), .B2(new_n815_), .ZN(new_n816_));
  INV_X1    g615(.A(new_n757_), .ZN(new_n817_));
  NAND2_X1  g616(.A1(new_n816_), .A2(new_n817_), .ZN(new_n818_));
  XOR2_X1   g617(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n819_));
  NAND3_X1  g618(.A1(new_n818_), .A2(new_n809_), .A3(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(KEYINPUT120), .ZN(new_n821_));
  OAI21_X1  g620(.A(KEYINPUT59), .B1(new_n808_), .B2(new_n810_), .ZN(new_n822_));
  AND3_X1   g621(.A1(new_n820_), .A2(new_n821_), .A3(new_n822_), .ZN(new_n823_));
  AOI21_X1  g622(.A(new_n821_), .B1(new_n820_), .B2(new_n822_), .ZN(new_n824_));
  NOR3_X1   g623(.A1(new_n823_), .A2(new_n824_), .A3(new_n602_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n813_), .B1(new_n825_), .B2(new_n812_), .ZN(G1340gat));
  NAND2_X1  g625(.A1(new_n820_), .A2(new_n822_), .ZN(new_n827_));
  OAI21_X1  g626(.A(G120gat), .B1(new_n827_), .B2(new_n551_), .ZN(new_n828_));
  NAND2_X1  g627(.A1(new_n818_), .A2(new_n809_), .ZN(new_n829_));
  INV_X1    g628(.A(G120gat), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n830_), .B1(new_n551_), .B2(KEYINPUT60), .ZN(new_n831_));
  OAI21_X1  g630(.A(new_n831_), .B1(KEYINPUT60), .B2(new_n830_), .ZN(new_n832_));
  OAI21_X1  g631(.A(new_n828_), .B1(new_n829_), .B2(new_n832_), .ZN(G1341gat));
  INV_X1    g632(.A(G127gat), .ZN(new_n834_));
  NAND3_X1  g633(.A1(new_n811_), .A2(new_n834_), .A3(new_n567_), .ZN(new_n835_));
  NOR3_X1   g634(.A1(new_n823_), .A2(new_n824_), .A3(new_n566_), .ZN(new_n836_));
  OAI21_X1  g635(.A(new_n835_), .B1(new_n836_), .B2(new_n834_), .ZN(G1342gat));
  INV_X1    g636(.A(G134gat), .ZN(new_n838_));
  NOR2_X1   g637(.A1(new_n595_), .A2(new_n838_), .ZN(new_n839_));
  INV_X1    g638(.A(new_n839_), .ZN(new_n840_));
  NOR3_X1   g639(.A1(new_n823_), .A2(new_n824_), .A3(new_n840_), .ZN(new_n841_));
  OAI21_X1  g640(.A(new_n838_), .B1(new_n829_), .B2(new_n593_), .ZN(new_n842_));
  INV_X1    g641(.A(KEYINPUT121), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n842_), .A2(new_n843_), .ZN(new_n844_));
  OAI211_X1 g643(.A(KEYINPUT121), .B(new_n838_), .C1(new_n829_), .C2(new_n593_), .ZN(new_n845_));
  NAND2_X1  g644(.A1(new_n844_), .A2(new_n845_), .ZN(new_n846_));
  OAI21_X1  g645(.A(KEYINPUT122), .B1(new_n841_), .B2(new_n846_), .ZN(new_n847_));
  NAND2_X1  g646(.A1(new_n827_), .A2(KEYINPUT120), .ZN(new_n848_));
  NAND3_X1  g647(.A1(new_n820_), .A2(new_n822_), .A3(new_n821_), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n848_), .A2(new_n849_), .A3(new_n839_), .ZN(new_n850_));
  INV_X1    g649(.A(KEYINPUT122), .ZN(new_n851_));
  NAND4_X1  g650(.A1(new_n850_), .A2(new_n851_), .A3(new_n844_), .A4(new_n845_), .ZN(new_n852_));
  NAND2_X1  g651(.A1(new_n847_), .A2(new_n852_), .ZN(G1343gat));
  NAND4_X1  g652(.A1(new_n342_), .A2(new_n633_), .A3(new_n410_), .A4(new_n264_), .ZN(new_n854_));
  NOR2_X1   g653(.A1(new_n808_), .A2(new_n854_), .ZN(new_n855_));
  XNOR2_X1  g654(.A(new_n855_), .B(KEYINPUT123), .ZN(new_n856_));
  NOR2_X1   g655(.A1(new_n856_), .A2(new_n602_), .ZN(new_n857_));
  XNOR2_X1  g656(.A(new_n857_), .B(new_n355_), .ZN(G1344gat));
  NOR2_X1   g657(.A1(new_n856_), .A2(new_n551_), .ZN(new_n859_));
  XNOR2_X1  g658(.A(new_n859_), .B(new_n356_), .ZN(G1345gat));
  NOR2_X1   g659(.A1(new_n856_), .A2(new_n566_), .ZN(new_n861_));
  XOR2_X1   g660(.A(KEYINPUT61), .B(G155gat), .Z(new_n862_));
  XNOR2_X1  g661(.A(new_n861_), .B(new_n862_), .ZN(G1346gat));
  NAND3_X1  g662(.A1(new_n646_), .A2(G162gat), .A3(new_n648_), .ZN(new_n864_));
  NOR2_X1   g663(.A1(new_n856_), .A2(new_n864_), .ZN(new_n865_));
  INV_X1    g664(.A(new_n854_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n818_), .A2(new_n866_), .ZN(new_n867_));
  NAND2_X1  g666(.A1(new_n867_), .A2(KEYINPUT123), .ZN(new_n868_));
  INV_X1    g667(.A(KEYINPUT123), .ZN(new_n869_));
  NAND2_X1  g668(.A1(new_n855_), .A2(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n593_), .B1(new_n868_), .B2(new_n870_), .ZN(new_n871_));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n872_));
  OR3_X1    g671(.A1(new_n871_), .A2(new_n872_), .A3(G162gat), .ZN(new_n873_));
  OAI21_X1  g672(.A(new_n872_), .B1(new_n871_), .B2(G162gat), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n865_), .B1(new_n873_), .B2(new_n874_), .ZN(G1347gat));
  NOR2_X1   g674(.A1(new_n808_), .A2(new_n342_), .ZN(new_n876_));
  NOR2_X1   g675(.A1(new_n657_), .A2(new_n633_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n876_), .A2(new_n877_), .ZN(new_n878_));
  INV_X1    g677(.A(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n879_), .A2(new_n463_), .ZN(new_n880_));
  INV_X1    g679(.A(KEYINPUT62), .ZN(new_n881_));
  AND3_X1   g680(.A1(new_n880_), .A2(new_n881_), .A3(G169gat), .ZN(new_n882_));
  AOI21_X1  g681(.A(new_n881_), .B1(new_n880_), .B2(G169gat), .ZN(new_n883_));
  OR2_X1    g682(.A1(new_n878_), .A2(KEYINPUT125), .ZN(new_n884_));
  NAND2_X1  g683(.A1(new_n878_), .A2(KEYINPUT125), .ZN(new_n885_));
  NAND2_X1  g684(.A1(new_n884_), .A2(new_n885_), .ZN(new_n886_));
  INV_X1    g685(.A(new_n886_), .ZN(new_n887_));
  NOR2_X1   g686(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n888_));
  AND2_X1   g687(.A1(KEYINPUT22), .A2(G169gat), .ZN(new_n889_));
  OAI21_X1  g688(.A(new_n463_), .B1(new_n888_), .B2(new_n889_), .ZN(new_n890_));
  OAI22_X1  g689(.A1(new_n882_), .A2(new_n883_), .B1(new_n887_), .B2(new_n890_), .ZN(G1348gat));
  OAI21_X1  g690(.A(G176gat), .B1(new_n878_), .B2(new_n551_), .ZN(new_n892_));
  OR2_X1    g691(.A1(new_n551_), .A2(G176gat), .ZN(new_n893_));
  OAI21_X1  g692(.A(new_n892_), .B1(new_n887_), .B2(new_n893_), .ZN(G1349gat));
  NAND2_X1  g693(.A1(new_n567_), .A2(new_n288_), .ZN(new_n895_));
  INV_X1    g694(.A(new_n895_), .ZN(new_n896_));
  NAND2_X1  g695(.A1(new_n879_), .A2(new_n567_), .ZN(new_n897_));
  AOI22_X1  g696(.A1(new_n886_), .A2(new_n896_), .B1(new_n207_), .B2(new_n897_), .ZN(G1350gat));
  OR2_X1    g697(.A1(new_n593_), .A2(new_n221_), .ZN(new_n899_));
  AOI21_X1  g698(.A(new_n595_), .B1(new_n884_), .B2(new_n885_), .ZN(new_n900_));
  OAI22_X1  g699(.A1(new_n887_), .A2(new_n899_), .B1(new_n900_), .B2(new_n208_), .ZN(G1351gat));
  AND2_X1   g700(.A1(new_n264_), .A2(new_n413_), .ZN(new_n902_));
  AND2_X1   g701(.A1(new_n876_), .A2(new_n902_), .ZN(new_n903_));
  NAND2_X1  g702(.A1(new_n903_), .A2(new_n463_), .ZN(new_n904_));
  XNOR2_X1  g703(.A(new_n904_), .B(G197gat), .ZN(G1352gat));
  NAND2_X1  g704(.A1(new_n903_), .A2(new_n601_), .ZN(new_n906_));
  XNOR2_X1  g705(.A(new_n906_), .B(G204gat), .ZN(G1353gat));
  XNOR2_X1  g706(.A(KEYINPUT63), .B(G211gat), .ZN(new_n908_));
  NAND3_X1  g707(.A1(new_n903_), .A2(new_n567_), .A3(new_n908_), .ZN(new_n909_));
  NAND2_X1  g708(.A1(new_n876_), .A2(new_n902_), .ZN(new_n910_));
  OAI22_X1  g709(.A1(new_n910_), .A2(new_n566_), .B1(KEYINPUT63), .B2(G211gat), .ZN(new_n911_));
  NAND2_X1  g710(.A1(new_n909_), .A2(new_n911_), .ZN(new_n912_));
  INV_X1    g711(.A(KEYINPUT126), .ZN(new_n913_));
  XNOR2_X1  g712(.A(new_n912_), .B(new_n913_), .ZN(G1354gat));
  OR3_X1    g713(.A1(new_n910_), .A2(G218gat), .A3(new_n593_), .ZN(new_n915_));
  OAI21_X1  g714(.A(G218gat), .B1(new_n910_), .B2(new_n595_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n915_), .A2(new_n916_), .ZN(G1355gat));
endmodule


