//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 0 1 1 0 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:27:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n749_,
    new_n750_, new_n751_, new_n752_, new_n753_, new_n754_, new_n755_,
    new_n756_, new_n757_, new_n758_, new_n759_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n794_, new_n795_, new_n796_, new_n797_,
    new_n798_, new_n799_, new_n801_, new_n802_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n835_,
    new_n836_, new_n837_, new_n838_, new_n839_, new_n840_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n850_, new_n851_, new_n852_, new_n853_,
    new_n854_, new_n855_, new_n856_, new_n857_, new_n858_, new_n859_,
    new_n860_, new_n861_, new_n862_, new_n863_, new_n864_, new_n865_,
    new_n866_, new_n867_, new_n868_, new_n869_, new_n870_, new_n871_,
    new_n872_, new_n873_, new_n874_, new_n875_, new_n876_, new_n877_,
    new_n878_, new_n879_, new_n880_, new_n881_, new_n882_, new_n883_,
    new_n884_, new_n885_, new_n886_, new_n887_, new_n888_, new_n889_,
    new_n890_, new_n891_, new_n892_, new_n893_, new_n894_, new_n895_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n916_, new_n917_, new_n918_, new_n920_, new_n921_, new_n922_,
    new_n924_, new_n925_, new_n926_, new_n928_, new_n930_, new_n931_,
    new_n933_, new_n934_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n958_, new_n959_,
    new_n960_, new_n961_, new_n963_, new_n964_, new_n966_, new_n967_,
    new_n968_, new_n970_, new_n971_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n978_, new_n979_;
  NAND2_X1  g000(.A1(G226gat), .A2(G233gat), .ZN(new_n202_));
  XNOR2_X1  g001(.A(new_n202_), .B(KEYINPUT19), .ZN(new_n203_));
  INV_X1    g002(.A(new_n203_), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n204_), .A2(KEYINPUT20), .ZN(new_n205_));
  INV_X1    g004(.A(new_n205_), .ZN(new_n206_));
  XOR2_X1   g005(.A(G211gat), .B(G218gat), .Z(new_n207_));
  INV_X1    g006(.A(new_n207_), .ZN(new_n208_));
  INV_X1    g007(.A(G197gat), .ZN(new_n209_));
  INV_X1    g008(.A(G204gat), .ZN(new_n210_));
  NAND2_X1  g009(.A1(new_n209_), .A2(new_n210_), .ZN(new_n211_));
  NAND2_X1  g010(.A1(G197gat), .A2(G204gat), .ZN(new_n212_));
  NAND3_X1  g011(.A1(new_n211_), .A2(KEYINPUT21), .A3(new_n212_), .ZN(new_n213_));
  NOR2_X1   g012(.A1(new_n208_), .A2(new_n213_), .ZN(new_n214_));
  INV_X1    g013(.A(new_n214_), .ZN(new_n215_));
  INV_X1    g014(.A(KEYINPUT86), .ZN(new_n216_));
  NAND2_X1  g015(.A1(new_n213_), .A2(new_n216_), .ZN(new_n217_));
  NAND4_X1  g016(.A1(new_n211_), .A2(KEYINPUT86), .A3(KEYINPUT21), .A4(new_n212_), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n217_), .A2(new_n218_), .ZN(new_n219_));
  AOI21_X1  g018(.A(KEYINPUT21), .B1(new_n211_), .B2(new_n212_), .ZN(new_n220_));
  NOR2_X1   g019(.A1(new_n220_), .A2(new_n207_), .ZN(new_n221_));
  AND3_X1   g020(.A1(new_n219_), .A2(KEYINPUT87), .A3(new_n221_), .ZN(new_n222_));
  AOI21_X1  g021(.A(KEYINPUT87), .B1(new_n219_), .B2(new_n221_), .ZN(new_n223_));
  OAI21_X1  g022(.A(new_n215_), .B1(new_n222_), .B2(new_n223_), .ZN(new_n224_));
  INV_X1    g023(.A(G169gat), .ZN(new_n225_));
  INV_X1    g024(.A(G176gat), .ZN(new_n226_));
  NOR2_X1   g025(.A1(new_n225_), .A2(new_n226_), .ZN(new_n227_));
  OAI21_X1  g026(.A(KEYINPUT24), .B1(G169gat), .B2(G176gat), .ZN(new_n228_));
  OR2_X1    g027(.A1(new_n227_), .A2(new_n228_), .ZN(new_n229_));
  NOR3_X1   g028(.A1(KEYINPUT24), .A2(G169gat), .A3(G176gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(G183gat), .A2(G190gat), .ZN(new_n231_));
  NAND2_X1  g030(.A1(new_n231_), .A2(KEYINPUT23), .ZN(new_n232_));
  INV_X1    g031(.A(KEYINPUT23), .ZN(new_n233_));
  NAND3_X1  g032(.A1(new_n233_), .A2(G183gat), .A3(G190gat), .ZN(new_n234_));
  AOI21_X1  g033(.A(new_n230_), .B1(new_n232_), .B2(new_n234_), .ZN(new_n235_));
  XNOR2_X1  g034(.A(KEYINPUT25), .B(G183gat), .ZN(new_n236_));
  XNOR2_X1  g035(.A(KEYINPUT26), .B(G190gat), .ZN(new_n237_));
  NAND2_X1  g036(.A1(new_n236_), .A2(new_n237_), .ZN(new_n238_));
  NAND3_X1  g037(.A1(new_n229_), .A2(new_n235_), .A3(new_n238_), .ZN(new_n239_));
  NOR2_X1   g038(.A1(KEYINPUT22), .A2(G176gat), .ZN(new_n240_));
  XNOR2_X1  g039(.A(new_n240_), .B(G169gat), .ZN(new_n241_));
  AND2_X1   g040(.A1(new_n232_), .A2(new_n234_), .ZN(new_n242_));
  NOR2_X1   g041(.A1(G183gat), .A2(G190gat), .ZN(new_n243_));
  OAI21_X1  g042(.A(new_n241_), .B1(new_n242_), .B2(new_n243_), .ZN(new_n244_));
  NAND2_X1  g043(.A1(new_n239_), .A2(new_n244_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n206_), .B1(new_n224_), .B2(new_n245_), .ZN(new_n246_));
  INV_X1    g045(.A(KEYINPUT90), .ZN(new_n247_));
  NAND2_X1  g046(.A1(new_n219_), .A2(new_n221_), .ZN(new_n248_));
  INV_X1    g047(.A(KEYINPUT87), .ZN(new_n249_));
  NAND2_X1  g048(.A1(new_n248_), .A2(new_n249_), .ZN(new_n250_));
  NAND3_X1  g049(.A1(new_n219_), .A2(KEYINPUT87), .A3(new_n221_), .ZN(new_n251_));
  AOI21_X1  g050(.A(new_n214_), .B1(new_n250_), .B2(new_n251_), .ZN(new_n252_));
  AOI21_X1  g051(.A(new_n243_), .B1(new_n233_), .B2(new_n231_), .ZN(new_n253_));
  OAI21_X1  g052(.A(new_n253_), .B1(new_n233_), .B2(new_n231_), .ZN(new_n254_));
  NAND2_X1  g053(.A1(new_n254_), .A2(new_n241_), .ZN(new_n255_));
  NAND2_X1  g054(.A1(new_n229_), .A2(KEYINPUT79), .ZN(new_n256_));
  NAND2_X1  g055(.A1(new_n256_), .A2(new_n235_), .ZN(new_n257_));
  INV_X1    g056(.A(G183gat), .ZN(new_n258_));
  OAI21_X1  g057(.A(KEYINPUT78), .B1(new_n258_), .B2(KEYINPUT25), .ZN(new_n259_));
  OAI211_X1 g058(.A(new_n259_), .B(new_n237_), .C1(new_n236_), .C2(KEYINPUT78), .ZN(new_n260_));
  OR3_X1    g059(.A1(new_n227_), .A2(new_n228_), .A3(KEYINPUT79), .ZN(new_n261_));
  NAND2_X1  g060(.A1(new_n260_), .A2(new_n261_), .ZN(new_n262_));
  OAI21_X1  g061(.A(new_n255_), .B1(new_n257_), .B2(new_n262_), .ZN(new_n263_));
  INV_X1    g062(.A(new_n263_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n247_), .B1(new_n252_), .B2(new_n264_), .ZN(new_n265_));
  NAND3_X1  g064(.A1(new_n224_), .A2(KEYINPUT90), .A3(new_n263_), .ZN(new_n266_));
  AOI21_X1  g065(.A(new_n246_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n252_), .A2(new_n264_), .ZN(new_n268_));
  NAND2_X1  g067(.A1(new_n224_), .A2(new_n245_), .ZN(new_n269_));
  NAND3_X1  g068(.A1(new_n268_), .A2(new_n269_), .A3(KEYINPUT20), .ZN(new_n270_));
  AOI22_X1  g069(.A1(new_n267_), .A2(KEYINPUT91), .B1(new_n203_), .B2(new_n270_), .ZN(new_n271_));
  XOR2_X1   g070(.A(G8gat), .B(G36gat), .Z(new_n272_));
  XNOR2_X1  g071(.A(KEYINPUT92), .B(KEYINPUT18), .ZN(new_n273_));
  XNOR2_X1  g072(.A(new_n272_), .B(new_n273_), .ZN(new_n274_));
  XNOR2_X1  g073(.A(G64gat), .B(G92gat), .ZN(new_n275_));
  XNOR2_X1  g074(.A(new_n274_), .B(new_n275_), .ZN(new_n276_));
  NAND2_X1  g075(.A1(new_n265_), .A2(new_n266_), .ZN(new_n277_));
  INV_X1    g076(.A(new_n245_), .ZN(new_n278_));
  AOI21_X1  g077(.A(new_n205_), .B1(new_n252_), .B2(new_n278_), .ZN(new_n279_));
  NAND2_X1  g078(.A1(new_n277_), .A2(new_n279_), .ZN(new_n280_));
  INV_X1    g079(.A(KEYINPUT91), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n280_), .A2(new_n281_), .ZN(new_n282_));
  NAND3_X1  g081(.A1(new_n271_), .A2(new_n276_), .A3(new_n282_), .ZN(new_n283_));
  INV_X1    g082(.A(new_n276_), .ZN(new_n284_));
  NOR3_X1   g083(.A1(new_n252_), .A2(new_n264_), .A3(new_n247_), .ZN(new_n285_));
  AOI21_X1  g084(.A(KEYINPUT90), .B1(new_n224_), .B2(new_n263_), .ZN(new_n286_));
  OAI211_X1 g085(.A(KEYINPUT91), .B(new_n279_), .C1(new_n285_), .C2(new_n286_), .ZN(new_n287_));
  NAND2_X1  g086(.A1(new_n270_), .A2(new_n203_), .ZN(new_n288_));
  NAND2_X1  g087(.A1(new_n287_), .A2(new_n288_), .ZN(new_n289_));
  AOI21_X1  g088(.A(KEYINPUT91), .B1(new_n277_), .B2(new_n279_), .ZN(new_n290_));
  OAI21_X1  g089(.A(new_n284_), .B1(new_n289_), .B2(new_n290_), .ZN(new_n291_));
  NAND2_X1  g090(.A1(new_n283_), .A2(new_n291_), .ZN(new_n292_));
  XOR2_X1   g091(.A(KEYINPUT100), .B(KEYINPUT27), .Z(new_n293_));
  INV_X1    g092(.A(KEYINPUT27), .ZN(new_n294_));
  NAND4_X1  g093(.A1(new_n268_), .A2(new_n269_), .A3(KEYINPUT20), .A4(new_n204_), .ZN(new_n295_));
  XOR2_X1   g094(.A(KEYINPUT97), .B(KEYINPUT20), .Z(new_n296_));
  INV_X1    g095(.A(KEYINPUT98), .ZN(new_n297_));
  XNOR2_X1  g096(.A(new_n245_), .B(new_n297_), .ZN(new_n298_));
  OAI21_X1  g097(.A(new_n296_), .B1(new_n298_), .B2(new_n224_), .ZN(new_n299_));
  AOI21_X1  g098(.A(new_n299_), .B1(new_n265_), .B2(new_n266_), .ZN(new_n300_));
  OAI21_X1  g099(.A(new_n295_), .B1(new_n300_), .B2(new_n204_), .ZN(new_n301_));
  AOI21_X1  g100(.A(new_n294_), .B1(new_n301_), .B2(new_n284_), .ZN(new_n302_));
  AOI22_X1  g101(.A1(new_n292_), .A2(new_n293_), .B1(new_n302_), .B2(new_n283_), .ZN(new_n303_));
  NAND2_X1  g102(.A1(G227gat), .A2(G233gat), .ZN(new_n304_));
  XNOR2_X1  g103(.A(new_n304_), .B(G15gat), .ZN(new_n305_));
  XNOR2_X1  g104(.A(new_n305_), .B(G71gat), .ZN(new_n306_));
  XNOR2_X1  g105(.A(KEYINPUT80), .B(G43gat), .ZN(new_n307_));
  INV_X1    g106(.A(G99gat), .ZN(new_n308_));
  XNOR2_X1  g107(.A(new_n307_), .B(new_n308_), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n306_), .B(new_n309_), .ZN(new_n310_));
  INV_X1    g109(.A(KEYINPUT30), .ZN(new_n311_));
  NAND2_X1  g110(.A1(new_n263_), .A2(new_n311_), .ZN(new_n312_));
  OAI211_X1 g111(.A(KEYINPUT30), .B(new_n255_), .C1(new_n257_), .C2(new_n262_), .ZN(new_n313_));
  NAND2_X1  g112(.A1(new_n312_), .A2(new_n313_), .ZN(new_n314_));
  NAND2_X1  g113(.A1(new_n314_), .A2(KEYINPUT81), .ZN(new_n315_));
  INV_X1    g114(.A(KEYINPUT81), .ZN(new_n316_));
  NAND3_X1  g115(.A1(new_n312_), .A2(new_n316_), .A3(new_n313_), .ZN(new_n317_));
  AOI21_X1  g116(.A(new_n310_), .B1(new_n315_), .B2(new_n317_), .ZN(new_n318_));
  INV_X1    g117(.A(new_n317_), .ZN(new_n319_));
  INV_X1    g118(.A(new_n310_), .ZN(new_n320_));
  NOR2_X1   g119(.A1(new_n319_), .A2(new_n320_), .ZN(new_n321_));
  XNOR2_X1  g120(.A(G127gat), .B(G134gat), .ZN(new_n322_));
  XNOR2_X1  g121(.A(G113gat), .B(G120gat), .ZN(new_n323_));
  AND2_X1   g122(.A1(new_n322_), .A2(new_n323_), .ZN(new_n324_));
  NOR2_X1   g123(.A1(new_n322_), .A2(new_n323_), .ZN(new_n325_));
  NOR2_X1   g124(.A1(new_n324_), .A2(new_n325_), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT31), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  OR3_X1    g127(.A1(new_n318_), .A2(new_n321_), .A3(new_n328_), .ZN(new_n329_));
  OAI21_X1  g128(.A(new_n328_), .B1(new_n318_), .B2(new_n321_), .ZN(new_n330_));
  NAND2_X1  g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  INV_X1    g130(.A(new_n331_), .ZN(new_n332_));
  INV_X1    g131(.A(KEYINPUT99), .ZN(new_n333_));
  NAND2_X1  g132(.A1(G225gat), .A2(G233gat), .ZN(new_n334_));
  INV_X1    g133(.A(new_n334_), .ZN(new_n335_));
  INV_X1    g134(.A(KEYINPUT4), .ZN(new_n336_));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n337_));
  INV_X1    g136(.A(G141gat), .ZN(new_n338_));
  INV_X1    g137(.A(G148gat), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n337_), .A2(new_n338_), .A3(new_n339_), .ZN(new_n340_));
  NAND2_X1  g139(.A1(G141gat), .A2(G148gat), .ZN(new_n341_));
  INV_X1    g140(.A(KEYINPUT2), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n341_), .A2(new_n342_), .ZN(new_n343_));
  NAND3_X1  g142(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n344_));
  OAI21_X1  g143(.A(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n345_));
  NAND4_X1  g144(.A1(new_n340_), .A2(new_n343_), .A3(new_n344_), .A4(new_n345_), .ZN(new_n346_));
  OR2_X1    g145(.A1(G155gat), .A2(G162gat), .ZN(new_n347_));
  NAND2_X1  g146(.A1(G155gat), .A2(G162gat), .ZN(new_n348_));
  AND2_X1   g147(.A1(new_n347_), .A2(new_n348_), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n346_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(new_n348_), .A2(KEYINPUT1), .ZN(new_n351_));
  INV_X1    g150(.A(KEYINPUT1), .ZN(new_n352_));
  NAND3_X1  g151(.A1(new_n352_), .A2(G155gat), .A3(G162gat), .ZN(new_n353_));
  NAND3_X1  g152(.A1(new_n351_), .A2(new_n353_), .A3(new_n347_), .ZN(new_n354_));
  XOR2_X1   g153(.A(G141gat), .B(G148gat), .Z(new_n355_));
  NAND2_X1  g154(.A1(new_n354_), .A2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n350_), .A2(new_n356_), .ZN(new_n357_));
  NAND2_X1  g156(.A1(new_n357_), .A2(new_n326_), .ZN(new_n358_));
  INV_X1    g157(.A(new_n322_), .ZN(new_n359_));
  XOR2_X1   g158(.A(G113gat), .B(G120gat), .Z(new_n360_));
  NAND2_X1  g159(.A1(new_n359_), .A2(new_n360_), .ZN(new_n361_));
  NAND2_X1  g160(.A1(new_n322_), .A2(new_n323_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  AOI22_X1  g162(.A1(new_n346_), .A2(new_n349_), .B1(new_n354_), .B2(new_n355_), .ZN(new_n364_));
  NAND2_X1  g163(.A1(new_n363_), .A2(new_n364_), .ZN(new_n365_));
  INV_X1    g164(.A(KEYINPUT93), .ZN(new_n366_));
  NAND3_X1  g165(.A1(new_n358_), .A2(new_n365_), .A3(new_n366_), .ZN(new_n367_));
  NAND3_X1  g166(.A1(new_n363_), .A2(new_n364_), .A3(KEYINPUT93), .ZN(new_n368_));
  AOI21_X1  g167(.A(new_n336_), .B1(new_n367_), .B2(new_n368_), .ZN(new_n369_));
  NAND3_X1  g168(.A1(new_n357_), .A2(new_n326_), .A3(new_n336_), .ZN(new_n370_));
  INV_X1    g169(.A(new_n370_), .ZN(new_n371_));
  OAI21_X1  g170(.A(new_n335_), .B1(new_n369_), .B2(new_n371_), .ZN(new_n372_));
  XNOR2_X1  g171(.A(G1gat), .B(G29gat), .ZN(new_n373_));
  XNOR2_X1  g172(.A(new_n373_), .B(G85gat), .ZN(new_n374_));
  XNOR2_X1  g173(.A(KEYINPUT0), .B(G57gat), .ZN(new_n375_));
  XOR2_X1   g174(.A(new_n374_), .B(new_n375_), .Z(new_n376_));
  INV_X1    g175(.A(new_n376_), .ZN(new_n377_));
  NAND3_X1  g176(.A1(new_n367_), .A2(new_n368_), .A3(new_n334_), .ZN(new_n378_));
  NAND3_X1  g177(.A1(new_n372_), .A2(new_n377_), .A3(new_n378_), .ZN(new_n379_));
  INV_X1    g178(.A(new_n379_), .ZN(new_n380_));
  AOI21_X1  g179(.A(new_n377_), .B1(new_n372_), .B2(new_n378_), .ZN(new_n381_));
  OAI21_X1  g180(.A(new_n333_), .B1(new_n380_), .B2(new_n381_), .ZN(new_n382_));
  INV_X1    g181(.A(new_n381_), .ZN(new_n383_));
  NAND3_X1  g182(.A1(new_n383_), .A2(KEYINPUT99), .A3(new_n379_), .ZN(new_n384_));
  NAND2_X1  g183(.A1(new_n382_), .A2(new_n384_), .ZN(new_n385_));
  NOR2_X1   g184(.A1(new_n332_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387_));
  AOI21_X1  g186(.A(KEYINPUT82), .B1(new_n364_), .B2(new_n387_), .ZN(new_n388_));
  INV_X1    g187(.A(new_n388_), .ZN(new_n389_));
  NAND3_X1  g188(.A1(new_n364_), .A2(KEYINPUT82), .A3(new_n387_), .ZN(new_n390_));
  XOR2_X1   g189(.A(KEYINPUT83), .B(KEYINPUT28), .Z(new_n391_));
  INV_X1    g190(.A(new_n391_), .ZN(new_n392_));
  AND3_X1   g191(.A1(new_n389_), .A2(new_n390_), .A3(new_n392_), .ZN(new_n393_));
  AOI21_X1  g192(.A(new_n392_), .B1(new_n389_), .B2(new_n390_), .ZN(new_n394_));
  XNOR2_X1  g193(.A(G22gat), .B(G50gat), .ZN(new_n395_));
  INV_X1    g194(.A(new_n395_), .ZN(new_n396_));
  OR3_X1    g195(.A1(new_n393_), .A2(new_n394_), .A3(new_n396_), .ZN(new_n397_));
  OAI21_X1  g196(.A(new_n396_), .B1(new_n393_), .B2(new_n394_), .ZN(new_n398_));
  AND2_X1   g197(.A1(new_n397_), .A2(new_n398_), .ZN(new_n399_));
  XNOR2_X1  g198(.A(G78gat), .B(G106gat), .ZN(new_n400_));
  NAND2_X1  g199(.A1(new_n357_), .A2(KEYINPUT29), .ZN(new_n401_));
  NAND2_X1  g200(.A1(new_n224_), .A2(new_n401_), .ZN(new_n402_));
  INV_X1    g201(.A(G228gat), .ZN(new_n403_));
  INV_X1    g202(.A(G233gat), .ZN(new_n404_));
  OR2_X1    g203(.A1(new_n404_), .A2(KEYINPUT84), .ZN(new_n405_));
  NAND2_X1  g204(.A1(new_n404_), .A2(KEYINPUT84), .ZN(new_n406_));
  AOI21_X1  g205(.A(new_n403_), .B1(new_n405_), .B2(new_n406_), .ZN(new_n407_));
  XNOR2_X1  g206(.A(new_n407_), .B(KEYINPUT85), .ZN(new_n408_));
  INV_X1    g207(.A(new_n408_), .ZN(new_n409_));
  NAND2_X1  g208(.A1(new_n402_), .A2(new_n409_), .ZN(new_n410_));
  NAND3_X1  g209(.A1(new_n224_), .A2(new_n401_), .A3(new_n408_), .ZN(new_n411_));
  AOI21_X1  g210(.A(new_n400_), .B1(new_n410_), .B2(new_n411_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(new_n411_), .ZN(new_n413_));
  INV_X1    g212(.A(new_n400_), .ZN(new_n414_));
  NOR2_X1   g213(.A1(new_n413_), .A2(new_n414_), .ZN(new_n415_));
  OAI21_X1  g214(.A(new_n399_), .B1(new_n412_), .B2(new_n415_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n413_), .A2(KEYINPUT88), .ZN(new_n417_));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n410_), .A2(new_n418_), .A3(new_n411_), .ZN(new_n419_));
  NAND4_X1  g218(.A1(new_n417_), .A2(KEYINPUT89), .A3(new_n400_), .A4(new_n419_), .ZN(new_n420_));
  AOI21_X1  g219(.A(new_n412_), .B1(new_n397_), .B2(new_n398_), .ZN(new_n421_));
  NAND2_X1  g220(.A1(new_n420_), .A2(new_n421_), .ZN(new_n422_));
  AOI21_X1  g221(.A(new_n414_), .B1(new_n413_), .B2(KEYINPUT88), .ZN(new_n423_));
  AOI21_X1  g222(.A(KEYINPUT89), .B1(new_n423_), .B2(new_n419_), .ZN(new_n424_));
  OAI21_X1  g223(.A(new_n416_), .B1(new_n422_), .B2(new_n424_), .ZN(new_n425_));
  INV_X1    g224(.A(new_n425_), .ZN(new_n426_));
  AND3_X1   g225(.A1(new_n303_), .A2(new_n386_), .A3(new_n426_), .ZN(new_n427_));
  NAND2_X1  g226(.A1(new_n276_), .A2(KEYINPUT32), .ZN(new_n428_));
  INV_X1    g227(.A(new_n428_), .ZN(new_n429_));
  NAND2_X1  g228(.A1(new_n301_), .A2(new_n429_), .ZN(new_n430_));
  NAND3_X1  g229(.A1(new_n271_), .A2(new_n282_), .A3(new_n428_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n383_), .A2(new_n379_), .ZN(new_n432_));
  NAND3_X1  g231(.A1(new_n430_), .A2(new_n431_), .A3(new_n432_), .ZN(new_n433_));
  INV_X1    g232(.A(KEYINPUT94), .ZN(new_n434_));
  NAND3_X1  g233(.A1(new_n367_), .A2(new_n434_), .A3(new_n368_), .ZN(new_n435_));
  AND2_X1   g234(.A1(new_n435_), .A2(new_n335_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n367_), .A2(new_n368_), .ZN(new_n437_));
  NAND2_X1  g236(.A1(new_n437_), .A2(KEYINPUT94), .ZN(new_n438_));
  AOI21_X1  g237(.A(new_n376_), .B1(new_n436_), .B2(new_n438_), .ZN(new_n439_));
  NAND2_X1  g238(.A1(new_n437_), .A2(KEYINPUT4), .ZN(new_n440_));
  INV_X1    g239(.A(KEYINPUT95), .ZN(new_n441_));
  NAND2_X1  g240(.A1(new_n370_), .A2(new_n334_), .ZN(new_n442_));
  INV_X1    g241(.A(new_n442_), .ZN(new_n443_));
  NAND3_X1  g242(.A1(new_n440_), .A2(new_n441_), .A3(new_n443_), .ZN(new_n444_));
  OAI21_X1  g243(.A(KEYINPUT95), .B1(new_n369_), .B2(new_n442_), .ZN(new_n445_));
  NAND2_X1  g244(.A1(new_n444_), .A2(new_n445_), .ZN(new_n446_));
  AND3_X1   g245(.A1(new_n439_), .A2(new_n446_), .A3(KEYINPUT96), .ZN(new_n447_));
  AOI21_X1  g246(.A(KEYINPUT96), .B1(new_n439_), .B2(new_n446_), .ZN(new_n448_));
  INV_X1    g247(.A(KEYINPUT33), .ZN(new_n449_));
  NOR2_X1   g248(.A1(new_n381_), .A2(new_n449_), .ZN(new_n450_));
  AOI211_X1 g249(.A(KEYINPUT33), .B(new_n377_), .C1(new_n372_), .C2(new_n378_), .ZN(new_n451_));
  OAI22_X1  g250(.A1(new_n447_), .A2(new_n448_), .B1(new_n450_), .B2(new_n451_), .ZN(new_n452_));
  OAI21_X1  g251(.A(new_n433_), .B1(new_n452_), .B2(new_n292_), .ZN(new_n453_));
  NAND2_X1  g252(.A1(new_n453_), .A2(new_n426_), .ZN(new_n454_));
  INV_X1    g253(.A(new_n385_), .ZN(new_n455_));
  AOI21_X1  g254(.A(new_n276_), .B1(new_n271_), .B2(new_n282_), .ZN(new_n456_));
  NOR3_X1   g255(.A1(new_n289_), .A2(new_n290_), .A3(new_n284_), .ZN(new_n457_));
  OAI21_X1  g256(.A(new_n293_), .B1(new_n456_), .B2(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n302_), .A2(new_n283_), .ZN(new_n459_));
  NAND4_X1  g258(.A1(new_n455_), .A2(new_n458_), .A3(new_n425_), .A4(new_n459_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n454_), .A2(new_n460_), .ZN(new_n461_));
  AOI21_X1  g260(.A(new_n427_), .B1(new_n461_), .B2(new_n332_), .ZN(new_n462_));
  INV_X1    g261(.A(KEYINPUT77), .ZN(new_n463_));
  NAND2_X1  g262(.A1(G229gat), .A2(G233gat), .ZN(new_n464_));
  INV_X1    g263(.A(KEYINPUT75), .ZN(new_n465_));
  XOR2_X1   g264(.A(G1gat), .B(G8gat), .Z(new_n466_));
  INV_X1    g265(.A(new_n466_), .ZN(new_n467_));
  XNOR2_X1  g266(.A(G15gat), .B(G22gat), .ZN(new_n468_));
  INV_X1    g267(.A(KEYINPUT73), .ZN(new_n469_));
  INV_X1    g268(.A(G1gat), .ZN(new_n470_));
  INV_X1    g269(.A(G8gat), .ZN(new_n471_));
  OAI21_X1  g270(.A(KEYINPUT14), .B1(new_n470_), .B2(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n468_), .A2(new_n469_), .A3(new_n472_), .ZN(new_n473_));
  INV_X1    g272(.A(new_n473_), .ZN(new_n474_));
  AOI21_X1  g273(.A(new_n469_), .B1(new_n468_), .B2(new_n472_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n467_), .B1(new_n474_), .B2(new_n475_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G43gat), .B(G50gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  INV_X1    g277(.A(G36gat), .ZN(new_n479_));
  NAND2_X1  g278(.A1(new_n479_), .A2(G29gat), .ZN(new_n480_));
  INV_X1    g279(.A(G29gat), .ZN(new_n481_));
  NAND2_X1  g280(.A1(new_n481_), .A2(G36gat), .ZN(new_n482_));
  AND3_X1   g281(.A1(new_n480_), .A2(new_n482_), .A3(KEYINPUT71), .ZN(new_n483_));
  AOI21_X1  g282(.A(KEYINPUT71), .B1(new_n480_), .B2(new_n482_), .ZN(new_n484_));
  OAI21_X1  g283(.A(new_n478_), .B1(new_n483_), .B2(new_n484_), .ZN(new_n485_));
  NAND2_X1  g284(.A1(new_n480_), .A2(new_n482_), .ZN(new_n486_));
  INV_X1    g285(.A(KEYINPUT71), .ZN(new_n487_));
  NAND2_X1  g286(.A1(new_n486_), .A2(new_n487_), .ZN(new_n488_));
  NAND3_X1  g287(.A1(new_n480_), .A2(new_n482_), .A3(KEYINPUT71), .ZN(new_n489_));
  NAND3_X1  g288(.A1(new_n488_), .A2(new_n489_), .A3(new_n477_), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n485_), .A2(new_n490_), .ZN(new_n491_));
  AND2_X1   g290(.A1(G15gat), .A2(G22gat), .ZN(new_n492_));
  NOR2_X1   g291(.A1(G15gat), .A2(G22gat), .ZN(new_n493_));
  NOR2_X1   g292(.A1(new_n492_), .A2(new_n493_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT14), .ZN(new_n495_));
  AOI21_X1  g294(.A(new_n495_), .B1(G1gat), .B2(G8gat), .ZN(new_n496_));
  OAI21_X1  g295(.A(KEYINPUT73), .B1(new_n494_), .B2(new_n496_), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n497_), .A2(new_n466_), .A3(new_n473_), .ZN(new_n498_));
  AND3_X1   g297(.A1(new_n476_), .A2(new_n491_), .A3(new_n498_), .ZN(new_n499_));
  AOI21_X1  g298(.A(new_n491_), .B1(new_n498_), .B2(new_n476_), .ZN(new_n500_));
  OAI21_X1  g299(.A(new_n465_), .B1(new_n499_), .B2(new_n500_), .ZN(new_n501_));
  AND3_X1   g300(.A1(new_n497_), .A2(new_n466_), .A3(new_n473_), .ZN(new_n502_));
  AOI21_X1  g301(.A(new_n466_), .B1(new_n497_), .B2(new_n473_), .ZN(new_n503_));
  OAI211_X1 g302(.A(new_n490_), .B(new_n485_), .C1(new_n502_), .C2(new_n503_), .ZN(new_n504_));
  NAND3_X1  g303(.A1(new_n476_), .A2(new_n491_), .A3(new_n498_), .ZN(new_n505_));
  NAND3_X1  g304(.A1(new_n504_), .A2(KEYINPUT75), .A3(new_n505_), .ZN(new_n506_));
  AOI21_X1  g305(.A(new_n464_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n507_));
  NAND2_X1  g306(.A1(new_n476_), .A2(new_n498_), .ZN(new_n508_));
  INV_X1    g307(.A(KEYINPUT15), .ZN(new_n509_));
  NAND2_X1  g308(.A1(new_n491_), .A2(new_n509_), .ZN(new_n510_));
  NAND3_X1  g309(.A1(new_n485_), .A2(new_n490_), .A3(KEYINPUT15), .ZN(new_n511_));
  NAND3_X1  g310(.A1(new_n508_), .A2(new_n510_), .A3(new_n511_), .ZN(new_n512_));
  XOR2_X1   g311(.A(new_n464_), .B(KEYINPUT76), .Z(new_n513_));
  NAND3_X1  g312(.A1(new_n512_), .A2(new_n505_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(new_n514_), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n463_), .B1(new_n507_), .B2(new_n515_), .ZN(new_n516_));
  XNOR2_X1  g315(.A(G113gat), .B(G141gat), .ZN(new_n517_));
  XNOR2_X1  g316(.A(G169gat), .B(G197gat), .ZN(new_n518_));
  XOR2_X1   g317(.A(new_n517_), .B(new_n518_), .Z(new_n519_));
  INV_X1    g318(.A(new_n519_), .ZN(new_n520_));
  NAND2_X1  g319(.A1(new_n516_), .A2(new_n520_), .ZN(new_n521_));
  OAI211_X1 g320(.A(new_n463_), .B(new_n519_), .C1(new_n507_), .C2(new_n515_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n521_), .A2(new_n522_), .ZN(new_n523_));
  NOR2_X1   g322(.A1(new_n462_), .A2(new_n523_), .ZN(new_n524_));
  INV_X1    g323(.A(G85gat), .ZN(new_n525_));
  INV_X1    g324(.A(G92gat), .ZN(new_n526_));
  NAND2_X1  g325(.A1(new_n525_), .A2(new_n526_), .ZN(new_n527_));
  NAND2_X1  g326(.A1(G85gat), .A2(G92gat), .ZN(new_n528_));
  AND2_X1   g327(.A1(new_n527_), .A2(new_n528_), .ZN(new_n529_));
  NAND2_X1  g328(.A1(new_n529_), .A2(KEYINPUT9), .ZN(new_n530_));
  XOR2_X1   g329(.A(KEYINPUT10), .B(G99gat), .Z(new_n531_));
  INV_X1    g330(.A(G106gat), .ZN(new_n532_));
  NAND2_X1  g331(.A1(new_n531_), .A2(new_n532_), .ZN(new_n533_));
  NAND2_X1  g332(.A1(G99gat), .A2(G106gat), .ZN(new_n534_));
  INV_X1    g333(.A(KEYINPUT6), .ZN(new_n535_));
  NAND2_X1  g334(.A1(new_n534_), .A2(new_n535_), .ZN(new_n536_));
  NAND3_X1  g335(.A1(KEYINPUT6), .A2(G99gat), .A3(G106gat), .ZN(new_n537_));
  AND2_X1   g336(.A1(new_n536_), .A2(new_n537_), .ZN(new_n538_));
  OR2_X1    g337(.A1(new_n528_), .A2(KEYINPUT9), .ZN(new_n539_));
  NAND4_X1  g338(.A1(new_n530_), .A2(new_n533_), .A3(new_n538_), .A4(new_n539_), .ZN(new_n540_));
  INV_X1    g339(.A(KEYINPUT8), .ZN(new_n541_));
  NAND3_X1  g340(.A1(new_n527_), .A2(new_n541_), .A3(new_n528_), .ZN(new_n542_));
  INV_X1    g341(.A(KEYINPUT7), .ZN(new_n543_));
  NAND3_X1  g342(.A1(new_n543_), .A2(new_n308_), .A3(new_n532_), .ZN(new_n544_));
  OAI21_X1  g343(.A(KEYINPUT7), .B1(G99gat), .B2(G106gat), .ZN(new_n545_));
  NAND4_X1  g344(.A1(new_n544_), .A2(new_n536_), .A3(new_n545_), .A4(new_n537_), .ZN(new_n546_));
  AOI21_X1  g345(.A(new_n542_), .B1(new_n546_), .B2(KEYINPUT64), .ZN(new_n547_));
  AND2_X1   g346(.A1(new_n544_), .A2(new_n545_), .ZN(new_n548_));
  INV_X1    g347(.A(KEYINPUT64), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n548_), .A2(new_n538_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n547_), .A2(new_n550_), .ZN(new_n551_));
  INV_X1    g350(.A(new_n551_), .ZN(new_n552_));
  XNOR2_X1  g351(.A(KEYINPUT65), .B(KEYINPUT6), .ZN(new_n553_));
  NAND2_X1  g352(.A1(new_n553_), .A2(new_n534_), .ZN(new_n554_));
  INV_X1    g353(.A(new_n534_), .ZN(new_n555_));
  INV_X1    g354(.A(KEYINPUT65), .ZN(new_n556_));
  NOR2_X1   g355(.A1(new_n556_), .A2(KEYINPUT6), .ZN(new_n557_));
  NOR2_X1   g356(.A1(new_n535_), .A2(KEYINPUT65), .ZN(new_n558_));
  OAI21_X1  g357(.A(new_n555_), .B1(new_n557_), .B2(new_n558_), .ZN(new_n559_));
  NAND3_X1  g358(.A1(new_n548_), .A2(new_n554_), .A3(new_n559_), .ZN(new_n560_));
  AOI21_X1  g359(.A(new_n541_), .B1(new_n560_), .B2(new_n529_), .ZN(new_n561_));
  OAI211_X1 g360(.A(new_n491_), .B(new_n540_), .C1(new_n552_), .C2(new_n561_), .ZN(new_n562_));
  NAND2_X1  g361(.A1(G232gat), .A2(G233gat), .ZN(new_n563_));
  XNOR2_X1  g362(.A(new_n563_), .B(KEYINPUT34), .ZN(new_n564_));
  OR2_X1    g363(.A1(new_n564_), .A2(KEYINPUT35), .ZN(new_n565_));
  INV_X1    g364(.A(new_n540_), .ZN(new_n566_));
  OAI211_X1 g365(.A(new_n544_), .B(new_n545_), .C1(new_n553_), .C2(new_n534_), .ZN(new_n567_));
  NOR3_X1   g366(.A1(new_n557_), .A2(new_n558_), .A3(new_n555_), .ZN(new_n568_));
  OAI21_X1  g367(.A(new_n529_), .B1(new_n567_), .B2(new_n568_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT8), .ZN(new_n570_));
  AOI21_X1  g369(.A(new_n566_), .B1(new_n570_), .B2(new_n551_), .ZN(new_n571_));
  NAND2_X1  g370(.A1(new_n510_), .A2(new_n511_), .ZN(new_n572_));
  OAI211_X1 g371(.A(new_n562_), .B(new_n565_), .C1(new_n571_), .C2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n564_), .A2(KEYINPUT35), .ZN(new_n574_));
  XOR2_X1   g373(.A(new_n574_), .B(KEYINPUT70), .Z(new_n575_));
  INV_X1    g374(.A(new_n575_), .ZN(new_n576_));
  NAND2_X1  g375(.A1(new_n573_), .A2(new_n576_), .ZN(new_n577_));
  OAI21_X1  g376(.A(new_n540_), .B1(new_n552_), .B2(new_n561_), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n578_), .A2(new_n511_), .A3(new_n510_), .ZN(new_n579_));
  NAND4_X1  g378(.A1(new_n579_), .A2(new_n562_), .A3(new_n565_), .A4(new_n575_), .ZN(new_n580_));
  NAND3_X1  g379(.A1(new_n577_), .A2(new_n580_), .A3(KEYINPUT72), .ZN(new_n581_));
  XNOR2_X1  g380(.A(G190gat), .B(G218gat), .ZN(new_n582_));
  XNOR2_X1  g381(.A(G134gat), .B(G162gat), .ZN(new_n583_));
  XNOR2_X1  g382(.A(new_n582_), .B(new_n583_), .ZN(new_n584_));
  NOR2_X1   g383(.A1(new_n584_), .A2(KEYINPUT36), .ZN(new_n585_));
  INV_X1    g384(.A(new_n585_), .ZN(new_n586_));
  NAND2_X1  g385(.A1(new_n581_), .A2(new_n586_), .ZN(new_n587_));
  NAND4_X1  g386(.A1(new_n577_), .A2(new_n580_), .A3(KEYINPUT72), .A4(new_n585_), .ZN(new_n588_));
  NAND2_X1  g387(.A1(new_n587_), .A2(new_n588_), .ZN(new_n589_));
  INV_X1    g388(.A(KEYINPUT37), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n577_), .A2(new_n580_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n591_), .A2(KEYINPUT36), .A3(new_n584_), .ZN(new_n592_));
  AND3_X1   g391(.A1(new_n589_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n593_));
  AOI21_X1  g392(.A(new_n590_), .B1(new_n589_), .B2(new_n592_), .ZN(new_n594_));
  NOR2_X1   g393(.A1(new_n593_), .A2(new_n594_), .ZN(new_n595_));
  XNOR2_X1  g394(.A(G57gat), .B(G64gat), .ZN(new_n596_));
  NAND2_X1  g395(.A1(new_n596_), .A2(KEYINPUT11), .ZN(new_n597_));
  XOR2_X1   g396(.A(G71gat), .B(G78gat), .Z(new_n598_));
  NOR2_X1   g397(.A1(new_n597_), .A2(new_n598_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n599_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n596_), .A2(KEYINPUT11), .ZN(new_n601_));
  NAND2_X1  g400(.A1(new_n597_), .A2(new_n598_), .ZN(new_n602_));
  OAI21_X1  g401(.A(new_n600_), .B1(new_n601_), .B2(new_n602_), .ZN(new_n603_));
  NAND2_X1  g402(.A1(G231gat), .A2(G233gat), .ZN(new_n604_));
  XNOR2_X1  g403(.A(new_n603_), .B(new_n604_), .ZN(new_n605_));
  XNOR2_X1  g404(.A(new_n605_), .B(new_n508_), .ZN(new_n606_));
  INV_X1    g405(.A(KEYINPUT74), .ZN(new_n607_));
  OR2_X1    g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  XNOR2_X1  g407(.A(G127gat), .B(G155gat), .ZN(new_n609_));
  XNOR2_X1  g408(.A(new_n609_), .B(KEYINPUT16), .ZN(new_n610_));
  XNOR2_X1  g409(.A(G183gat), .B(G211gat), .ZN(new_n611_));
  XNOR2_X1  g410(.A(new_n610_), .B(new_n611_), .ZN(new_n612_));
  NAND2_X1  g411(.A1(new_n608_), .A2(new_n612_), .ZN(new_n613_));
  OAI21_X1  g412(.A(KEYINPUT17), .B1(new_n606_), .B2(new_n612_), .ZN(new_n614_));
  NAND2_X1  g413(.A1(new_n613_), .A2(new_n614_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n608_), .A2(KEYINPUT17), .A3(new_n612_), .ZN(new_n616_));
  NAND2_X1  g415(.A1(new_n615_), .A2(new_n616_), .ZN(new_n617_));
  NAND2_X1  g416(.A1(new_n595_), .A2(new_n617_), .ZN(new_n618_));
  INV_X1    g417(.A(new_n603_), .ZN(new_n619_));
  AOI22_X1  g418(.A1(new_n569_), .A2(KEYINPUT8), .B1(new_n550_), .B2(new_n547_), .ZN(new_n620_));
  OAI21_X1  g419(.A(new_n619_), .B1(new_n620_), .B2(new_n566_), .ZN(new_n621_));
  OAI211_X1 g420(.A(new_n603_), .B(new_n540_), .C1(new_n552_), .C2(new_n561_), .ZN(new_n622_));
  NAND3_X1  g421(.A1(new_n621_), .A2(KEYINPUT12), .A3(new_n622_), .ZN(new_n623_));
  INV_X1    g422(.A(KEYINPUT12), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n578_), .A2(new_n624_), .A3(new_n619_), .ZN(new_n625_));
  NAND2_X1  g424(.A1(new_n623_), .A2(new_n625_), .ZN(new_n626_));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627_));
  NAND2_X1  g426(.A1(new_n626_), .A2(new_n627_), .ZN(new_n628_));
  NAND2_X1  g427(.A1(new_n621_), .A2(new_n622_), .ZN(new_n629_));
  NAND3_X1  g428(.A1(new_n629_), .A2(G230gat), .A3(G233gat), .ZN(new_n630_));
  NAND2_X1  g429(.A1(new_n628_), .A2(new_n630_), .ZN(new_n631_));
  XOR2_X1   g430(.A(G120gat), .B(G148gat), .Z(new_n632_));
  XNOR2_X1  g431(.A(G176gat), .B(G204gat), .ZN(new_n633_));
  XNOR2_X1  g432(.A(new_n632_), .B(new_n633_), .ZN(new_n634_));
  XNOR2_X1  g433(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n635_));
  XNOR2_X1  g434(.A(new_n634_), .B(new_n635_), .ZN(new_n636_));
  NAND2_X1  g435(.A1(new_n636_), .A2(KEYINPUT66), .ZN(new_n637_));
  XOR2_X1   g436(.A(new_n637_), .B(KEYINPUT68), .Z(new_n638_));
  INV_X1    g437(.A(new_n638_), .ZN(new_n639_));
  NAND2_X1  g438(.A1(new_n631_), .A2(new_n639_), .ZN(new_n640_));
  NAND3_X1  g439(.A1(new_n638_), .A2(new_n628_), .A3(new_n630_), .ZN(new_n641_));
  NAND2_X1  g440(.A1(new_n640_), .A2(new_n641_), .ZN(new_n642_));
  INV_X1    g441(.A(KEYINPUT13), .ZN(new_n643_));
  NAND2_X1  g442(.A1(new_n642_), .A2(new_n643_), .ZN(new_n644_));
  NAND3_X1  g443(.A1(new_n640_), .A2(new_n641_), .A3(KEYINPUT13), .ZN(new_n645_));
  AND2_X1   g444(.A1(new_n644_), .A2(new_n645_), .ZN(new_n646_));
  OR2_X1    g445(.A1(new_n646_), .A2(KEYINPUT69), .ZN(new_n647_));
  NAND2_X1  g446(.A1(new_n646_), .A2(KEYINPUT69), .ZN(new_n648_));
  AOI21_X1  g447(.A(new_n618_), .B1(new_n647_), .B2(new_n648_), .ZN(new_n649_));
  NAND4_X1  g448(.A1(new_n524_), .A2(new_n470_), .A3(new_n385_), .A4(new_n649_), .ZN(new_n650_));
  INV_X1    g449(.A(KEYINPUT38), .ZN(new_n651_));
  NOR2_X1   g450(.A1(new_n650_), .A2(new_n651_), .ZN(new_n652_));
  XNOR2_X1  g451(.A(new_n652_), .B(KEYINPUT101), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n650_), .A2(new_n651_), .ZN(new_n654_));
  NAND2_X1  g453(.A1(new_n458_), .A2(new_n459_), .ZN(new_n655_));
  NOR2_X1   g454(.A1(new_n655_), .A2(new_n425_), .ZN(new_n656_));
  NAND2_X1  g455(.A1(new_n656_), .A2(new_n386_), .ZN(new_n657_));
  AND2_X1   g456(.A1(new_n420_), .A2(new_n421_), .ZN(new_n658_));
  INV_X1    g457(.A(new_n424_), .ZN(new_n659_));
  NAND2_X1  g458(.A1(new_n658_), .A2(new_n659_), .ZN(new_n660_));
  AOI21_X1  g459(.A(new_n385_), .B1(new_n660_), .B2(new_n416_), .ZN(new_n661_));
  AOI22_X1  g460(.A1(new_n661_), .A2(new_n303_), .B1(new_n453_), .B2(new_n426_), .ZN(new_n662_));
  OAI21_X1  g461(.A(new_n657_), .B1(new_n662_), .B2(new_n331_), .ZN(new_n663_));
  NAND2_X1  g462(.A1(new_n589_), .A2(new_n592_), .ZN(new_n664_));
  INV_X1    g463(.A(new_n664_), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n644_), .A2(new_n645_), .ZN(new_n666_));
  AND2_X1   g465(.A1(new_n615_), .A2(new_n616_), .ZN(new_n667_));
  NOR3_X1   g466(.A1(new_n666_), .A2(new_n667_), .A3(new_n523_), .ZN(new_n668_));
  NAND3_X1  g467(.A1(new_n663_), .A2(new_n665_), .A3(new_n668_), .ZN(new_n669_));
  OAI21_X1  g468(.A(G1gat), .B1(new_n669_), .B2(new_n455_), .ZN(new_n670_));
  NAND3_X1  g469(.A1(new_n653_), .A2(new_n654_), .A3(new_n670_), .ZN(G1324gat));
  XNOR2_X1  g470(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n672_));
  NOR2_X1   g471(.A1(new_n303_), .A2(G8gat), .ZN(new_n673_));
  NAND3_X1  g472(.A1(new_n524_), .A2(new_n649_), .A3(new_n673_), .ZN(new_n674_));
  XNOR2_X1  g473(.A(new_n674_), .B(KEYINPUT102), .ZN(new_n675_));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n676_));
  OAI21_X1  g475(.A(new_n676_), .B1(new_n669_), .B2(new_n303_), .ZN(new_n677_));
  NOR2_X1   g476(.A1(new_n462_), .A2(new_n664_), .ZN(new_n678_));
  NAND4_X1  g477(.A1(new_n678_), .A2(KEYINPUT103), .A3(new_n655_), .A4(new_n668_), .ZN(new_n679_));
  NAND4_X1  g478(.A1(new_n677_), .A2(new_n679_), .A3(KEYINPUT39), .A4(G8gat), .ZN(new_n680_));
  AND2_X1   g479(.A1(new_n675_), .A2(new_n680_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n677_), .A2(new_n679_), .A3(G8gat), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT39), .ZN(new_n683_));
  NAND2_X1  g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  AOI21_X1  g483(.A(new_n672_), .B1(new_n681_), .B2(new_n684_), .ZN(new_n685_));
  AND4_X1   g484(.A1(new_n684_), .A2(new_n675_), .A3(new_n680_), .A4(new_n672_), .ZN(new_n686_));
  NOR2_X1   g485(.A1(new_n685_), .A2(new_n686_), .ZN(G1325gat));
  OAI21_X1  g486(.A(G15gat), .B1(new_n669_), .B2(new_n332_), .ZN(new_n688_));
  XNOR2_X1  g487(.A(new_n688_), .B(KEYINPUT41), .ZN(new_n689_));
  NAND2_X1  g488(.A1(new_n524_), .A2(new_n649_), .ZN(new_n690_));
  NOR3_X1   g489(.A1(new_n690_), .A2(G15gat), .A3(new_n332_), .ZN(new_n691_));
  OR2_X1    g490(.A1(new_n689_), .A2(new_n691_), .ZN(G1326gat));
  OAI21_X1  g491(.A(G22gat), .B1(new_n669_), .B2(new_n426_), .ZN(new_n693_));
  XNOR2_X1  g492(.A(new_n693_), .B(KEYINPUT42), .ZN(new_n694_));
  OR2_X1    g493(.A1(new_n426_), .A2(G22gat), .ZN(new_n695_));
  OAI21_X1  g494(.A(new_n694_), .B1(new_n690_), .B2(new_n695_), .ZN(G1327gat));
  NOR3_X1   g495(.A1(new_n666_), .A2(new_n617_), .A3(new_n665_), .ZN(new_n697_));
  NAND2_X1  g496(.A1(new_n524_), .A2(new_n697_), .ZN(new_n698_));
  INV_X1    g497(.A(new_n698_), .ZN(new_n699_));
  AOI21_X1  g498(.A(G29gat), .B1(new_n699_), .B2(new_n385_), .ZN(new_n700_));
  OAI21_X1  g499(.A(KEYINPUT106), .B1(KEYINPUT105), .B2(KEYINPUT44), .ZN(new_n701_));
  INV_X1    g500(.A(new_n701_), .ZN(new_n702_));
  INV_X1    g501(.A(KEYINPUT43), .ZN(new_n703_));
  NAND2_X1  g502(.A1(new_n664_), .A2(KEYINPUT37), .ZN(new_n704_));
  NAND3_X1  g503(.A1(new_n589_), .A2(new_n590_), .A3(new_n592_), .ZN(new_n705_));
  NAND2_X1  g504(.A1(new_n704_), .A2(new_n705_), .ZN(new_n706_));
  AOI21_X1  g505(.A(new_n703_), .B1(new_n663_), .B2(new_n706_), .ZN(new_n707_));
  AOI21_X1  g506(.A(new_n331_), .B1(new_n454_), .B2(new_n460_), .ZN(new_n708_));
  OAI211_X1 g507(.A(new_n703_), .B(new_n706_), .C1(new_n708_), .C2(new_n427_), .ZN(new_n709_));
  INV_X1    g508(.A(new_n709_), .ZN(new_n710_));
  NOR2_X1   g509(.A1(new_n707_), .A2(new_n710_), .ZN(new_n711_));
  NOR2_X1   g510(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n712_));
  NOR2_X1   g511(.A1(new_n617_), .A2(new_n712_), .ZN(new_n713_));
  INV_X1    g512(.A(new_n523_), .ZN(new_n714_));
  NAND3_X1  g513(.A1(new_n713_), .A2(new_n646_), .A3(new_n714_), .ZN(new_n715_));
  OAI21_X1  g514(.A(new_n702_), .B1(new_n711_), .B2(new_n715_), .ZN(new_n716_));
  OAI21_X1  g515(.A(KEYINPUT43), .B1(new_n462_), .B2(new_n595_), .ZN(new_n717_));
  NAND2_X1  g516(.A1(new_n717_), .A2(new_n709_), .ZN(new_n718_));
  INV_X1    g517(.A(new_n715_), .ZN(new_n719_));
  NAND3_X1  g518(.A1(new_n718_), .A2(new_n719_), .A3(new_n701_), .ZN(new_n720_));
  NAND2_X1  g519(.A1(new_n716_), .A2(new_n720_), .ZN(new_n721_));
  NOR2_X1   g520(.A1(new_n455_), .A2(new_n481_), .ZN(new_n722_));
  AOI21_X1  g521(.A(new_n700_), .B1(new_n721_), .B2(new_n722_), .ZN(G1328gat));
  AND4_X1   g522(.A1(new_n479_), .A2(new_n524_), .A3(new_n655_), .A4(new_n697_), .ZN(new_n724_));
  XNOR2_X1  g523(.A(KEYINPUT107), .B(KEYINPUT45), .ZN(new_n725_));
  XNOR2_X1  g524(.A(new_n724_), .B(new_n725_), .ZN(new_n726_));
  AOI21_X1  g525(.A(new_n303_), .B1(new_n716_), .B2(new_n720_), .ZN(new_n727_));
  OAI21_X1  g526(.A(new_n726_), .B1(new_n727_), .B2(new_n479_), .ZN(new_n728_));
  INV_X1    g527(.A(KEYINPUT46), .ZN(new_n729_));
  NAND2_X1  g528(.A1(new_n728_), .A2(new_n729_), .ZN(new_n730_));
  OAI211_X1 g529(.A(new_n726_), .B(KEYINPUT46), .C1(new_n727_), .C2(new_n479_), .ZN(new_n731_));
  NAND2_X1  g530(.A1(new_n730_), .A2(new_n731_), .ZN(G1329gat));
  INV_X1    g531(.A(KEYINPUT47), .ZN(new_n733_));
  AOI21_X1  g532(.A(new_n701_), .B1(new_n718_), .B2(new_n719_), .ZN(new_n734_));
  AOI211_X1 g533(.A(new_n715_), .B(new_n702_), .C1(new_n717_), .C2(new_n709_), .ZN(new_n735_));
  OAI21_X1  g534(.A(new_n331_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n736_));
  NAND2_X1  g535(.A1(new_n736_), .A2(G43gat), .ZN(new_n737_));
  NOR3_X1   g536(.A1(new_n698_), .A2(G43gat), .A3(new_n332_), .ZN(new_n738_));
  INV_X1    g537(.A(new_n738_), .ZN(new_n739_));
  AOI21_X1  g538(.A(new_n733_), .B1(new_n737_), .B2(new_n739_), .ZN(new_n740_));
  AOI211_X1 g539(.A(KEYINPUT47), .B(new_n738_), .C1(new_n736_), .C2(G43gat), .ZN(new_n741_));
  NOR2_X1   g540(.A1(new_n740_), .A2(new_n741_), .ZN(G1330gat));
  OR3_X1    g541(.A1(new_n698_), .A2(G50gat), .A3(new_n426_), .ZN(new_n743_));
  OAI21_X1  g542(.A(new_n425_), .B1(new_n734_), .B2(new_n735_), .ZN(new_n744_));
  INV_X1    g543(.A(KEYINPUT108), .ZN(new_n745_));
  AND3_X1   g544(.A1(new_n744_), .A2(new_n745_), .A3(G50gat), .ZN(new_n746_));
  AOI21_X1  g545(.A(new_n745_), .B1(new_n744_), .B2(G50gat), .ZN(new_n747_));
  OAI21_X1  g546(.A(new_n743_), .B1(new_n746_), .B2(new_n747_), .ZN(G1331gat));
  AND2_X1   g547(.A1(new_n647_), .A2(new_n648_), .ZN(new_n749_));
  NAND4_X1  g548(.A1(new_n678_), .A2(new_n523_), .A3(new_n749_), .A4(new_n617_), .ZN(new_n750_));
  INV_X1    g549(.A(G57gat), .ZN(new_n751_));
  NOR3_X1   g550(.A1(new_n750_), .A2(new_n751_), .A3(new_n455_), .ZN(new_n752_));
  NOR2_X1   g551(.A1(new_n706_), .A2(new_n667_), .ZN(new_n753_));
  NAND2_X1  g552(.A1(new_n753_), .A2(new_n666_), .ZN(new_n754_));
  XNOR2_X1  g553(.A(new_n754_), .B(KEYINPUT109), .ZN(new_n755_));
  NAND3_X1  g554(.A1(new_n755_), .A2(new_n663_), .A3(new_n523_), .ZN(new_n756_));
  OR2_X1    g555(.A1(new_n756_), .A2(KEYINPUT110), .ZN(new_n757_));
  NAND2_X1  g556(.A1(new_n756_), .A2(KEYINPUT110), .ZN(new_n758_));
  NAND3_X1  g557(.A1(new_n757_), .A2(new_n385_), .A3(new_n758_), .ZN(new_n759_));
  AOI21_X1  g558(.A(new_n752_), .B1(new_n759_), .B2(new_n751_), .ZN(G1332gat));
  OR3_X1    g559(.A1(new_n756_), .A2(G64gat), .A3(new_n303_), .ZN(new_n761_));
  OAI21_X1  g560(.A(G64gat), .B1(new_n750_), .B2(new_n303_), .ZN(new_n762_));
  OR2_X1    g561(.A1(new_n762_), .A2(KEYINPUT48), .ZN(new_n763_));
  INV_X1    g562(.A(new_n763_), .ZN(new_n764_));
  AND2_X1   g563(.A1(new_n762_), .A2(KEYINPUT48), .ZN(new_n765_));
  OAI21_X1  g564(.A(new_n761_), .B1(new_n764_), .B2(new_n765_), .ZN(G1333gat));
  OR3_X1    g565(.A1(new_n756_), .A2(G71gat), .A3(new_n332_), .ZN(new_n767_));
  OR2_X1    g566(.A1(new_n750_), .A2(new_n332_), .ZN(new_n768_));
  XOR2_X1   g567(.A(KEYINPUT111), .B(KEYINPUT49), .Z(new_n769_));
  NAND3_X1  g568(.A1(new_n768_), .A2(G71gat), .A3(new_n769_), .ZN(new_n770_));
  INV_X1    g569(.A(new_n770_), .ZN(new_n771_));
  AOI21_X1  g570(.A(new_n769_), .B1(new_n768_), .B2(G71gat), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n767_), .B1(new_n771_), .B2(new_n772_), .ZN(G1334gat));
  OR3_X1    g572(.A1(new_n756_), .A2(G78gat), .A3(new_n426_), .ZN(new_n774_));
  OAI21_X1  g573(.A(G78gat), .B1(new_n750_), .B2(new_n426_), .ZN(new_n775_));
  OR2_X1    g574(.A1(new_n775_), .A2(KEYINPUT50), .ZN(new_n776_));
  INV_X1    g575(.A(new_n776_), .ZN(new_n777_));
  AND2_X1   g576(.A1(new_n775_), .A2(KEYINPUT50), .ZN(new_n778_));
  OAI21_X1  g577(.A(new_n774_), .B1(new_n777_), .B2(new_n778_), .ZN(G1335gat));
  NOR2_X1   g578(.A1(new_n617_), .A2(new_n665_), .ZN(new_n780_));
  NAND4_X1  g579(.A1(new_n749_), .A2(new_n663_), .A3(new_n523_), .A4(new_n780_), .ZN(new_n781_));
  OR2_X1    g580(.A1(new_n781_), .A2(KEYINPUT112), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(KEYINPUT112), .ZN(new_n783_));
  NAND2_X1  g582(.A1(new_n782_), .A2(new_n783_), .ZN(new_n784_));
  NAND3_X1  g583(.A1(new_n784_), .A2(new_n525_), .A3(new_n385_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n667_), .A2(new_n666_), .A3(new_n523_), .ZN(new_n786_));
  AOI21_X1  g585(.A(new_n786_), .B1(new_n717_), .B2(new_n709_), .ZN(new_n787_));
  INV_X1    g586(.A(new_n787_), .ZN(new_n788_));
  OAI21_X1  g587(.A(G85gat), .B1(new_n788_), .B2(new_n455_), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n785_), .A2(new_n789_), .ZN(G1336gat));
  NAND3_X1  g589(.A1(new_n784_), .A2(new_n526_), .A3(new_n655_), .ZN(new_n791_));
  OAI21_X1  g590(.A(G92gat), .B1(new_n788_), .B2(new_n303_), .ZN(new_n792_));
  NAND2_X1  g591(.A1(new_n791_), .A2(new_n792_), .ZN(G1337gat));
  NAND2_X1  g592(.A1(new_n331_), .A2(new_n531_), .ZN(new_n794_));
  AOI21_X1  g593(.A(new_n794_), .B1(new_n782_), .B2(new_n783_), .ZN(new_n795_));
  AOI21_X1  g594(.A(new_n308_), .B1(new_n787_), .B2(new_n331_), .ZN(new_n796_));
  INV_X1    g595(.A(KEYINPUT113), .ZN(new_n797_));
  OAI22_X1  g596(.A1(new_n795_), .A2(new_n796_), .B1(new_n797_), .B2(KEYINPUT51), .ZN(new_n798_));
  NAND2_X1  g597(.A1(new_n797_), .A2(KEYINPUT51), .ZN(new_n799_));
  XNOR2_X1  g598(.A(new_n798_), .B(new_n799_), .ZN(G1338gat));
  NAND3_X1  g599(.A1(new_n784_), .A2(new_n532_), .A3(new_n425_), .ZN(new_n801_));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802_));
  NAND2_X1  g601(.A1(new_n787_), .A2(new_n425_), .ZN(new_n803_));
  AOI21_X1  g602(.A(new_n802_), .B1(new_n803_), .B2(G106gat), .ZN(new_n804_));
  AOI211_X1 g603(.A(KEYINPUT52), .B(new_n532_), .C1(new_n787_), .C2(new_n425_), .ZN(new_n805_));
  OAI21_X1  g604(.A(new_n801_), .B1(new_n804_), .B2(new_n805_), .ZN(new_n806_));
  NAND2_X1  g605(.A1(new_n806_), .A2(KEYINPUT53), .ZN(new_n807_));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n808_));
  OAI211_X1 g607(.A(new_n801_), .B(new_n808_), .C1(new_n804_), .C2(new_n805_), .ZN(new_n809_));
  NAND2_X1  g608(.A1(new_n807_), .A2(new_n809_), .ZN(G1339gat));
  NOR2_X1   g609(.A1(new_n455_), .A2(new_n332_), .ZN(new_n811_));
  NAND2_X1  g610(.A1(new_n656_), .A2(new_n811_), .ZN(new_n812_));
  INV_X1    g611(.A(new_n636_), .ZN(new_n813_));
  NAND3_X1  g612(.A1(new_n628_), .A2(new_n630_), .A3(new_n813_), .ZN(new_n814_));
  AND3_X1   g613(.A1(new_n521_), .A2(new_n814_), .A3(new_n522_), .ZN(new_n815_));
  NAND2_X1  g614(.A1(new_n626_), .A2(KEYINPUT55), .ZN(new_n816_));
  NAND3_X1  g615(.A1(KEYINPUT114), .A2(G230gat), .A3(G233gat), .ZN(new_n817_));
  AOI22_X1  g616(.A1(new_n623_), .A2(new_n625_), .B1(G230gat), .B2(G233gat), .ZN(new_n818_));
  OAI211_X1 g617(.A(new_n816_), .B(new_n817_), .C1(KEYINPUT55), .C2(new_n818_), .ZN(new_n819_));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820_));
  AOI21_X1  g619(.A(new_n820_), .B1(new_n623_), .B2(new_n625_), .ZN(new_n821_));
  INV_X1    g620(.A(new_n817_), .ZN(new_n822_));
  AOI21_X1  g621(.A(new_n813_), .B1(new_n821_), .B2(new_n822_), .ZN(new_n823_));
  AND3_X1   g622(.A1(new_n819_), .A2(KEYINPUT56), .A3(new_n823_), .ZN(new_n824_));
  AOI21_X1  g623(.A(KEYINPUT56), .B1(new_n819_), .B2(new_n823_), .ZN(new_n825_));
  OAI21_X1  g624(.A(new_n815_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n826_));
  AND3_X1   g625(.A1(new_n504_), .A2(KEYINPUT75), .A3(new_n505_), .ZN(new_n827_));
  AOI21_X1  g626(.A(KEYINPUT75), .B1(new_n504_), .B2(new_n505_), .ZN(new_n828_));
  OAI21_X1  g627(.A(new_n513_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n829_));
  INV_X1    g628(.A(new_n513_), .ZN(new_n830_));
  NAND3_X1  g629(.A1(new_n512_), .A2(new_n505_), .A3(new_n830_), .ZN(new_n831_));
  AOI21_X1  g630(.A(new_n519_), .B1(new_n829_), .B2(new_n831_), .ZN(new_n832_));
  INV_X1    g631(.A(new_n464_), .ZN(new_n833_));
  OAI21_X1  g632(.A(new_n833_), .B1(new_n827_), .B2(new_n828_), .ZN(new_n834_));
  AOI21_X1  g633(.A(new_n520_), .B1(new_n834_), .B2(new_n514_), .ZN(new_n835_));
  OAI21_X1  g634(.A(KEYINPUT115), .B1(new_n832_), .B2(new_n835_), .ZN(new_n836_));
  AOI21_X1  g635(.A(new_n830_), .B1(new_n501_), .B2(new_n506_), .ZN(new_n837_));
  INV_X1    g636(.A(new_n831_), .ZN(new_n838_));
  OAI21_X1  g637(.A(new_n520_), .B1(new_n837_), .B2(new_n838_), .ZN(new_n839_));
  OAI21_X1  g638(.A(new_n519_), .B1(new_n507_), .B2(new_n515_), .ZN(new_n840_));
  INV_X1    g639(.A(KEYINPUT115), .ZN(new_n841_));
  NAND3_X1  g640(.A1(new_n839_), .A2(new_n840_), .A3(new_n841_), .ZN(new_n842_));
  NAND3_X1  g641(.A1(new_n642_), .A2(new_n836_), .A3(new_n842_), .ZN(new_n843_));
  NAND2_X1  g642(.A1(new_n826_), .A2(new_n843_), .ZN(new_n844_));
  NAND2_X1  g643(.A1(new_n844_), .A2(new_n665_), .ZN(new_n845_));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846_));
  NAND2_X1  g645(.A1(new_n845_), .A2(new_n846_), .ZN(new_n847_));
  NAND3_X1  g646(.A1(new_n844_), .A2(KEYINPUT57), .A3(new_n665_), .ZN(new_n848_));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849_));
  NAND3_X1  g648(.A1(new_n836_), .A2(new_n814_), .A3(new_n842_), .ZN(new_n850_));
  NAND2_X1  g649(.A1(new_n816_), .A2(new_n817_), .ZN(new_n851_));
  AOI21_X1  g650(.A(KEYINPUT55), .B1(new_n626_), .B2(new_n627_), .ZN(new_n852_));
  OAI21_X1  g651(.A(new_n823_), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n854_));
  NAND2_X1  g653(.A1(new_n853_), .A2(new_n854_), .ZN(new_n855_));
  NAND3_X1  g654(.A1(new_n819_), .A2(KEYINPUT56), .A3(new_n823_), .ZN(new_n856_));
  AOI21_X1  g655(.A(new_n850_), .B1(new_n855_), .B2(new_n856_), .ZN(new_n857_));
  OAI211_X1 g656(.A(new_n706_), .B(new_n849_), .C1(new_n857_), .C2(KEYINPUT58), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(KEYINPUT58), .ZN(new_n859_));
  NAND2_X1  g658(.A1(new_n858_), .A2(new_n859_), .ZN(new_n860_));
  AND3_X1   g659(.A1(new_n836_), .A2(new_n814_), .A3(new_n842_), .ZN(new_n861_));
  OAI21_X1  g660(.A(new_n861_), .B1(new_n824_), .B2(new_n825_), .ZN(new_n862_));
  INV_X1    g661(.A(KEYINPUT58), .ZN(new_n863_));
  NAND2_X1  g662(.A1(new_n862_), .A2(new_n863_), .ZN(new_n864_));
  AOI21_X1  g663(.A(new_n849_), .B1(new_n864_), .B2(new_n706_), .ZN(new_n865_));
  OAI211_X1 g664(.A(new_n847_), .B(new_n848_), .C1(new_n860_), .C2(new_n865_), .ZN(new_n866_));
  NAND2_X1  g665(.A1(new_n866_), .A2(new_n667_), .ZN(new_n867_));
  INV_X1    g666(.A(KEYINPUT54), .ZN(new_n868_));
  NAND3_X1  g667(.A1(new_n644_), .A2(new_n523_), .A3(new_n645_), .ZN(new_n869_));
  INV_X1    g668(.A(new_n869_), .ZN(new_n870_));
  AOI21_X1  g669(.A(new_n868_), .B1(new_n753_), .B2(new_n870_), .ZN(new_n871_));
  NOR3_X1   g670(.A1(new_n618_), .A2(KEYINPUT54), .A3(new_n869_), .ZN(new_n872_));
  NOR2_X1   g671(.A1(new_n871_), .A2(new_n872_), .ZN(new_n873_));
  INV_X1    g672(.A(new_n873_), .ZN(new_n874_));
  AOI21_X1  g673(.A(new_n812_), .B1(new_n867_), .B2(new_n874_), .ZN(new_n875_));
  INV_X1    g674(.A(KEYINPUT59), .ZN(new_n876_));
  OAI21_X1  g675(.A(KEYINPUT117), .B1(new_n875_), .B2(new_n876_), .ZN(new_n877_));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n878_));
  AOI21_X1  g677(.A(new_n873_), .B1(new_n866_), .B2(new_n667_), .ZN(new_n879_));
  OAI211_X1 g678(.A(new_n878_), .B(KEYINPUT59), .C1(new_n879_), .C2(new_n812_), .ZN(new_n880_));
  NAND2_X1  g679(.A1(new_n877_), .A2(new_n880_), .ZN(new_n881_));
  INV_X1    g680(.A(new_n879_), .ZN(new_n882_));
  INV_X1    g681(.A(new_n812_), .ZN(new_n883_));
  AND2_X1   g682(.A1(new_n883_), .A2(KEYINPUT118), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n883_), .A2(KEYINPUT118), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n884_), .A2(new_n885_), .A3(KEYINPUT59), .ZN(new_n886_));
  NAND2_X1  g685(.A1(new_n882_), .A2(new_n886_), .ZN(new_n887_));
  NAND3_X1  g686(.A1(new_n881_), .A2(new_n714_), .A3(new_n887_), .ZN(new_n888_));
  NAND2_X1  g687(.A1(new_n888_), .A2(G113gat), .ZN(new_n889_));
  AOI21_X1  g688(.A(KEYINPUT57), .B1(new_n844_), .B2(new_n665_), .ZN(new_n890_));
  AOI211_X1 g689(.A(new_n846_), .B(new_n664_), .C1(new_n826_), .C2(new_n843_), .ZN(new_n891_));
  NOR2_X1   g690(.A1(new_n890_), .A2(new_n891_), .ZN(new_n892_));
  NAND2_X1  g691(.A1(new_n855_), .A2(new_n856_), .ZN(new_n893_));
  AOI21_X1  g692(.A(KEYINPUT58), .B1(new_n893_), .B2(new_n861_), .ZN(new_n894_));
  OAI21_X1  g693(.A(KEYINPUT116), .B1(new_n894_), .B2(new_n595_), .ZN(new_n895_));
  NAND3_X1  g694(.A1(new_n895_), .A2(new_n859_), .A3(new_n858_), .ZN(new_n896_));
  AOI21_X1  g695(.A(new_n617_), .B1(new_n892_), .B2(new_n896_), .ZN(new_n897_));
  OAI21_X1  g696(.A(new_n883_), .B1(new_n897_), .B2(new_n873_), .ZN(new_n898_));
  OR3_X1    g697(.A1(new_n898_), .A2(G113gat), .A3(new_n523_), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n889_), .A2(new_n899_), .ZN(G1340gat));
  XOR2_X1   g699(.A(KEYINPUT119), .B(G120gat), .Z(new_n901_));
  INV_X1    g700(.A(new_n901_), .ZN(new_n902_));
  INV_X1    g701(.A(KEYINPUT60), .ZN(new_n903_));
  AOI21_X1  g702(.A(new_n902_), .B1(new_n666_), .B2(new_n903_), .ZN(new_n904_));
  OAI22_X1  g703(.A1(new_n904_), .A2(KEYINPUT120), .B1(KEYINPUT60), .B2(new_n901_), .ZN(new_n905_));
  AOI21_X1  g704(.A(new_n905_), .B1(KEYINPUT120), .B2(new_n904_), .ZN(new_n906_));
  NAND2_X1  g705(.A1(new_n875_), .A2(new_n906_), .ZN(new_n907_));
  INV_X1    g706(.A(new_n749_), .ZN(new_n908_));
  AOI21_X1  g707(.A(new_n908_), .B1(new_n882_), .B2(new_n886_), .ZN(new_n909_));
  INV_X1    g708(.A(new_n880_), .ZN(new_n910_));
  AOI21_X1  g709(.A(new_n878_), .B1(new_n898_), .B2(KEYINPUT59), .ZN(new_n911_));
  OAI211_X1 g710(.A(KEYINPUT121), .B(new_n909_), .C1(new_n910_), .C2(new_n911_), .ZN(new_n912_));
  NAND2_X1  g711(.A1(new_n912_), .A2(new_n902_), .ZN(new_n913_));
  AOI21_X1  g712(.A(KEYINPUT121), .B1(new_n881_), .B2(new_n909_), .ZN(new_n914_));
  OAI21_X1  g713(.A(new_n907_), .B1(new_n913_), .B2(new_n914_), .ZN(G1341gat));
  NAND3_X1  g714(.A1(new_n881_), .A2(new_n617_), .A3(new_n887_), .ZN(new_n916_));
  NAND2_X1  g715(.A1(new_n916_), .A2(G127gat), .ZN(new_n917_));
  OR3_X1    g716(.A1(new_n898_), .A2(G127gat), .A3(new_n667_), .ZN(new_n918_));
  NAND2_X1  g717(.A1(new_n917_), .A2(new_n918_), .ZN(G1342gat));
  NAND3_X1  g718(.A1(new_n881_), .A2(new_n706_), .A3(new_n887_), .ZN(new_n920_));
  NAND2_X1  g719(.A1(new_n920_), .A2(G134gat), .ZN(new_n921_));
  OR3_X1    g720(.A1(new_n898_), .A2(G134gat), .A3(new_n665_), .ZN(new_n922_));
  NAND2_X1  g721(.A1(new_n921_), .A2(new_n922_), .ZN(G1343gat));
  NOR3_X1   g722(.A1(new_n426_), .A2(new_n455_), .A3(new_n331_), .ZN(new_n924_));
  NAND3_X1  g723(.A1(new_n882_), .A2(new_n303_), .A3(new_n924_), .ZN(new_n925_));
  NOR2_X1   g724(.A1(new_n925_), .A2(new_n523_), .ZN(new_n926_));
  XNOR2_X1  g725(.A(new_n926_), .B(new_n338_), .ZN(G1344gat));
  NOR2_X1   g726(.A1(new_n925_), .A2(new_n908_), .ZN(new_n928_));
  XNOR2_X1  g727(.A(new_n928_), .B(new_n339_), .ZN(G1345gat));
  NOR2_X1   g728(.A1(new_n925_), .A2(new_n667_), .ZN(new_n930_));
  XOR2_X1   g729(.A(KEYINPUT61), .B(G155gat), .Z(new_n931_));
  XNOR2_X1  g730(.A(new_n930_), .B(new_n931_), .ZN(G1346gat));
  OAI21_X1  g731(.A(G162gat), .B1(new_n925_), .B2(new_n595_), .ZN(new_n933_));
  OR2_X1    g732(.A1(new_n665_), .A2(G162gat), .ZN(new_n934_));
  OAI21_X1  g733(.A(new_n933_), .B1(new_n925_), .B2(new_n934_), .ZN(G1347gat));
  XOR2_X1   g734(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n936_));
  NOR3_X1   g735(.A1(new_n425_), .A2(new_n385_), .A3(new_n332_), .ZN(new_n937_));
  OAI211_X1 g736(.A(new_n655_), .B(new_n937_), .C1(new_n897_), .C2(new_n873_), .ZN(new_n938_));
  NOR2_X1   g737(.A1(new_n938_), .A2(new_n523_), .ZN(new_n939_));
  INV_X1    g738(.A(KEYINPUT22), .ZN(new_n940_));
  AOI21_X1  g739(.A(new_n936_), .B1(new_n939_), .B2(new_n940_), .ZN(new_n941_));
  NAND2_X1  g740(.A1(new_n941_), .A2(G169gat), .ZN(new_n942_));
  AOI21_X1  g741(.A(new_n225_), .B1(new_n939_), .B2(new_n936_), .ZN(new_n943_));
  OAI21_X1  g742(.A(new_n942_), .B1(new_n941_), .B2(new_n943_), .ZN(G1348gat));
  NOR2_X1   g743(.A1(new_n879_), .A2(new_n303_), .ZN(new_n945_));
  NOR2_X1   g744(.A1(new_n908_), .A2(new_n226_), .ZN(new_n946_));
  NAND4_X1  g745(.A1(new_n945_), .A2(KEYINPUT123), .A3(new_n937_), .A4(new_n946_), .ZN(new_n947_));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n948_));
  INV_X1    g747(.A(new_n946_), .ZN(new_n949_));
  OAI21_X1  g748(.A(new_n948_), .B1(new_n938_), .B2(new_n949_), .ZN(new_n950_));
  NAND2_X1  g749(.A1(new_n947_), .A2(new_n950_), .ZN(new_n951_));
  OAI21_X1  g750(.A(new_n226_), .B1(new_n938_), .B2(new_n646_), .ZN(new_n952_));
  NAND2_X1  g751(.A1(new_n951_), .A2(new_n952_), .ZN(new_n953_));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n954_));
  NAND2_X1  g753(.A1(new_n953_), .A2(new_n954_), .ZN(new_n955_));
  NAND3_X1  g754(.A1(new_n951_), .A2(KEYINPUT124), .A3(new_n952_), .ZN(new_n956_));
  NAND2_X1  g755(.A1(new_n955_), .A2(new_n956_), .ZN(G1349gat));
  NOR2_X1   g756(.A1(new_n938_), .A2(new_n667_), .ZN(new_n958_));
  NAND2_X1  g757(.A1(new_n258_), .A2(KEYINPUT125), .ZN(new_n959_));
  NAND3_X1  g758(.A1(new_n958_), .A2(new_n236_), .A3(new_n959_), .ZN(new_n960_));
  NOR2_X1   g759(.A1(KEYINPUT125), .A2(G183gat), .ZN(new_n961_));
  OAI21_X1  g760(.A(new_n960_), .B1(new_n958_), .B2(new_n961_), .ZN(G1350gat));
  OAI21_X1  g761(.A(G190gat), .B1(new_n938_), .B2(new_n595_), .ZN(new_n963_));
  NAND2_X1  g762(.A1(new_n664_), .A2(new_n237_), .ZN(new_n964_));
  OAI21_X1  g763(.A(new_n963_), .B1(new_n938_), .B2(new_n964_), .ZN(G1351gat));
  NAND3_X1  g764(.A1(new_n945_), .A2(new_n661_), .A3(new_n332_), .ZN(new_n966_));
  NOR2_X1   g765(.A1(new_n966_), .A2(new_n523_), .ZN(new_n967_));
  XNOR2_X1  g766(.A(KEYINPUT126), .B(G197gat), .ZN(new_n968_));
  XNOR2_X1  g767(.A(new_n967_), .B(new_n968_), .ZN(G1352gat));
  NOR2_X1   g768(.A1(new_n966_), .A2(new_n908_), .ZN(new_n970_));
  NAND2_X1  g769(.A1(KEYINPUT127), .A2(G204gat), .ZN(new_n971_));
  XNOR2_X1  g770(.A(new_n970_), .B(new_n971_), .ZN(G1353gat));
  NOR2_X1   g771(.A1(new_n966_), .A2(new_n667_), .ZN(new_n973_));
  NOR3_X1   g772(.A1(new_n973_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n974_));
  XNOR2_X1  g773(.A(KEYINPUT63), .B(G211gat), .ZN(new_n975_));
  NOR3_X1   g774(.A1(new_n966_), .A2(new_n667_), .A3(new_n975_), .ZN(new_n976_));
  NOR2_X1   g775(.A1(new_n974_), .A2(new_n976_), .ZN(G1354gat));
  OAI21_X1  g776(.A(G218gat), .B1(new_n966_), .B2(new_n595_), .ZN(new_n978_));
  OR2_X1    g777(.A1(new_n665_), .A2(G218gat), .ZN(new_n979_));
  OAI21_X1  g778(.A(new_n978_), .B1(new_n966_), .B2(new_n979_), .ZN(G1355gat));
endmodule


