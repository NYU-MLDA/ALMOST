//Secret key is'1 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Mar 25 21:34:04 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n639_, new_n640_, new_n641_, new_n642_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n730_, new_n731_,
    new_n732_, new_n733_, new_n734_, new_n735_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n825_,
    new_n826_, new_n827_, new_n829_, new_n830_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n839_, new_n841_,
    new_n842_, new_n843_, new_n844_, new_n845_, new_n846_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n884_, new_n885_, new_n886_,
    new_n888_, new_n889_, new_n891_, new_n892_, new_n893_, new_n894_,
    new_n896_, new_n897_, new_n898_, new_n899_, new_n900_, new_n901_,
    new_n902_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n919_, new_n920_, new_n921_;
  INV_X1    g000(.A(KEYINPUT68), .ZN(new_n202_));
  XOR2_X1   g001(.A(KEYINPUT10), .B(G99gat), .Z(new_n203_));
  INV_X1    g002(.A(G106gat), .ZN(new_n204_));
  NAND2_X1  g003(.A1(new_n203_), .A2(new_n204_), .ZN(new_n205_));
  XOR2_X1   g004(.A(G85gat), .B(G92gat), .Z(new_n206_));
  NAND2_X1  g005(.A1(new_n206_), .A2(KEYINPUT9), .ZN(new_n207_));
  INV_X1    g006(.A(G85gat), .ZN(new_n208_));
  INV_X1    g007(.A(G92gat), .ZN(new_n209_));
  OR3_X1    g008(.A1(new_n208_), .A2(new_n209_), .A3(KEYINPUT9), .ZN(new_n210_));
  NAND2_X1  g009(.A1(G99gat), .A2(G106gat), .ZN(new_n211_));
  NAND2_X1  g010(.A1(new_n211_), .A2(KEYINPUT6), .ZN(new_n212_));
  INV_X1    g011(.A(KEYINPUT6), .ZN(new_n213_));
  NAND3_X1  g012(.A1(new_n213_), .A2(G99gat), .A3(G106gat), .ZN(new_n214_));
  NAND2_X1  g013(.A1(new_n212_), .A2(new_n214_), .ZN(new_n215_));
  NAND4_X1  g014(.A1(new_n205_), .A2(new_n207_), .A3(new_n210_), .A4(new_n215_), .ZN(new_n216_));
  INV_X1    g015(.A(G99gat), .ZN(new_n217_));
  NAND3_X1  g016(.A1(new_n217_), .A2(new_n204_), .A3(KEYINPUT64), .ZN(new_n218_));
  NAND2_X1  g017(.A1(new_n218_), .A2(KEYINPUT7), .ZN(new_n219_));
  INV_X1    g018(.A(KEYINPUT7), .ZN(new_n220_));
  NAND4_X1  g019(.A1(new_n220_), .A2(new_n217_), .A3(new_n204_), .A4(KEYINPUT64), .ZN(new_n221_));
  NAND3_X1  g020(.A1(new_n219_), .A2(new_n215_), .A3(new_n221_), .ZN(new_n222_));
  INV_X1    g021(.A(KEYINPUT8), .ZN(new_n223_));
  AND3_X1   g022(.A1(new_n222_), .A2(new_n223_), .A3(new_n206_), .ZN(new_n224_));
  AOI21_X1  g023(.A(new_n223_), .B1(new_n222_), .B2(new_n206_), .ZN(new_n225_));
  OAI21_X1  g024(.A(new_n216_), .B1(new_n224_), .B2(new_n225_), .ZN(new_n226_));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n227_));
  NAND2_X1  g026(.A1(new_n226_), .A2(new_n227_), .ZN(new_n228_));
  OAI211_X1 g027(.A(KEYINPUT65), .B(new_n216_), .C1(new_n224_), .C2(new_n225_), .ZN(new_n229_));
  XNOR2_X1  g028(.A(G57gat), .B(G64gat), .ZN(new_n230_));
  NAND2_X1  g029(.A1(new_n230_), .A2(KEYINPUT11), .ZN(new_n231_));
  XOR2_X1   g030(.A(G71gat), .B(G78gat), .Z(new_n232_));
  NOR2_X1   g031(.A1(new_n231_), .A2(new_n232_), .ZN(new_n233_));
  AND2_X1   g032(.A1(new_n231_), .A2(new_n232_), .ZN(new_n234_));
  OR2_X1    g033(.A1(new_n230_), .A2(KEYINPUT11), .ZN(new_n235_));
  AOI21_X1  g034(.A(new_n233_), .B1(new_n234_), .B2(new_n235_), .ZN(new_n236_));
  INV_X1    g035(.A(new_n236_), .ZN(new_n237_));
  NAND3_X1  g036(.A1(new_n228_), .A2(new_n229_), .A3(new_n237_), .ZN(new_n238_));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n239_));
  NAND2_X1  g038(.A1(new_n238_), .A2(new_n239_), .ZN(new_n240_));
  INV_X1    g039(.A(new_n225_), .ZN(new_n241_));
  NAND3_X1  g040(.A1(new_n222_), .A2(new_n223_), .A3(new_n206_), .ZN(new_n242_));
  NAND2_X1  g041(.A1(new_n241_), .A2(new_n242_), .ZN(new_n243_));
  AOI21_X1  g042(.A(KEYINPUT65), .B1(new_n243_), .B2(new_n216_), .ZN(new_n244_));
  INV_X1    g043(.A(new_n229_), .ZN(new_n245_));
  OAI21_X1  g044(.A(new_n236_), .B1(new_n244_), .B2(new_n245_), .ZN(new_n246_));
  NAND4_X1  g045(.A1(new_n228_), .A2(KEYINPUT66), .A3(new_n229_), .A4(new_n237_), .ZN(new_n247_));
  NAND3_X1  g046(.A1(new_n240_), .A2(new_n246_), .A3(new_n247_), .ZN(new_n248_));
  NAND2_X1  g047(.A1(G230gat), .A2(G233gat), .ZN(new_n249_));
  INV_X1    g048(.A(new_n249_), .ZN(new_n250_));
  NAND2_X1  g049(.A1(new_n248_), .A2(new_n250_), .ZN(new_n251_));
  INV_X1    g050(.A(KEYINPUT12), .ZN(new_n252_));
  NAND2_X1  g051(.A1(new_n246_), .A2(new_n252_), .ZN(new_n253_));
  NAND3_X1  g052(.A1(new_n226_), .A2(KEYINPUT12), .A3(new_n236_), .ZN(new_n254_));
  AND2_X1   g053(.A1(new_n238_), .A2(new_n254_), .ZN(new_n255_));
  NAND3_X1  g054(.A1(new_n253_), .A2(new_n255_), .A3(new_n249_), .ZN(new_n256_));
  XOR2_X1   g055(.A(G120gat), .B(G148gat), .Z(new_n257_));
  XNOR2_X1  g056(.A(KEYINPUT67), .B(KEYINPUT5), .ZN(new_n258_));
  XNOR2_X1  g057(.A(new_n257_), .B(new_n258_), .ZN(new_n259_));
  XNOR2_X1  g058(.A(G176gat), .B(G204gat), .ZN(new_n260_));
  XNOR2_X1  g059(.A(new_n259_), .B(new_n260_), .ZN(new_n261_));
  NAND3_X1  g060(.A1(new_n251_), .A2(new_n256_), .A3(new_n261_), .ZN(new_n262_));
  INV_X1    g061(.A(new_n262_), .ZN(new_n263_));
  AOI21_X1  g062(.A(new_n261_), .B1(new_n251_), .B2(new_n256_), .ZN(new_n264_));
  OAI21_X1  g063(.A(new_n202_), .B1(new_n263_), .B2(new_n264_), .ZN(new_n265_));
  NAND2_X1  g064(.A1(new_n251_), .A2(new_n256_), .ZN(new_n266_));
  INV_X1    g065(.A(new_n261_), .ZN(new_n267_));
  NAND2_X1  g066(.A1(new_n266_), .A2(new_n267_), .ZN(new_n268_));
  NAND3_X1  g067(.A1(new_n268_), .A2(KEYINPUT68), .A3(new_n262_), .ZN(new_n269_));
  INV_X1    g068(.A(KEYINPUT13), .ZN(new_n270_));
  AND3_X1   g069(.A1(new_n265_), .A2(new_n269_), .A3(new_n270_), .ZN(new_n271_));
  AOI21_X1  g070(.A(new_n270_), .B1(new_n265_), .B2(new_n269_), .ZN(new_n272_));
  NOR2_X1   g071(.A1(new_n271_), .A2(new_n272_), .ZN(new_n273_));
  XOR2_X1   g072(.A(G127gat), .B(G155gat), .Z(new_n274_));
  XNOR2_X1  g073(.A(new_n274_), .B(KEYINPUT16), .ZN(new_n275_));
  XNOR2_X1  g074(.A(G183gat), .B(G211gat), .ZN(new_n276_));
  XNOR2_X1  g075(.A(new_n275_), .B(new_n276_), .ZN(new_n277_));
  XNOR2_X1  g076(.A(G15gat), .B(G22gat), .ZN(new_n278_));
  INV_X1    g077(.A(G1gat), .ZN(new_n279_));
  INV_X1    g078(.A(G8gat), .ZN(new_n280_));
  OAI21_X1  g079(.A(KEYINPUT14), .B1(new_n279_), .B2(new_n280_), .ZN(new_n281_));
  NAND2_X1  g080(.A1(new_n278_), .A2(new_n281_), .ZN(new_n282_));
  XNOR2_X1  g081(.A(G1gat), .B(G8gat), .ZN(new_n283_));
  XOR2_X1   g082(.A(new_n282_), .B(new_n283_), .Z(new_n284_));
  NAND2_X1  g083(.A1(G231gat), .A2(G233gat), .ZN(new_n285_));
  XOR2_X1   g084(.A(new_n284_), .B(new_n285_), .Z(new_n286_));
  XNOR2_X1  g085(.A(new_n286_), .B(new_n237_), .ZN(new_n287_));
  INV_X1    g086(.A(new_n287_), .ZN(new_n288_));
  OAI21_X1  g087(.A(new_n277_), .B1(new_n288_), .B2(KEYINPUT17), .ZN(new_n289_));
  OAI21_X1  g088(.A(new_n289_), .B1(KEYINPUT17), .B2(new_n277_), .ZN(new_n290_));
  NAND2_X1  g089(.A1(new_n287_), .A2(KEYINPUT74), .ZN(new_n291_));
  XNOR2_X1  g090(.A(new_n290_), .B(new_n291_), .ZN(new_n292_));
  XNOR2_X1  g091(.A(G29gat), .B(G36gat), .ZN(new_n293_));
  XNOR2_X1  g092(.A(G43gat), .B(G50gat), .ZN(new_n294_));
  XNOR2_X1  g093(.A(new_n293_), .B(new_n294_), .ZN(new_n295_));
  NAND2_X1  g094(.A1(new_n284_), .A2(new_n295_), .ZN(new_n296_));
  NAND2_X1  g095(.A1(new_n296_), .A2(KEYINPUT75), .ZN(new_n297_));
  OR2_X1    g096(.A1(new_n284_), .A2(new_n295_), .ZN(new_n298_));
  XNOR2_X1  g097(.A(new_n297_), .B(new_n298_), .ZN(new_n299_));
  NAND2_X1  g098(.A1(G229gat), .A2(G233gat), .ZN(new_n300_));
  INV_X1    g099(.A(new_n300_), .ZN(new_n301_));
  NAND2_X1  g100(.A1(new_n299_), .A2(new_n301_), .ZN(new_n302_));
  INV_X1    g101(.A(new_n296_), .ZN(new_n303_));
  XNOR2_X1  g102(.A(new_n295_), .B(KEYINPUT15), .ZN(new_n304_));
  INV_X1    g103(.A(new_n284_), .ZN(new_n305_));
  AOI21_X1  g104(.A(new_n303_), .B1(new_n304_), .B2(new_n305_), .ZN(new_n306_));
  NAND2_X1  g105(.A1(new_n306_), .A2(new_n300_), .ZN(new_n307_));
  NAND2_X1  g106(.A1(new_n302_), .A2(new_n307_), .ZN(new_n308_));
  XNOR2_X1  g107(.A(G113gat), .B(G141gat), .ZN(new_n309_));
  XNOR2_X1  g108(.A(new_n309_), .B(KEYINPUT76), .ZN(new_n310_));
  XNOR2_X1  g109(.A(G169gat), .B(G197gat), .ZN(new_n311_));
  XOR2_X1   g110(.A(new_n310_), .B(new_n311_), .Z(new_n312_));
  XNOR2_X1  g111(.A(new_n308_), .B(new_n312_), .ZN(new_n313_));
  NAND3_X1  g112(.A1(new_n273_), .A2(new_n292_), .A3(new_n313_), .ZN(new_n314_));
  XNOR2_X1  g113(.A(new_n314_), .B(KEYINPUT96), .ZN(new_n315_));
  NAND3_X1  g114(.A1(new_n228_), .A2(new_n295_), .A3(new_n229_), .ZN(new_n316_));
  NAND2_X1  g115(.A1(new_n316_), .A2(KEYINPUT71), .ZN(new_n317_));
  NAND2_X1  g116(.A1(new_n304_), .A2(new_n226_), .ZN(new_n318_));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n319_));
  NAND4_X1  g118(.A1(new_n228_), .A2(new_n319_), .A3(new_n295_), .A4(new_n229_), .ZN(new_n320_));
  NAND2_X1  g119(.A1(G232gat), .A2(G233gat), .ZN(new_n321_));
  XNOR2_X1  g120(.A(new_n321_), .B(KEYINPUT34), .ZN(new_n322_));
  OR2_X1    g121(.A1(new_n322_), .A2(KEYINPUT35), .ZN(new_n323_));
  NAND4_X1  g122(.A1(new_n317_), .A2(new_n318_), .A3(new_n320_), .A4(new_n323_), .ZN(new_n324_));
  NAND4_X1  g123(.A1(new_n317_), .A2(KEYINPUT70), .A3(new_n320_), .A4(new_n323_), .ZN(new_n325_));
  NAND2_X1  g124(.A1(new_n322_), .A2(KEYINPUT35), .ZN(new_n326_));
  XNOR2_X1  g125(.A(new_n326_), .B(KEYINPUT69), .ZN(new_n327_));
  INV_X1    g126(.A(new_n327_), .ZN(new_n328_));
  AND3_X1   g127(.A1(new_n324_), .A2(new_n325_), .A3(new_n328_), .ZN(new_n329_));
  AOI21_X1  g128(.A(new_n324_), .B1(new_n325_), .B2(new_n328_), .ZN(new_n330_));
  NOR2_X1   g129(.A1(new_n329_), .A2(new_n330_), .ZN(new_n331_));
  XNOR2_X1  g130(.A(G190gat), .B(G218gat), .ZN(new_n332_));
  XNOR2_X1  g131(.A(G134gat), .B(G162gat), .ZN(new_n333_));
  XNOR2_X1  g132(.A(new_n332_), .B(new_n333_), .ZN(new_n334_));
  NOR2_X1   g133(.A1(new_n334_), .A2(KEYINPUT36), .ZN(new_n335_));
  NAND3_X1  g134(.A1(new_n331_), .A2(KEYINPUT72), .A3(new_n335_), .ZN(new_n336_));
  AND3_X1   g135(.A1(new_n317_), .A2(new_n320_), .A3(new_n323_), .ZN(new_n337_));
  OAI211_X1 g136(.A(new_n337_), .B(new_n318_), .C1(KEYINPUT70), .C2(new_n327_), .ZN(new_n338_));
  NAND3_X1  g137(.A1(new_n324_), .A2(new_n325_), .A3(new_n328_), .ZN(new_n339_));
  NAND3_X1  g138(.A1(new_n338_), .A2(new_n335_), .A3(new_n339_), .ZN(new_n340_));
  INV_X1    g139(.A(KEYINPUT72), .ZN(new_n341_));
  NAND2_X1  g140(.A1(new_n340_), .A2(new_n341_), .ZN(new_n342_));
  NAND2_X1  g141(.A1(new_n336_), .A2(new_n342_), .ZN(new_n343_));
  XOR2_X1   g142(.A(new_n334_), .B(KEYINPUT36), .Z(new_n344_));
  OAI21_X1  g143(.A(new_n344_), .B1(new_n329_), .B2(new_n330_), .ZN(new_n345_));
  NAND2_X1  g144(.A1(new_n343_), .A2(new_n345_), .ZN(new_n346_));
  INV_X1    g145(.A(KEYINPUT95), .ZN(new_n347_));
  INV_X1    g146(.A(G197gat), .ZN(new_n348_));
  INV_X1    g147(.A(G204gat), .ZN(new_n349_));
  NAND2_X1  g148(.A1(new_n348_), .A2(new_n349_), .ZN(new_n350_));
  NAND2_X1  g149(.A1(G197gat), .A2(G204gat), .ZN(new_n351_));
  AND3_X1   g150(.A1(new_n350_), .A2(KEYINPUT21), .A3(new_n351_), .ZN(new_n352_));
  XNOR2_X1  g151(.A(G211gat), .B(G218gat), .ZN(new_n353_));
  OR2_X1    g152(.A1(new_n352_), .A2(new_n353_), .ZN(new_n354_));
  AOI21_X1  g153(.A(KEYINPUT21), .B1(new_n350_), .B2(new_n351_), .ZN(new_n355_));
  OAI21_X1  g154(.A(new_n353_), .B1(new_n352_), .B2(new_n355_), .ZN(new_n356_));
  NAND2_X1  g155(.A1(new_n354_), .A2(new_n356_), .ZN(new_n357_));
  INV_X1    g156(.A(G183gat), .ZN(new_n358_));
  INV_X1    g157(.A(G190gat), .ZN(new_n359_));
  NOR3_X1   g158(.A1(new_n358_), .A2(new_n359_), .A3(KEYINPUT23), .ZN(new_n360_));
  INV_X1    g159(.A(new_n360_), .ZN(new_n361_));
  OAI21_X1  g160(.A(KEYINPUT23), .B1(new_n358_), .B2(new_n359_), .ZN(new_n362_));
  NAND2_X1  g161(.A1(new_n361_), .A2(new_n362_), .ZN(new_n363_));
  OR2_X1    g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364_));
  NAND2_X1  g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365_));
  NAND3_X1  g164(.A1(new_n364_), .A2(KEYINPUT24), .A3(new_n365_), .ZN(new_n366_));
  OR2_X1    g165(.A1(new_n364_), .A2(KEYINPUT24), .ZN(new_n367_));
  XNOR2_X1  g166(.A(KEYINPUT25), .B(G183gat), .ZN(new_n368_));
  XNOR2_X1  g167(.A(KEYINPUT26), .B(G190gat), .ZN(new_n369_));
  NAND2_X1  g168(.A1(new_n368_), .A2(new_n369_), .ZN(new_n370_));
  NAND4_X1  g169(.A1(new_n363_), .A2(new_n366_), .A3(new_n367_), .A4(new_n370_), .ZN(new_n371_));
  AND2_X1   g170(.A1(new_n357_), .A2(new_n371_), .ZN(new_n372_));
  INV_X1    g171(.A(KEYINPUT90), .ZN(new_n373_));
  XNOR2_X1  g172(.A(KEYINPUT22), .B(G169gat), .ZN(new_n374_));
  INV_X1    g173(.A(G176gat), .ZN(new_n375_));
  NAND2_X1  g174(.A1(new_n374_), .A2(new_n375_), .ZN(new_n376_));
  NAND2_X1  g175(.A1(new_n376_), .A2(new_n365_), .ZN(new_n377_));
  INV_X1    g176(.A(KEYINPUT23), .ZN(new_n378_));
  AOI21_X1  g177(.A(new_n378_), .B1(G183gat), .B2(G190gat), .ZN(new_n379_));
  INV_X1    g178(.A(KEYINPUT79), .ZN(new_n380_));
  NOR2_X1   g179(.A1(new_n379_), .A2(new_n380_), .ZN(new_n381_));
  NOR2_X1   g180(.A1(new_n362_), .A2(KEYINPUT79), .ZN(new_n382_));
  OAI21_X1  g181(.A(new_n361_), .B1(new_n381_), .B2(new_n382_), .ZN(new_n383_));
  NOR2_X1   g182(.A1(G183gat), .A2(G190gat), .ZN(new_n384_));
  INV_X1    g183(.A(new_n384_), .ZN(new_n385_));
  NAND2_X1  g184(.A1(new_n383_), .A2(new_n385_), .ZN(new_n386_));
  INV_X1    g185(.A(KEYINPUT89), .ZN(new_n387_));
  AOI21_X1  g186(.A(new_n377_), .B1(new_n386_), .B2(new_n387_), .ZN(new_n388_));
  NAND3_X1  g187(.A1(new_n383_), .A2(KEYINPUT89), .A3(new_n385_), .ZN(new_n389_));
  AOI21_X1  g188(.A(new_n373_), .B1(new_n388_), .B2(new_n389_), .ZN(new_n390_));
  NAND2_X1  g189(.A1(new_n379_), .A2(new_n380_), .ZN(new_n391_));
  NAND2_X1  g190(.A1(new_n362_), .A2(KEYINPUT79), .ZN(new_n392_));
  AOI21_X1  g191(.A(new_n360_), .B1(new_n391_), .B2(new_n392_), .ZN(new_n393_));
  OAI21_X1  g192(.A(new_n387_), .B1(new_n393_), .B2(new_n384_), .ZN(new_n394_));
  INV_X1    g193(.A(new_n377_), .ZN(new_n395_));
  AND4_X1   g194(.A1(new_n373_), .A2(new_n389_), .A3(new_n394_), .A4(new_n395_), .ZN(new_n396_));
  OAI21_X1  g195(.A(new_n372_), .B1(new_n390_), .B2(new_n396_), .ZN(new_n397_));
  NAND2_X1  g196(.A1(G226gat), .A2(G233gat), .ZN(new_n398_));
  XNOR2_X1  g197(.A(new_n398_), .B(KEYINPUT19), .ZN(new_n399_));
  INV_X1    g198(.A(new_n399_), .ZN(new_n400_));
  NOR2_X1   g199(.A1(KEYINPUT26), .A2(G190gat), .ZN(new_n401_));
  XNOR2_X1  g200(.A(KEYINPUT77), .B(G190gat), .ZN(new_n402_));
  AOI21_X1  g201(.A(new_n401_), .B1(new_n402_), .B2(KEYINPUT26), .ZN(new_n403_));
  INV_X1    g202(.A(new_n368_), .ZN(new_n404_));
  OAI21_X1  g203(.A(new_n366_), .B1(new_n403_), .B2(new_n404_), .ZN(new_n405_));
  INV_X1    g204(.A(KEYINPUT78), .ZN(new_n406_));
  NAND2_X1  g205(.A1(new_n405_), .A2(new_n406_), .ZN(new_n407_));
  OAI211_X1 g206(.A(KEYINPUT78), .B(new_n366_), .C1(new_n403_), .C2(new_n404_), .ZN(new_n408_));
  NAND4_X1  g207(.A1(new_n407_), .A2(new_n408_), .A3(new_n367_), .A4(new_n383_), .ZN(new_n409_));
  INV_X1    g208(.A(new_n376_), .ZN(new_n410_));
  OR2_X1    g209(.A1(new_n410_), .A2(KEYINPUT80), .ZN(new_n411_));
  OAI21_X1  g210(.A(new_n363_), .B1(G183gat), .B2(new_n402_), .ZN(new_n412_));
  NAND2_X1  g211(.A1(new_n410_), .A2(KEYINPUT80), .ZN(new_n413_));
  NAND4_X1  g212(.A1(new_n411_), .A2(new_n365_), .A3(new_n412_), .A4(new_n413_), .ZN(new_n414_));
  NAND2_X1  g213(.A1(new_n409_), .A2(new_n414_), .ZN(new_n415_));
  INV_X1    g214(.A(new_n357_), .ZN(new_n416_));
  NAND2_X1  g215(.A1(new_n415_), .A2(new_n416_), .ZN(new_n417_));
  NAND4_X1  g216(.A1(new_n397_), .A2(KEYINPUT20), .A3(new_n400_), .A4(new_n417_), .ZN(new_n418_));
  NAND3_X1  g217(.A1(new_n409_), .A2(new_n414_), .A3(new_n357_), .ZN(new_n419_));
  NAND2_X1  g218(.A1(new_n419_), .A2(KEYINPUT20), .ZN(new_n420_));
  OAI21_X1  g219(.A(new_n371_), .B1(new_n390_), .B2(new_n396_), .ZN(new_n421_));
  AOI21_X1  g220(.A(new_n420_), .B1(new_n421_), .B2(new_n416_), .ZN(new_n422_));
  OAI21_X1  g221(.A(new_n418_), .B1(new_n422_), .B2(new_n400_), .ZN(new_n423_));
  XNOR2_X1  g222(.A(G8gat), .B(G36gat), .ZN(new_n424_));
  XNOR2_X1  g223(.A(new_n424_), .B(KEYINPUT18), .ZN(new_n425_));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426_));
  XOR2_X1   g225(.A(new_n425_), .B(new_n426_), .Z(new_n427_));
  INV_X1    g226(.A(new_n427_), .ZN(new_n428_));
  NAND2_X1  g227(.A1(new_n423_), .A2(new_n428_), .ZN(new_n429_));
  OAI211_X1 g228(.A(new_n427_), .B(new_n418_), .C1(new_n422_), .C2(new_n400_), .ZN(new_n430_));
  AOI21_X1  g229(.A(KEYINPUT27), .B1(new_n429_), .B2(new_n430_), .ZN(new_n431_));
  NAND2_X1  g230(.A1(new_n430_), .A2(KEYINPUT27), .ZN(new_n432_));
  NAND2_X1  g231(.A1(new_n422_), .A2(new_n400_), .ZN(new_n433_));
  NAND2_X1  g232(.A1(new_n388_), .A2(new_n389_), .ZN(new_n434_));
  NAND2_X1  g233(.A1(new_n434_), .A2(new_n372_), .ZN(new_n435_));
  NAND3_X1  g234(.A1(new_n417_), .A2(KEYINPUT20), .A3(new_n435_), .ZN(new_n436_));
  NAND2_X1  g235(.A1(new_n436_), .A2(new_n399_), .ZN(new_n437_));
  AOI21_X1  g236(.A(new_n427_), .B1(new_n433_), .B2(new_n437_), .ZN(new_n438_));
  NOR2_X1   g237(.A1(new_n432_), .A2(new_n438_), .ZN(new_n439_));
  INV_X1    g238(.A(KEYINPUT3), .ZN(new_n440_));
  INV_X1    g239(.A(G141gat), .ZN(new_n441_));
  INV_X1    g240(.A(G148gat), .ZN(new_n442_));
  NAND4_X1  g241(.A1(new_n440_), .A2(new_n441_), .A3(new_n442_), .A4(KEYINPUT87), .ZN(new_n443_));
  INV_X1    g242(.A(KEYINPUT87), .ZN(new_n444_));
  OAI22_X1  g243(.A1(new_n444_), .A2(KEYINPUT3), .B1(G141gat), .B2(G148gat), .ZN(new_n445_));
  NAND2_X1  g244(.A1(G141gat), .A2(G148gat), .ZN(new_n446_));
  INV_X1    g245(.A(KEYINPUT2), .ZN(new_n447_));
  NAND2_X1  g246(.A1(new_n446_), .A2(new_n447_), .ZN(new_n448_));
  NAND3_X1  g247(.A1(KEYINPUT2), .A2(G141gat), .A3(G148gat), .ZN(new_n449_));
  NAND4_X1  g248(.A1(new_n443_), .A2(new_n445_), .A3(new_n448_), .A4(new_n449_), .ZN(new_n450_));
  OR3_X1    g249(.A1(KEYINPUT86), .A2(G155gat), .A3(G162gat), .ZN(new_n451_));
  OAI21_X1  g250(.A(KEYINPUT86), .B1(G155gat), .B2(G162gat), .ZN(new_n452_));
  NAND2_X1  g251(.A1(G155gat), .A2(G162gat), .ZN(new_n453_));
  NAND4_X1  g252(.A1(new_n450_), .A2(new_n451_), .A3(new_n452_), .A4(new_n453_), .ZN(new_n454_));
  NAND2_X1  g253(.A1(new_n453_), .A2(KEYINPUT1), .ZN(new_n455_));
  INV_X1    g254(.A(KEYINPUT1), .ZN(new_n456_));
  NAND3_X1  g255(.A1(new_n456_), .A2(G155gat), .A3(G162gat), .ZN(new_n457_));
  NAND4_X1  g256(.A1(new_n451_), .A2(new_n452_), .A3(new_n455_), .A4(new_n457_), .ZN(new_n458_));
  NAND2_X1  g257(.A1(new_n441_), .A2(new_n442_), .ZN(new_n459_));
  NAND3_X1  g258(.A1(new_n458_), .A2(new_n459_), .A3(new_n446_), .ZN(new_n460_));
  NAND2_X1  g259(.A1(new_n454_), .A2(new_n460_), .ZN(new_n461_));
  NOR2_X1   g260(.A1(new_n461_), .A2(KEYINPUT29), .ZN(new_n462_));
  XOR2_X1   g261(.A(new_n462_), .B(KEYINPUT28), .Z(new_n463_));
  AND2_X1   g262(.A1(G228gat), .A2(G233gat), .ZN(new_n464_));
  NOR2_X1   g263(.A1(new_n464_), .A2(KEYINPUT88), .ZN(new_n465_));
  XNOR2_X1  g264(.A(new_n463_), .B(new_n465_), .ZN(new_n466_));
  INV_X1    g265(.A(G78gat), .ZN(new_n467_));
  AND2_X1   g266(.A1(new_n464_), .A2(KEYINPUT88), .ZN(new_n468_));
  NOR2_X1   g267(.A1(new_n357_), .A2(new_n468_), .ZN(new_n469_));
  NAND2_X1  g268(.A1(new_n461_), .A2(KEYINPUT29), .ZN(new_n470_));
  AOI21_X1  g269(.A(new_n467_), .B1(new_n469_), .B2(new_n470_), .ZN(new_n471_));
  INV_X1    g270(.A(new_n471_), .ZN(new_n472_));
  NAND3_X1  g271(.A1(new_n469_), .A2(new_n470_), .A3(new_n467_), .ZN(new_n473_));
  NAND3_X1  g272(.A1(new_n472_), .A2(G106gat), .A3(new_n473_), .ZN(new_n474_));
  INV_X1    g273(.A(new_n473_), .ZN(new_n475_));
  OAI21_X1  g274(.A(new_n204_), .B1(new_n475_), .B2(new_n471_), .ZN(new_n476_));
  XNOR2_X1  g275(.A(G22gat), .B(G50gat), .ZN(new_n477_));
  INV_X1    g276(.A(new_n477_), .ZN(new_n478_));
  NAND3_X1  g277(.A1(new_n474_), .A2(new_n476_), .A3(new_n478_), .ZN(new_n479_));
  INV_X1    g278(.A(new_n479_), .ZN(new_n480_));
  AOI21_X1  g279(.A(new_n478_), .B1(new_n474_), .B2(new_n476_), .ZN(new_n481_));
  OAI21_X1  g280(.A(new_n466_), .B1(new_n480_), .B2(new_n481_), .ZN(new_n482_));
  NAND2_X1  g281(.A1(G225gat), .A2(G233gat), .ZN(new_n483_));
  XNOR2_X1  g282(.A(G113gat), .B(G120gat), .ZN(new_n484_));
  INV_X1    g283(.A(new_n484_), .ZN(new_n485_));
  XNOR2_X1  g284(.A(G127gat), .B(G134gat), .ZN(new_n486_));
  NOR2_X1   g285(.A1(new_n486_), .A2(KEYINPUT84), .ZN(new_n487_));
  INV_X1    g286(.A(G134gat), .ZN(new_n488_));
  NAND2_X1  g287(.A1(new_n488_), .A2(G127gat), .ZN(new_n489_));
  INV_X1    g288(.A(G127gat), .ZN(new_n490_));
  NAND2_X1  g289(.A1(new_n490_), .A2(G134gat), .ZN(new_n491_));
  AND3_X1   g290(.A1(new_n489_), .A2(new_n491_), .A3(KEYINPUT84), .ZN(new_n492_));
  OAI21_X1  g291(.A(new_n485_), .B1(new_n487_), .B2(new_n492_), .ZN(new_n493_));
  NAND2_X1  g292(.A1(new_n489_), .A2(new_n491_), .ZN(new_n494_));
  INV_X1    g293(.A(KEYINPUT84), .ZN(new_n495_));
  NAND2_X1  g294(.A1(new_n494_), .A2(new_n495_), .ZN(new_n496_));
  NAND2_X1  g295(.A1(new_n486_), .A2(KEYINPUT84), .ZN(new_n497_));
  NAND3_X1  g296(.A1(new_n496_), .A2(new_n497_), .A3(new_n484_), .ZN(new_n498_));
  NAND2_X1  g297(.A1(new_n493_), .A2(new_n498_), .ZN(new_n499_));
  NAND2_X1  g298(.A1(new_n461_), .A2(new_n499_), .ZN(new_n500_));
  NAND4_X1  g299(.A1(new_n454_), .A2(new_n493_), .A3(new_n460_), .A4(new_n498_), .ZN(new_n501_));
  NAND3_X1  g300(.A1(new_n500_), .A2(KEYINPUT4), .A3(new_n501_), .ZN(new_n502_));
  INV_X1    g301(.A(KEYINPUT4), .ZN(new_n503_));
  NAND3_X1  g302(.A1(new_n461_), .A2(new_n499_), .A3(new_n503_), .ZN(new_n504_));
  AOI21_X1  g303(.A(new_n483_), .B1(new_n502_), .B2(new_n504_), .ZN(new_n505_));
  XNOR2_X1  g304(.A(G1gat), .B(G29gat), .ZN(new_n506_));
  XNOR2_X1  g305(.A(KEYINPUT91), .B(KEYINPUT0), .ZN(new_n507_));
  XNOR2_X1  g306(.A(new_n506_), .B(new_n507_), .ZN(new_n508_));
  XNOR2_X1  g307(.A(G57gat), .B(G85gat), .ZN(new_n509_));
  XNOR2_X1  g308(.A(new_n508_), .B(new_n509_), .ZN(new_n510_));
  INV_X1    g309(.A(new_n510_), .ZN(new_n511_));
  INV_X1    g310(.A(new_n483_), .ZN(new_n512_));
  AOI21_X1  g311(.A(new_n512_), .B1(new_n500_), .B2(new_n501_), .ZN(new_n513_));
  OR3_X1    g312(.A1(new_n505_), .A2(new_n511_), .A3(new_n513_), .ZN(new_n514_));
  INV_X1    g313(.A(KEYINPUT94), .ZN(new_n515_));
  OAI21_X1  g314(.A(new_n511_), .B1(new_n505_), .B2(new_n513_), .ZN(new_n516_));
  NAND3_X1  g315(.A1(new_n514_), .A2(new_n515_), .A3(new_n516_), .ZN(new_n517_));
  OAI211_X1 g316(.A(KEYINPUT94), .B(new_n511_), .C1(new_n505_), .C2(new_n513_), .ZN(new_n518_));
  NAND2_X1  g317(.A1(new_n517_), .A2(new_n518_), .ZN(new_n519_));
  INV_X1    g318(.A(new_n465_), .ZN(new_n520_));
  XNOR2_X1  g319(.A(new_n463_), .B(new_n520_), .ZN(new_n521_));
  NAND2_X1  g320(.A1(new_n474_), .A2(new_n476_), .ZN(new_n522_));
  NAND2_X1  g321(.A1(new_n522_), .A2(new_n477_), .ZN(new_n523_));
  NAND3_X1  g322(.A1(new_n521_), .A2(new_n523_), .A3(new_n479_), .ZN(new_n524_));
  NAND3_X1  g323(.A1(new_n482_), .A2(new_n519_), .A3(new_n524_), .ZN(new_n525_));
  NOR3_X1   g324(.A1(new_n431_), .A2(new_n439_), .A3(new_n525_), .ZN(new_n526_));
  INV_X1    g325(.A(KEYINPUT93), .ZN(new_n527_));
  NAND2_X1  g326(.A1(new_n429_), .A2(new_n430_), .ZN(new_n528_));
  OAI211_X1 g327(.A(KEYINPUT33), .B(new_n511_), .C1(new_n505_), .C2(new_n513_), .ZN(new_n529_));
  NAND3_X1  g328(.A1(new_n502_), .A2(new_n483_), .A3(new_n504_), .ZN(new_n530_));
  NAND2_X1  g329(.A1(new_n500_), .A2(new_n501_), .ZN(new_n531_));
  OAI211_X1 g330(.A(new_n530_), .B(new_n510_), .C1(new_n483_), .C2(new_n531_), .ZN(new_n532_));
  INV_X1    g331(.A(KEYINPUT92), .ZN(new_n533_));
  INV_X1    g332(.A(KEYINPUT33), .ZN(new_n534_));
  NAND3_X1  g333(.A1(new_n516_), .A2(new_n533_), .A3(new_n534_), .ZN(new_n535_));
  INV_X1    g334(.A(new_n535_), .ZN(new_n536_));
  AOI21_X1  g335(.A(new_n533_), .B1(new_n516_), .B2(new_n534_), .ZN(new_n537_));
  OAI211_X1 g336(.A(new_n529_), .B(new_n532_), .C1(new_n536_), .C2(new_n537_), .ZN(new_n538_));
  OAI21_X1  g337(.A(new_n527_), .B1(new_n528_), .B2(new_n538_), .ZN(new_n539_));
  NAND2_X1  g338(.A1(new_n427_), .A2(KEYINPUT32), .ZN(new_n540_));
  AOI21_X1  g339(.A(new_n540_), .B1(new_n433_), .B2(new_n437_), .ZN(new_n541_));
  NOR2_X1   g340(.A1(new_n541_), .A2(new_n519_), .ZN(new_n542_));
  OAI211_X1 g341(.A(new_n418_), .B(new_n540_), .C1(new_n422_), .C2(new_n400_), .ZN(new_n543_));
  NAND2_X1  g342(.A1(new_n542_), .A2(new_n543_), .ZN(new_n544_));
  NAND2_X1  g343(.A1(new_n529_), .A2(new_n532_), .ZN(new_n545_));
  NAND2_X1  g344(.A1(new_n516_), .A2(new_n534_), .ZN(new_n546_));
  NAND2_X1  g345(.A1(new_n546_), .A2(KEYINPUT92), .ZN(new_n547_));
  AOI21_X1  g346(.A(new_n545_), .B1(new_n547_), .B2(new_n535_), .ZN(new_n548_));
  NAND4_X1  g347(.A1(new_n548_), .A2(KEYINPUT93), .A3(new_n430_), .A4(new_n429_), .ZN(new_n549_));
  NAND3_X1  g348(.A1(new_n539_), .A2(new_n544_), .A3(new_n549_), .ZN(new_n550_));
  NAND2_X1  g349(.A1(new_n482_), .A2(new_n524_), .ZN(new_n551_));
  AOI21_X1  g350(.A(new_n526_), .B1(new_n550_), .B2(new_n551_), .ZN(new_n552_));
  NAND3_X1  g351(.A1(new_n409_), .A2(KEYINPUT30), .A3(new_n414_), .ZN(new_n553_));
  INV_X1    g352(.A(new_n553_), .ZN(new_n554_));
  AOI21_X1  g353(.A(KEYINPUT30), .B1(new_n409_), .B2(new_n414_), .ZN(new_n555_));
  NOR2_X1   g354(.A1(new_n554_), .A2(new_n555_), .ZN(new_n556_));
  XNOR2_X1  g355(.A(G15gat), .B(G43gat), .ZN(new_n557_));
  XNOR2_X1  g356(.A(new_n557_), .B(KEYINPUT81), .ZN(new_n558_));
  XNOR2_X1  g357(.A(new_n558_), .B(G99gat), .ZN(new_n559_));
  NAND2_X1  g358(.A1(G227gat), .A2(G233gat), .ZN(new_n560_));
  XOR2_X1   g359(.A(new_n560_), .B(G71gat), .Z(new_n561_));
  XNOR2_X1  g360(.A(new_n559_), .B(new_n561_), .ZN(new_n562_));
  OAI21_X1  g361(.A(KEYINPUT82), .B1(new_n556_), .B2(new_n562_), .ZN(new_n563_));
  INV_X1    g362(.A(new_n562_), .ZN(new_n564_));
  INV_X1    g363(.A(KEYINPUT82), .ZN(new_n565_));
  OAI211_X1 g364(.A(new_n564_), .B(new_n565_), .C1(new_n555_), .C2(new_n554_), .ZN(new_n566_));
  NAND2_X1  g365(.A1(new_n563_), .A2(new_n566_), .ZN(new_n567_));
  INV_X1    g366(.A(new_n555_), .ZN(new_n568_));
  NAND3_X1  g367(.A1(new_n562_), .A2(new_n568_), .A3(new_n553_), .ZN(new_n569_));
  NAND2_X1  g368(.A1(new_n569_), .A2(KEYINPUT83), .ZN(new_n570_));
  INV_X1    g369(.A(KEYINPUT83), .ZN(new_n571_));
  NAND3_X1  g370(.A1(new_n556_), .A2(new_n571_), .A3(new_n562_), .ZN(new_n572_));
  NAND2_X1  g371(.A1(new_n570_), .A2(new_n572_), .ZN(new_n573_));
  NAND2_X1  g372(.A1(new_n567_), .A2(new_n573_), .ZN(new_n574_));
  NAND2_X1  g373(.A1(new_n574_), .A2(KEYINPUT85), .ZN(new_n575_));
  INV_X1    g374(.A(KEYINPUT85), .ZN(new_n576_));
  NAND3_X1  g375(.A1(new_n567_), .A2(new_n573_), .A3(new_n576_), .ZN(new_n577_));
  XNOR2_X1  g376(.A(new_n499_), .B(KEYINPUT31), .ZN(new_n578_));
  NAND3_X1  g377(.A1(new_n575_), .A2(new_n577_), .A3(new_n578_), .ZN(new_n579_));
  INV_X1    g378(.A(new_n578_), .ZN(new_n580_));
  NAND4_X1  g379(.A1(new_n567_), .A2(new_n573_), .A3(new_n576_), .A4(new_n580_), .ZN(new_n581_));
  NAND2_X1  g380(.A1(new_n579_), .A2(new_n581_), .ZN(new_n582_));
  INV_X1    g381(.A(new_n582_), .ZN(new_n583_));
  OAI21_X1  g382(.A(new_n347_), .B1(new_n552_), .B2(new_n583_), .ZN(new_n584_));
  INV_X1    g383(.A(new_n551_), .ZN(new_n585_));
  NAND3_X1  g384(.A1(new_n548_), .A2(new_n430_), .A3(new_n429_), .ZN(new_n586_));
  AOI22_X1  g385(.A1(new_n586_), .A2(new_n527_), .B1(new_n542_), .B2(new_n543_), .ZN(new_n587_));
  AOI21_X1  g386(.A(new_n585_), .B1(new_n587_), .B2(new_n549_), .ZN(new_n588_));
  OAI211_X1 g387(.A(KEYINPUT95), .B(new_n582_), .C1(new_n588_), .C2(new_n526_), .ZN(new_n589_));
  NOR2_X1   g388(.A1(new_n431_), .A2(new_n439_), .ZN(new_n590_));
  NAND2_X1  g389(.A1(new_n590_), .A2(new_n551_), .ZN(new_n591_));
  NAND3_X1  g390(.A1(new_n579_), .A2(new_n581_), .A3(new_n519_), .ZN(new_n592_));
  OR2_X1    g391(.A1(new_n591_), .A2(new_n592_), .ZN(new_n593_));
  NAND3_X1  g392(.A1(new_n584_), .A2(new_n589_), .A3(new_n593_), .ZN(new_n594_));
  AND3_X1   g393(.A1(new_n315_), .A2(new_n346_), .A3(new_n594_), .ZN(new_n595_));
  INV_X1    g394(.A(new_n595_), .ZN(new_n596_));
  OAI21_X1  g395(.A(G1gat), .B1(new_n596_), .B2(new_n519_), .ZN(new_n597_));
  INV_X1    g396(.A(KEYINPUT38), .ZN(new_n598_));
  INV_X1    g397(.A(new_n273_), .ZN(new_n599_));
  INV_X1    g398(.A(new_n313_), .ZN(new_n600_));
  NOR2_X1   g399(.A1(new_n599_), .A2(new_n600_), .ZN(new_n601_));
  AND2_X1   g400(.A1(new_n594_), .A2(new_n601_), .ZN(new_n602_));
  NAND2_X1  g401(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n603_));
  AOI21_X1  g402(.A(KEYINPUT72), .B1(new_n331_), .B2(new_n335_), .ZN(new_n604_));
  AND4_X1   g403(.A1(KEYINPUT72), .A2(new_n338_), .A3(new_n335_), .A4(new_n339_), .ZN(new_n605_));
  OAI211_X1 g404(.A(new_n603_), .B(new_n345_), .C1(new_n604_), .C2(new_n605_), .ZN(new_n606_));
  NOR2_X1   g405(.A1(KEYINPUT73), .A2(KEYINPUT37), .ZN(new_n607_));
  NAND2_X1  g406(.A1(new_n606_), .A2(new_n607_), .ZN(new_n608_));
  INV_X1    g407(.A(new_n607_), .ZN(new_n609_));
  NAND4_X1  g408(.A1(new_n343_), .A2(new_n603_), .A3(new_n345_), .A4(new_n609_), .ZN(new_n610_));
  NAND2_X1  g409(.A1(new_n608_), .A2(new_n610_), .ZN(new_n611_));
  INV_X1    g410(.A(new_n292_), .ZN(new_n612_));
  NOR2_X1   g411(.A1(new_n611_), .A2(new_n612_), .ZN(new_n613_));
  AND2_X1   g412(.A1(new_n602_), .A2(new_n613_), .ZN(new_n614_));
  INV_X1    g413(.A(new_n519_), .ZN(new_n615_));
  NAND3_X1  g414(.A1(new_n614_), .A2(new_n279_), .A3(new_n615_), .ZN(new_n616_));
  AND3_X1   g415(.A1(new_n616_), .A2(KEYINPUT97), .A3(new_n598_), .ZN(new_n617_));
  AOI21_X1  g416(.A(KEYINPUT97), .B1(new_n616_), .B2(new_n598_), .ZN(new_n618_));
  OAI221_X1 g417(.A(new_n597_), .B1(new_n598_), .B2(new_n616_), .C1(new_n617_), .C2(new_n618_), .ZN(G1324gat));
  XNOR2_X1  g418(.A(KEYINPUT98), .B(KEYINPUT40), .ZN(new_n620_));
  INV_X1    g419(.A(new_n590_), .ZN(new_n621_));
  AOI21_X1  g420(.A(new_n280_), .B1(new_n595_), .B2(new_n621_), .ZN(new_n622_));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n623_));
  XNOR2_X1  g422(.A(new_n622_), .B(new_n623_), .ZN(new_n624_));
  NAND3_X1  g423(.A1(new_n614_), .A2(new_n280_), .A3(new_n621_), .ZN(new_n625_));
  AOI21_X1  g424(.A(new_n620_), .B1(new_n624_), .B2(new_n625_), .ZN(new_n626_));
  NOR2_X1   g425(.A1(new_n622_), .A2(new_n623_), .ZN(new_n627_));
  AOI211_X1 g426(.A(KEYINPUT39), .B(new_n280_), .C1(new_n595_), .C2(new_n621_), .ZN(new_n628_));
  OAI211_X1 g427(.A(new_n625_), .B(new_n620_), .C1(new_n627_), .C2(new_n628_), .ZN(new_n629_));
  INV_X1    g428(.A(new_n629_), .ZN(new_n630_));
  NOR2_X1   g429(.A1(new_n626_), .A2(new_n630_), .ZN(G1325gat));
  INV_X1    g430(.A(G15gat), .ZN(new_n632_));
  NAND3_X1  g431(.A1(new_n614_), .A2(new_n632_), .A3(new_n583_), .ZN(new_n633_));
  OAI21_X1  g432(.A(G15gat), .B1(new_n596_), .B2(new_n582_), .ZN(new_n634_));
  INV_X1    g433(.A(KEYINPUT41), .ZN(new_n635_));
  AND2_X1   g434(.A1(new_n634_), .A2(new_n635_), .ZN(new_n636_));
  NOR2_X1   g435(.A1(new_n634_), .A2(new_n635_), .ZN(new_n637_));
  OAI21_X1  g436(.A(new_n633_), .B1(new_n636_), .B2(new_n637_), .ZN(G1326gat));
  INV_X1    g437(.A(G22gat), .ZN(new_n639_));
  AOI21_X1  g438(.A(new_n639_), .B1(new_n595_), .B2(new_n585_), .ZN(new_n640_));
  XOR2_X1   g439(.A(new_n640_), .B(KEYINPUT42), .Z(new_n641_));
  NAND3_X1  g440(.A1(new_n614_), .A2(new_n639_), .A3(new_n585_), .ZN(new_n642_));
  NAND2_X1  g441(.A1(new_n641_), .A2(new_n642_), .ZN(G1327gat));
  NOR2_X1   g442(.A1(new_n346_), .A2(new_n292_), .ZN(new_n644_));
  NAND2_X1  g443(.A1(new_n602_), .A2(new_n644_), .ZN(new_n645_));
  OR3_X1    g444(.A1(new_n645_), .A2(G29gat), .A3(new_n519_), .ZN(new_n646_));
  NAND3_X1  g445(.A1(new_n273_), .A2(new_n612_), .A3(new_n313_), .ZN(new_n647_));
  XNOR2_X1  g446(.A(new_n647_), .B(KEYINPUT99), .ZN(new_n648_));
  INV_X1    g447(.A(KEYINPUT43), .ZN(new_n649_));
  AND3_X1   g448(.A1(new_n594_), .A2(new_n649_), .A3(new_n611_), .ZN(new_n650_));
  AOI21_X1  g449(.A(new_n649_), .B1(new_n594_), .B2(new_n611_), .ZN(new_n651_));
  OAI21_X1  g450(.A(new_n648_), .B1(new_n650_), .B2(new_n651_), .ZN(new_n652_));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653_));
  NAND2_X1  g452(.A1(new_n652_), .A2(new_n653_), .ZN(new_n654_));
  OAI211_X1 g453(.A(new_n648_), .B(KEYINPUT44), .C1(new_n650_), .C2(new_n651_), .ZN(new_n655_));
  NAND3_X1  g454(.A1(new_n654_), .A2(new_n615_), .A3(new_n655_), .ZN(new_n656_));
  INV_X1    g455(.A(KEYINPUT100), .ZN(new_n657_));
  AND3_X1   g456(.A1(new_n656_), .A2(new_n657_), .A3(G29gat), .ZN(new_n658_));
  AOI21_X1  g457(.A(new_n657_), .B1(new_n656_), .B2(G29gat), .ZN(new_n659_));
  OAI21_X1  g458(.A(new_n646_), .B1(new_n658_), .B2(new_n659_), .ZN(G1328gat));
  INV_X1    g459(.A(KEYINPUT46), .ZN(new_n661_));
  AOI21_X1  g460(.A(KEYINPUT102), .B1(new_n661_), .B2(KEYINPUT101), .ZN(new_n662_));
  INV_X1    g461(.A(new_n662_), .ZN(new_n663_));
  NAND3_X1  g462(.A1(new_n654_), .A2(new_n621_), .A3(new_n655_), .ZN(new_n664_));
  NAND2_X1  g463(.A1(new_n664_), .A2(G36gat), .ZN(new_n665_));
  NAND2_X1  g464(.A1(new_n661_), .A2(KEYINPUT102), .ZN(new_n666_));
  NOR2_X1   g465(.A1(new_n590_), .A2(G36gat), .ZN(new_n667_));
  NAND4_X1  g466(.A1(new_n594_), .A2(new_n601_), .A3(new_n644_), .A4(new_n667_), .ZN(new_n668_));
  AND2_X1   g467(.A1(new_n668_), .A2(KEYINPUT45), .ZN(new_n669_));
  NOR2_X1   g468(.A1(new_n668_), .A2(KEYINPUT45), .ZN(new_n670_));
  OAI21_X1  g469(.A(new_n666_), .B1(new_n669_), .B2(new_n670_), .ZN(new_n671_));
  INV_X1    g470(.A(new_n671_), .ZN(new_n672_));
  AOI21_X1  g471(.A(new_n663_), .B1(new_n665_), .B2(new_n672_), .ZN(new_n673_));
  AOI211_X1 g472(.A(new_n662_), .B(new_n671_), .C1(new_n664_), .C2(G36gat), .ZN(new_n674_));
  NOR2_X1   g473(.A1(new_n673_), .A2(new_n674_), .ZN(G1329gat));
  NAND4_X1  g474(.A1(new_n654_), .A2(G43gat), .A3(new_n583_), .A4(new_n655_), .ZN(new_n676_));
  INV_X1    g475(.A(G43gat), .ZN(new_n677_));
  OAI21_X1  g476(.A(new_n677_), .B1(new_n645_), .B2(new_n582_), .ZN(new_n678_));
  NAND2_X1  g477(.A1(new_n676_), .A2(new_n678_), .ZN(new_n679_));
  XNOR2_X1  g478(.A(new_n679_), .B(KEYINPUT47), .ZN(G1330gat));
  OR3_X1    g479(.A1(new_n645_), .A2(G50gat), .A3(new_n551_), .ZN(new_n681_));
  NAND3_X1  g480(.A1(new_n654_), .A2(new_n585_), .A3(new_n655_), .ZN(new_n682_));
  INV_X1    g481(.A(KEYINPUT103), .ZN(new_n683_));
  AND2_X1   g482(.A1(new_n682_), .A2(new_n683_), .ZN(new_n684_));
  OAI21_X1  g483(.A(G50gat), .B1(new_n682_), .B2(new_n683_), .ZN(new_n685_));
  OAI21_X1  g484(.A(new_n681_), .B1(new_n684_), .B2(new_n685_), .ZN(G1331gat));
  AND3_X1   g485(.A1(new_n594_), .A2(new_n600_), .A3(new_n599_), .ZN(new_n687_));
  INV_X1    g486(.A(new_n346_), .ZN(new_n688_));
  NOR2_X1   g487(.A1(new_n688_), .A2(new_n612_), .ZN(new_n689_));
  NAND4_X1  g488(.A1(new_n687_), .A2(G57gat), .A3(new_n615_), .A4(new_n689_), .ZN(new_n690_));
  XOR2_X1   g489(.A(new_n690_), .B(KEYINPUT104), .Z(new_n691_));
  NAND2_X1  g490(.A1(new_n687_), .A2(new_n613_), .ZN(new_n692_));
  INV_X1    g491(.A(new_n692_), .ZN(new_n693_));
  AOI21_X1  g492(.A(G57gat), .B1(new_n693_), .B2(new_n615_), .ZN(new_n694_));
  NOR2_X1   g493(.A1(new_n691_), .A2(new_n694_), .ZN(G1332gat));
  NAND2_X1  g494(.A1(new_n687_), .A2(new_n689_), .ZN(new_n696_));
  OAI21_X1  g495(.A(G64gat), .B1(new_n696_), .B2(new_n590_), .ZN(new_n697_));
  XNOR2_X1  g496(.A(new_n697_), .B(KEYINPUT48), .ZN(new_n698_));
  NOR2_X1   g497(.A1(new_n590_), .A2(G64gat), .ZN(new_n699_));
  XOR2_X1   g498(.A(new_n699_), .B(KEYINPUT105), .Z(new_n700_));
  OAI21_X1  g499(.A(new_n698_), .B1(new_n692_), .B2(new_n700_), .ZN(G1333gat));
  OR3_X1    g500(.A1(new_n692_), .A2(G71gat), .A3(new_n582_), .ZN(new_n702_));
  OAI21_X1  g501(.A(G71gat), .B1(new_n696_), .B2(new_n582_), .ZN(new_n703_));
  AND2_X1   g502(.A1(new_n703_), .A2(KEYINPUT49), .ZN(new_n704_));
  NOR2_X1   g503(.A1(new_n703_), .A2(KEYINPUT49), .ZN(new_n705_));
  OAI21_X1  g504(.A(new_n702_), .B1(new_n704_), .B2(new_n705_), .ZN(new_n706_));
  INV_X1    g505(.A(KEYINPUT106), .ZN(new_n707_));
  NAND2_X1  g506(.A1(new_n706_), .A2(new_n707_), .ZN(new_n708_));
  OAI211_X1 g507(.A(KEYINPUT106), .B(new_n702_), .C1(new_n704_), .C2(new_n705_), .ZN(new_n709_));
  NAND2_X1  g508(.A1(new_n708_), .A2(new_n709_), .ZN(G1334gat));
  OAI21_X1  g509(.A(G78gat), .B1(new_n696_), .B2(new_n551_), .ZN(new_n711_));
  XNOR2_X1  g510(.A(new_n711_), .B(KEYINPUT50), .ZN(new_n712_));
  NAND3_X1  g511(.A1(new_n693_), .A2(new_n467_), .A3(new_n585_), .ZN(new_n713_));
  NAND2_X1  g512(.A1(new_n712_), .A2(new_n713_), .ZN(G1335gat));
  AND2_X1   g513(.A1(new_n687_), .A2(new_n644_), .ZN(new_n715_));
  NAND3_X1  g514(.A1(new_n715_), .A2(new_n208_), .A3(new_n615_), .ZN(new_n716_));
  OR2_X1    g515(.A1(new_n650_), .A2(new_n651_), .ZN(new_n717_));
  NOR3_X1   g516(.A1(new_n273_), .A2(new_n292_), .A3(new_n313_), .ZN(new_n718_));
  NAND3_X1  g517(.A1(new_n717_), .A2(new_n615_), .A3(new_n718_), .ZN(new_n719_));
  INV_X1    g518(.A(new_n719_), .ZN(new_n720_));
  OAI21_X1  g519(.A(new_n716_), .B1(new_n720_), .B2(new_n208_), .ZN(G1336gat));
  NAND3_X1  g520(.A1(new_n717_), .A2(new_n621_), .A3(new_n718_), .ZN(new_n722_));
  NAND2_X1  g521(.A1(new_n722_), .A2(G92gat), .ZN(new_n723_));
  NAND3_X1  g522(.A1(new_n715_), .A2(new_n209_), .A3(new_n621_), .ZN(new_n724_));
  NAND2_X1  g523(.A1(new_n723_), .A2(new_n724_), .ZN(new_n725_));
  INV_X1    g524(.A(KEYINPUT107), .ZN(new_n726_));
  NAND2_X1  g525(.A1(new_n725_), .A2(new_n726_), .ZN(new_n727_));
  NAND3_X1  g526(.A1(new_n723_), .A2(KEYINPUT107), .A3(new_n724_), .ZN(new_n728_));
  NAND2_X1  g527(.A1(new_n727_), .A2(new_n728_), .ZN(G1337gat));
  OAI211_X1 g528(.A(new_n718_), .B(new_n583_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n730_));
  AND2_X1   g529(.A1(new_n583_), .A2(new_n203_), .ZN(new_n731_));
  AOI22_X1  g530(.A1(new_n730_), .A2(G99gat), .B1(new_n715_), .B2(new_n731_), .ZN(new_n732_));
  NOR2_X1   g531(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n733_));
  NOR2_X1   g532(.A1(new_n732_), .A2(new_n733_), .ZN(new_n734_));
  AND2_X1   g533(.A1(KEYINPUT108), .A2(KEYINPUT51), .ZN(new_n735_));
  XNOR2_X1  g534(.A(new_n734_), .B(new_n735_), .ZN(G1338gat));
  NAND3_X1  g535(.A1(new_n715_), .A2(new_n204_), .A3(new_n585_), .ZN(new_n737_));
  OAI211_X1 g536(.A(new_n718_), .B(new_n585_), .C1(new_n650_), .C2(new_n651_), .ZN(new_n738_));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739_));
  AND3_X1   g538(.A1(new_n738_), .A2(new_n739_), .A3(G106gat), .ZN(new_n740_));
  AOI21_X1  g539(.A(new_n739_), .B1(new_n738_), .B2(G106gat), .ZN(new_n741_));
  OAI21_X1  g540(.A(new_n737_), .B1(new_n740_), .B2(new_n741_), .ZN(new_n742_));
  NAND2_X1  g541(.A1(new_n742_), .A2(KEYINPUT53), .ZN(new_n743_));
  INV_X1    g542(.A(KEYINPUT53), .ZN(new_n744_));
  OAI211_X1 g543(.A(new_n744_), .B(new_n737_), .C1(new_n740_), .C2(new_n741_), .ZN(new_n745_));
  NAND2_X1  g544(.A1(new_n743_), .A2(new_n745_), .ZN(G1339gat));
  INV_X1    g545(.A(KEYINPUT113), .ZN(new_n747_));
  INV_X1    g546(.A(G113gat), .ZN(new_n748_));
  NOR3_X1   g547(.A1(new_n591_), .A2(new_n582_), .A3(new_n519_), .ZN(new_n749_));
  INV_X1    g548(.A(KEYINPUT59), .ZN(new_n750_));
  NAND2_X1  g549(.A1(new_n749_), .A2(new_n750_), .ZN(new_n751_));
  NAND2_X1  g550(.A1(new_n313_), .A2(new_n262_), .ZN(new_n752_));
  INV_X1    g551(.A(KEYINPUT55), .ZN(new_n753_));
  AOI21_X1  g552(.A(new_n237_), .B1(new_n228_), .B2(new_n229_), .ZN(new_n754_));
  OAI211_X1 g553(.A(new_n254_), .B(new_n238_), .C1(new_n754_), .C2(KEYINPUT12), .ZN(new_n755_));
  AOI21_X1  g554(.A(new_n753_), .B1(new_n755_), .B2(new_n250_), .ZN(new_n756_));
  NOR2_X1   g555(.A1(new_n755_), .A2(new_n250_), .ZN(new_n757_));
  NOR2_X1   g556(.A1(new_n756_), .A2(new_n757_), .ZN(new_n758_));
  NOR3_X1   g557(.A1(new_n755_), .A2(new_n753_), .A3(new_n250_), .ZN(new_n759_));
  OAI21_X1  g558(.A(new_n267_), .B1(new_n758_), .B2(new_n759_), .ZN(new_n760_));
  INV_X1    g559(.A(KEYINPUT56), .ZN(new_n761_));
  NAND2_X1  g560(.A1(new_n760_), .A2(new_n761_), .ZN(new_n762_));
  OAI211_X1 g561(.A(KEYINPUT56), .B(new_n267_), .C1(new_n758_), .C2(new_n759_), .ZN(new_n763_));
  AOI21_X1  g562(.A(new_n752_), .B1(new_n762_), .B2(new_n763_), .ZN(new_n764_));
  NOR2_X1   g563(.A1(new_n308_), .A2(new_n312_), .ZN(new_n765_));
  INV_X1    g564(.A(new_n312_), .ZN(new_n766_));
  AOI21_X1  g565(.A(new_n766_), .B1(new_n299_), .B2(new_n300_), .ZN(new_n767_));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n768_));
  OR2_X1    g567(.A1(new_n767_), .A2(new_n768_), .ZN(new_n769_));
  AOI22_X1  g568(.A1(new_n767_), .A2(new_n768_), .B1(new_n301_), .B2(new_n306_), .ZN(new_n770_));
  AOI21_X1  g569(.A(new_n765_), .B1(new_n769_), .B2(new_n770_), .ZN(new_n771_));
  AND3_X1   g570(.A1(new_n265_), .A2(new_n269_), .A3(new_n771_), .ZN(new_n772_));
  OAI21_X1  g571(.A(new_n346_), .B1(new_n764_), .B2(new_n772_), .ZN(new_n773_));
  INV_X1    g572(.A(KEYINPUT110), .ZN(new_n774_));
  OAI21_X1  g573(.A(new_n773_), .B1(new_n774_), .B2(KEYINPUT57), .ZN(new_n775_));
  NOR2_X1   g574(.A1(new_n774_), .A2(KEYINPUT57), .ZN(new_n776_));
  OAI211_X1 g575(.A(new_n346_), .B(new_n776_), .C1(new_n764_), .C2(new_n772_), .ZN(new_n777_));
  NAND2_X1  g576(.A1(new_n775_), .A2(new_n777_), .ZN(new_n778_));
  NAND2_X1  g577(.A1(new_n763_), .A2(KEYINPUT111), .ZN(new_n779_));
  AOI21_X1  g578(.A(new_n249_), .B1(new_n253_), .B2(new_n255_), .ZN(new_n780_));
  OAI21_X1  g579(.A(new_n256_), .B1(new_n780_), .B2(new_n753_), .ZN(new_n781_));
  INV_X1    g580(.A(new_n759_), .ZN(new_n782_));
  NAND2_X1  g581(.A1(new_n781_), .A2(new_n782_), .ZN(new_n783_));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n784_));
  NAND4_X1  g583(.A1(new_n783_), .A2(new_n784_), .A3(KEYINPUT56), .A4(new_n267_), .ZN(new_n785_));
  NAND3_X1  g584(.A1(new_n779_), .A2(new_n785_), .A3(new_n762_), .ZN(new_n786_));
  AND2_X1   g585(.A1(new_n771_), .A2(new_n262_), .ZN(new_n787_));
  NAND2_X1  g586(.A1(new_n786_), .A2(new_n787_), .ZN(new_n788_));
  INV_X1    g587(.A(KEYINPUT58), .ZN(new_n789_));
  NAND2_X1  g588(.A1(new_n788_), .A2(new_n789_), .ZN(new_n790_));
  NAND3_X1  g589(.A1(new_n786_), .A2(KEYINPUT58), .A3(new_n787_), .ZN(new_n791_));
  NAND3_X1  g590(.A1(new_n611_), .A2(new_n790_), .A3(new_n791_), .ZN(new_n792_));
  AOI21_X1  g591(.A(new_n292_), .B1(new_n778_), .B2(new_n792_), .ZN(new_n793_));
  INV_X1    g592(.A(new_n793_), .ZN(new_n794_));
  NOR3_X1   g593(.A1(new_n271_), .A2(new_n272_), .A3(new_n313_), .ZN(new_n795_));
  NAND4_X1  g594(.A1(new_n795_), .A2(new_n608_), .A3(new_n610_), .A4(new_n292_), .ZN(new_n796_));
  XNOR2_X1  g595(.A(new_n796_), .B(KEYINPUT54), .ZN(new_n797_));
  AOI21_X1  g596(.A(new_n751_), .B1(new_n794_), .B2(new_n797_), .ZN(new_n798_));
  AOI22_X1  g597(.A1(new_n792_), .A2(KEYINPUT112), .B1(new_n775_), .B2(new_n777_), .ZN(new_n799_));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800_));
  NAND4_X1  g599(.A1(new_n611_), .A2(new_n790_), .A3(new_n800_), .A4(new_n791_), .ZN(new_n801_));
  AOI21_X1  g600(.A(new_n292_), .B1(new_n799_), .B2(new_n801_), .ZN(new_n802_));
  INV_X1    g601(.A(KEYINPUT54), .ZN(new_n803_));
  XNOR2_X1  g602(.A(new_n796_), .B(new_n803_), .ZN(new_n804_));
  OAI21_X1  g603(.A(new_n749_), .B1(new_n802_), .B2(new_n804_), .ZN(new_n805_));
  AOI21_X1  g604(.A(new_n798_), .B1(new_n805_), .B2(KEYINPUT59), .ZN(new_n806_));
  AOI21_X1  g605(.A(new_n748_), .B1(new_n806_), .B2(new_n313_), .ZN(new_n807_));
  NOR3_X1   g606(.A1(new_n805_), .A2(G113gat), .A3(new_n600_), .ZN(new_n808_));
  OAI21_X1  g607(.A(new_n747_), .B1(new_n807_), .B2(new_n808_), .ZN(new_n809_));
  INV_X1    g608(.A(new_n808_), .ZN(new_n810_));
  AOI211_X1 g609(.A(new_n600_), .B(new_n798_), .C1(new_n805_), .C2(KEYINPUT59), .ZN(new_n811_));
  OAI211_X1 g610(.A(KEYINPUT113), .B(new_n810_), .C1(new_n811_), .C2(new_n748_), .ZN(new_n812_));
  NAND2_X1  g611(.A1(new_n809_), .A2(new_n812_), .ZN(G1340gat));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n814_));
  INV_X1    g613(.A(G120gat), .ZN(new_n815_));
  AOI21_X1  g614(.A(new_n815_), .B1(new_n806_), .B2(new_n599_), .ZN(new_n816_));
  OAI21_X1  g615(.A(new_n815_), .B1(new_n273_), .B2(KEYINPUT60), .ZN(new_n817_));
  OAI21_X1  g616(.A(new_n817_), .B1(KEYINPUT60), .B2(new_n815_), .ZN(new_n818_));
  NOR2_X1   g617(.A1(new_n805_), .A2(new_n818_), .ZN(new_n819_));
  OAI21_X1  g618(.A(new_n814_), .B1(new_n816_), .B2(new_n819_), .ZN(new_n820_));
  INV_X1    g619(.A(new_n819_), .ZN(new_n821_));
  AOI211_X1 g620(.A(new_n273_), .B(new_n798_), .C1(new_n805_), .C2(KEYINPUT59), .ZN(new_n822_));
  OAI211_X1 g621(.A(KEYINPUT114), .B(new_n821_), .C1(new_n822_), .C2(new_n815_), .ZN(new_n823_));
  NAND2_X1  g622(.A1(new_n820_), .A2(new_n823_), .ZN(G1341gat));
  INV_X1    g623(.A(new_n805_), .ZN(new_n825_));
  NAND3_X1  g624(.A1(new_n825_), .A2(new_n490_), .A3(new_n292_), .ZN(new_n826_));
  AND2_X1   g625(.A1(new_n806_), .A2(new_n292_), .ZN(new_n827_));
  OAI21_X1  g626(.A(new_n826_), .B1(new_n827_), .B2(new_n490_), .ZN(G1342gat));
  NAND3_X1  g627(.A1(new_n825_), .A2(new_n488_), .A3(new_n688_), .ZN(new_n829_));
  AND2_X1   g628(.A1(new_n806_), .A2(new_n611_), .ZN(new_n830_));
  OAI21_X1  g629(.A(new_n829_), .B1(new_n830_), .B2(new_n488_), .ZN(G1343gat));
  NOR2_X1   g630(.A1(new_n802_), .A2(new_n804_), .ZN(new_n832_));
  NAND4_X1  g631(.A1(new_n582_), .A2(new_n590_), .A3(new_n615_), .A4(new_n585_), .ZN(new_n833_));
  XOR2_X1   g632(.A(new_n833_), .B(KEYINPUT115), .Z(new_n834_));
  INV_X1    g633(.A(new_n834_), .ZN(new_n835_));
  NOR2_X1   g634(.A1(new_n832_), .A2(new_n835_), .ZN(new_n836_));
  NAND2_X1  g635(.A1(new_n836_), .A2(new_n313_), .ZN(new_n837_));
  XNOR2_X1  g636(.A(new_n837_), .B(G141gat), .ZN(G1344gat));
  NAND2_X1  g637(.A1(new_n836_), .A2(new_n599_), .ZN(new_n839_));
  XNOR2_X1  g638(.A(new_n839_), .B(G148gat), .ZN(G1345gat));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n841_));
  AOI21_X1  g640(.A(new_n841_), .B1(new_n836_), .B2(new_n292_), .ZN(new_n842_));
  INV_X1    g641(.A(new_n842_), .ZN(new_n843_));
  NOR4_X1   g642(.A1(new_n832_), .A2(KEYINPUT116), .A3(new_n612_), .A4(new_n835_), .ZN(new_n844_));
  INV_X1    g643(.A(new_n844_), .ZN(new_n845_));
  XNOR2_X1  g644(.A(KEYINPUT61), .B(G155gat), .ZN(new_n846_));
  NAND3_X1  g645(.A1(new_n843_), .A2(new_n845_), .A3(new_n846_), .ZN(new_n847_));
  INV_X1    g646(.A(new_n846_), .ZN(new_n848_));
  OAI21_X1  g647(.A(new_n848_), .B1(new_n842_), .B2(new_n844_), .ZN(new_n849_));
  NAND2_X1  g648(.A1(new_n847_), .A2(new_n849_), .ZN(G1346gat));
  INV_X1    g649(.A(new_n836_), .ZN(new_n851_));
  INV_X1    g650(.A(new_n611_), .ZN(new_n852_));
  OAI21_X1  g651(.A(G162gat), .B1(new_n851_), .B2(new_n852_), .ZN(new_n853_));
  OR2_X1    g652(.A1(new_n346_), .A2(G162gat), .ZN(new_n854_));
  OAI21_X1  g653(.A(new_n853_), .B1(new_n851_), .B2(new_n854_), .ZN(G1347gat));
  INV_X1    g654(.A(KEYINPUT121), .ZN(new_n856_));
  OR3_X1    g655(.A1(new_n592_), .A2(KEYINPUT117), .A3(new_n590_), .ZN(new_n857_));
  OAI21_X1  g656(.A(KEYINPUT117), .B1(new_n592_), .B2(new_n590_), .ZN(new_n858_));
  NAND2_X1  g657(.A1(new_n857_), .A2(new_n858_), .ZN(new_n859_));
  AOI21_X1  g658(.A(KEYINPUT118), .B1(new_n859_), .B2(new_n313_), .ZN(new_n860_));
  INV_X1    g659(.A(KEYINPUT118), .ZN(new_n861_));
  AOI211_X1 g660(.A(new_n861_), .B(new_n600_), .C1(new_n857_), .C2(new_n858_), .ZN(new_n862_));
  NOR2_X1   g661(.A1(new_n860_), .A2(new_n862_), .ZN(new_n863_));
  OAI211_X1 g662(.A(new_n863_), .B(new_n551_), .C1(new_n804_), .C2(new_n793_), .ZN(new_n864_));
  NAND3_X1  g663(.A1(new_n864_), .A2(KEYINPUT119), .A3(G169gat), .ZN(new_n865_));
  NAND2_X1  g664(.A1(new_n865_), .A2(KEYINPUT62), .ZN(new_n866_));
  AOI21_X1  g665(.A(KEYINPUT119), .B1(new_n864_), .B2(G169gat), .ZN(new_n867_));
  NOR2_X1   g666(.A1(new_n866_), .A2(new_n867_), .ZN(new_n868_));
  NAND2_X1  g667(.A1(new_n864_), .A2(G169gat), .ZN(new_n869_));
  INV_X1    g668(.A(KEYINPUT119), .ZN(new_n870_));
  INV_X1    g669(.A(KEYINPUT62), .ZN(new_n871_));
  NAND3_X1  g670(.A1(new_n869_), .A2(new_n870_), .A3(new_n871_), .ZN(new_n872_));
  INV_X1    g671(.A(new_n859_), .ZN(new_n873_));
  AOI211_X1 g672(.A(new_n585_), .B(new_n873_), .C1(new_n794_), .C2(new_n797_), .ZN(new_n874_));
  NAND2_X1  g673(.A1(new_n313_), .A2(new_n374_), .ZN(new_n875_));
  XNOR2_X1  g674(.A(new_n875_), .B(KEYINPUT120), .ZN(new_n876_));
  NAND2_X1  g675(.A1(new_n874_), .A2(new_n876_), .ZN(new_n877_));
  NAND2_X1  g676(.A1(new_n872_), .A2(new_n877_), .ZN(new_n878_));
  OAI21_X1  g677(.A(new_n856_), .B1(new_n868_), .B2(new_n878_), .ZN(new_n879_));
  NAND2_X1  g678(.A1(new_n869_), .A2(new_n870_), .ZN(new_n880_));
  NAND3_X1  g679(.A1(new_n880_), .A2(KEYINPUT62), .A3(new_n865_), .ZN(new_n881_));
  NAND4_X1  g680(.A1(new_n881_), .A2(KEYINPUT121), .A3(new_n872_), .A4(new_n877_), .ZN(new_n882_));
  NAND2_X1  g681(.A1(new_n879_), .A2(new_n882_), .ZN(G1348gat));
  AOI21_X1  g682(.A(G176gat), .B1(new_n874_), .B2(new_n599_), .ZN(new_n884_));
  NOR2_X1   g683(.A1(new_n832_), .A2(new_n585_), .ZN(new_n885_));
  NOR3_X1   g684(.A1(new_n873_), .A2(new_n375_), .A3(new_n273_), .ZN(new_n886_));
  AOI21_X1  g685(.A(new_n884_), .B1(new_n885_), .B2(new_n886_), .ZN(G1349gat));
  NAND3_X1  g686(.A1(new_n885_), .A2(new_n292_), .A3(new_n859_), .ZN(new_n888_));
  NOR2_X1   g687(.A1(new_n612_), .A2(new_n368_), .ZN(new_n889_));
  AOI22_X1  g688(.A1(new_n888_), .A2(new_n358_), .B1(new_n874_), .B2(new_n889_), .ZN(G1350gat));
  NAND3_X1  g689(.A1(new_n874_), .A2(new_n688_), .A3(new_n369_), .ZN(new_n891_));
  NAND2_X1  g690(.A1(new_n874_), .A2(new_n611_), .ZN(new_n892_));
  AND3_X1   g691(.A1(new_n892_), .A2(KEYINPUT122), .A3(G190gat), .ZN(new_n893_));
  AOI21_X1  g692(.A(KEYINPUT122), .B1(new_n892_), .B2(G190gat), .ZN(new_n894_));
  OAI21_X1  g693(.A(new_n891_), .B1(new_n893_), .B2(new_n894_), .ZN(G1351gat));
  NOR3_X1   g694(.A1(new_n583_), .A2(new_n590_), .A3(new_n525_), .ZN(new_n896_));
  OAI211_X1 g695(.A(new_n313_), .B(new_n896_), .C1(new_n802_), .C2(new_n804_), .ZN(new_n897_));
  AND2_X1   g696(.A1(new_n897_), .A2(new_n348_), .ZN(new_n898_));
  OR2_X1    g697(.A1(new_n898_), .A2(KEYINPUT124), .ZN(new_n899_));
  NAND2_X1  g698(.A1(new_n898_), .A2(KEYINPUT124), .ZN(new_n900_));
  OAI21_X1  g699(.A(KEYINPUT123), .B1(new_n897_), .B2(new_n348_), .ZN(new_n901_));
  OR3_X1    g700(.A1(new_n897_), .A2(KEYINPUT123), .A3(new_n348_), .ZN(new_n902_));
  AOI22_X1  g701(.A1(new_n899_), .A2(new_n900_), .B1(new_n901_), .B2(new_n902_), .ZN(G1352gat));
  INV_X1    g702(.A(new_n896_), .ZN(new_n904_));
  NOR2_X1   g703(.A1(new_n832_), .A2(new_n904_), .ZN(new_n905_));
  NAND2_X1  g704(.A1(new_n905_), .A2(new_n599_), .ZN(new_n906_));
  INV_X1    g705(.A(KEYINPUT125), .ZN(new_n907_));
  OAI21_X1  g706(.A(new_n906_), .B1(new_n907_), .B2(G204gat), .ZN(new_n908_));
  XNOR2_X1  g707(.A(KEYINPUT125), .B(G204gat), .ZN(new_n909_));
  OAI21_X1  g708(.A(new_n908_), .B1(new_n906_), .B2(new_n909_), .ZN(G1353gat));
  NOR3_X1   g709(.A1(new_n832_), .A2(new_n612_), .A3(new_n904_), .ZN(new_n911_));
  INV_X1    g710(.A(KEYINPUT126), .ZN(new_n912_));
  XOR2_X1   g711(.A(KEYINPUT63), .B(G211gat), .Z(new_n913_));
  NAND3_X1  g712(.A1(new_n911_), .A2(new_n912_), .A3(new_n913_), .ZN(new_n914_));
  NAND2_X1  g713(.A1(new_n911_), .A2(new_n913_), .ZN(new_n915_));
  NAND2_X1  g714(.A1(new_n915_), .A2(KEYINPUT126), .ZN(new_n916_));
  NOR3_X1   g715(.A1(new_n911_), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n917_));
  OAI21_X1  g716(.A(new_n914_), .B1(new_n916_), .B2(new_n917_), .ZN(G1354gat));
  AOI21_X1  g717(.A(G218gat), .B1(new_n905_), .B2(new_n688_), .ZN(new_n919_));
  NAND2_X1  g718(.A1(new_n611_), .A2(G218gat), .ZN(new_n920_));
  XNOR2_X1  g719(.A(new_n920_), .B(KEYINPUT127), .ZN(new_n921_));
  AOI21_X1  g720(.A(new_n919_), .B1(new_n905_), .B2(new_n921_), .ZN(G1355gat));
endmodule


